magic
tech sky130A
magscale 1 2
timestamp 1607618424
<< locali >>
rect 429485 666587 429519 684437
rect 494069 666587 494103 676141
rect 559297 666587 559331 684437
rect 429209 647275 429243 656829
rect 559205 647275 559239 656829
rect 37415 639557 37473 639591
rect 193263 639557 193413 639591
rect 212675 639557 212733 639591
rect 15209 639319 15243 639421
rect 24777 639319 24811 639489
rect 27629 639319 27663 639489
rect 37197 639319 37231 639489
rect 37289 639319 37323 639489
rect 46949 639319 46983 639489
rect 60657 639455 60691 639489
rect 60657 639421 60841 639455
rect 67649 639387 67683 639489
rect 75929 639319 75963 639489
rect 85497 639319 85531 639421
rect 86969 639387 87003 639489
rect 99297 639455 99331 639489
rect 99297 639421 99481 639455
rect 106289 639387 106323 639489
rect 118617 639455 118651 639489
rect 153243 639489 153611 639523
rect 118617 639421 118801 639455
rect 125609 639387 125643 639489
rect 153577 639455 153611 639489
rect 164249 639387 164283 639489
rect 176577 639455 176611 639489
rect 195931 639489 196023 639523
rect 176577 639421 176761 639455
rect 143583 639353 143641 639387
rect 183569 639387 183603 639489
rect 195989 639455 196023 639489
rect 212549 639455 212583 639489
rect 229661 639455 229695 639829
rect 229753 639591 229787 639761
rect 239321 639591 239355 639829
rect 239413 639591 239447 639761
rect 247601 639591 247635 639761
rect 251833 639591 251867 639829
rect 257905 639591 257939 639829
rect 257997 639591 258031 639761
rect 267749 639591 267783 639829
rect 267841 639591 267875 640033
rect 277225 639591 277259 640033
rect 277317 639591 277351 639829
rect 287069 639591 287103 640033
rect 287161 639591 287195 640101
rect 290565 639591 290599 640101
rect 292589 639591 292623 640033
rect 307033 639591 307067 640033
rect 307125 639591 307159 640237
rect 311817 639591 311851 640237
rect 325801 640203 325835 641665
rect 325801 640169 325927 640203
rect 311909 639591 311943 640033
rect 325801 639591 325835 640033
rect 325893 639591 325927 640169
rect 335185 639591 335219 641665
rect 336013 639591 336047 640033
rect 345029 639591 345063 641665
rect 354597 639591 354631 641665
rect 364349 639591 364383 641665
rect 373917 639591 373951 641665
rect 383669 639591 383703 641665
rect 393237 639591 393271 641665
rect 402989 639591 403023 641665
rect 408359 639625 408509 639659
rect 412557 639591 412591 641665
rect 441629 639591 441663 639693
rect 441721 639591 441755 640645
rect 445217 639591 445251 640645
rect 463709 639591 463743 639693
rect 473277 639591 473311 639693
rect 202889 639319 202923 639421
rect 212549 639421 212641 639455
rect 212457 639319 212491 639421
rect 234663 337705 235031 337739
rect 234997 337535 235031 337705
rect 237481 337603 237515 337705
rect 239413 337535 239447 337637
rect 228097 337399 228131 337501
rect 267473 337399 267507 337501
rect 228097 337365 228281 337399
rect 267565 328491 267599 337501
rect 230673 318835 230707 325533
rect 249993 317475 250027 321657
rect 252661 320127 252695 328389
rect 259653 318835 259687 321589
rect 230673 299523 230707 304249
rect 231961 298163 231995 315945
rect 267105 307819 267139 309145
rect 236285 289731 236319 298061
rect 241805 289867 241839 299421
rect 243001 298163 243035 307717
rect 270693 299523 270727 309077
rect 277593 306391 277627 311865
rect 288633 309179 288667 318733
rect 292773 317475 292807 327029
rect 294061 316047 294095 333897
rect 295625 328491 295659 338045
rect 326353 337195 326387 337909
rect 363245 337399 363279 337705
rect 363337 337467 363371 337705
rect 384221 337467 384255 337773
rect 384313 337603 384347 337909
rect 384405 337535 384439 337705
rect 363429 337399 363463 337433
rect 363245 337365 363463 337399
rect 355977 337127 356011 337297
rect 374561 336787 374595 337433
rect 381461 336787 381495 337433
rect 385049 337331 385083 338113
rect 395445 337943 395479 338113
rect 393881 336855 393915 337909
rect 398757 337331 398791 337909
rect 408509 336991 408543 337229
rect 412925 336923 412959 337433
rect 421021 337195 421055 338045
rect 422953 336855 422987 337841
rect 423045 337263 423079 337433
rect 427553 336855 427587 338045
rect 432153 337399 432187 337569
rect 430497 337059 430531 337161
rect 432613 337127 432647 337365
rect 433441 337331 433475 337501
rect 442181 337331 442215 337841
rect 444021 337535 444055 337841
rect 433349 337195 433383 337297
rect 432521 337025 432889 337059
rect 432521 336991 432555 337025
rect 435833 336787 435867 337025
rect 309425 328491 309459 331245
rect 342637 328491 342671 331245
rect 318993 317475 319027 326145
rect 356529 325703 356563 336685
rect 357633 325839 357667 335257
rect 370053 327131 370087 336685
rect 375573 327131 375607 336685
rect 393145 327131 393179 331245
rect 451473 330531 451507 338045
rect 486341 337399 486375 337773
rect 498945 337671 498979 338045
rect 499773 337331 499807 337637
rect 514033 336787 514067 336957
rect 523601 336855 523635 337501
rect 524061 337195 524095 337433
rect 526729 337195 526763 337569
rect 528695 337161 529857 337195
rect 523693 336991 523727 337161
rect 359013 318835 359047 321589
rect 392133 318835 392167 321589
rect 327273 309179 327307 318733
rect 332793 309179 332827 318733
rect 346593 309179 346627 311797
rect 249901 288439 249935 298061
rect 255513 288439 255547 298061
rect 230857 273275 230891 280109
rect 241805 270555 241839 280109
rect 249901 278783 249935 285821
rect 259653 282795 259687 289765
rect 265265 288439 265299 298061
rect 267013 280211 267047 298061
rect 277593 280211 277627 298061
rect 281641 289867 281675 299421
rect 292773 298231 292807 307717
rect 309333 299523 309367 309077
rect 334449 307819 334483 309145
rect 342453 299591 342487 309009
rect 287253 280211 287287 289765
rect 292681 288439 292715 298061
rect 295717 293267 295751 298061
rect 298385 287079 298419 296633
rect 305193 289867 305227 299421
rect 310713 289867 310747 299421
rect 324513 289867 324547 299353
rect 309333 280211 309367 289697
rect 331413 288439 331447 298061
rect 334265 282795 334299 298061
rect 346593 289867 346627 299421
rect 356529 298163 356563 315945
rect 371341 309315 371375 318733
rect 375757 309111 375791 317373
rect 376861 309315 376895 318733
rect 376861 299523 376895 309077
rect 381277 307819 381311 317373
rect 382289 302107 382323 317373
rect 387901 307819 387935 317373
rect 393237 309179 393271 324173
rect 416881 318835 416915 328389
rect 422401 318835 422435 328389
rect 427921 318835 427955 328389
rect 433717 318835 433751 328389
rect 466561 318835 466595 321589
rect 472081 318835 472115 328389
rect 397745 312171 397779 318733
rect 353493 288439 353527 298061
rect 370145 289731 370179 298061
rect 382473 289867 382507 299421
rect 387901 298163 387935 304861
rect 408785 298163 408819 302209
rect 416881 299523 416915 309077
rect 422493 299931 422527 309077
rect 428013 299523 428047 309077
rect 433441 299523 433475 309077
rect 451565 302107 451599 315945
rect 466561 299523 466595 309077
rect 472081 299523 472115 309077
rect 342545 280279 342579 282897
rect 408785 282795 408819 293029
rect 231869 259471 231903 263585
rect 252753 260899 252787 270453
rect 270601 269127 270635 278681
rect 277685 269127 277719 275077
rect 283113 270555 283147 280109
rect 230949 244171 230983 254405
rect 241805 251243 241839 260797
rect 267013 259471 267047 263585
rect 287253 260899 287287 270453
rect 295441 269127 295475 278681
rect 305193 270555 305227 280109
rect 310713 270555 310747 280109
rect 327273 272187 327307 280109
rect 334357 270623 334391 280109
rect 346593 270555 346627 280109
rect 364533 273207 364567 280109
rect 371433 270555 371467 280109
rect 309333 260899 309367 270385
rect 324421 260899 324455 263585
rect 342545 260899 342579 263585
rect 375481 263483 375515 278681
rect 376953 270555 376987 280109
rect 393237 270555 393271 280109
rect 400505 270555 400539 280109
rect 381093 260899 381127 270385
rect 392133 264299 392167 270453
rect 408785 263483 408819 278681
rect 416881 270555 416915 280109
rect 433625 270555 433659 280109
rect 451565 263483 451599 273717
rect 466561 270555 466595 280109
rect 472081 270555 472115 280109
rect 236285 240227 236319 244273
rect 252753 241519 252787 251141
rect 281917 241587 281951 259369
rect 283113 251243 283147 260797
rect 287253 241519 287287 251141
rect 292957 249747 292991 258009
rect 236285 230571 236319 240057
rect 281917 234583 281951 241417
rect 295441 240091 295475 259369
rect 305193 251243 305227 260797
rect 309333 251243 309367 260729
rect 310713 251243 310747 260797
rect 327273 251243 327307 260797
rect 334357 251311 334391 260797
rect 342453 251243 342487 260729
rect 346593 251243 346627 260797
rect 298201 242675 298235 251141
rect 334357 244171 334391 251141
rect 348065 241519 348099 254609
rect 353585 241519 353619 254609
rect 356437 251107 356471 253997
rect 359013 251311 359047 260797
rect 371433 251243 371467 260797
rect 375573 251243 375607 260797
rect 376953 251243 376987 260797
rect 400505 251243 400539 260797
rect 416881 251243 416915 260797
rect 433625 251243 433659 260797
rect 359013 244171 359047 251141
rect 369961 241519 369995 251141
rect 381093 241519 381127 251073
rect 451565 244171 451599 259369
rect 466561 251243 466595 260797
rect 472081 251243 472115 260797
rect 243185 224247 243219 231693
rect 259653 222207 259687 231761
rect 295533 227783 295567 237337
rect 348065 230367 348099 238697
rect 352021 230367 352055 234617
rect 356437 229211 356471 234685
rect 267105 220847 267139 224961
rect 324421 222275 324455 224961
rect 356437 224927 356471 229041
rect 281917 220847 281951 222173
rect 324421 219555 324455 222105
rect 236285 202895 236319 205581
rect 243093 201467 243127 217957
rect 267013 209831 267047 219385
rect 364441 218059 364475 235909
rect 381093 231863 381127 234685
rect 381185 222207 381219 224961
rect 392133 222207 392167 236725
rect 408693 222207 408727 231761
rect 295441 211123 295475 215373
rect 298293 211259 298327 215441
rect 309333 212551 309367 215305
rect 265173 202827 265207 209729
rect 281733 202827 281767 211089
rect 298293 205615 298327 211089
rect 309425 202895 309459 205649
rect 324421 202895 324455 205649
rect 331413 201535 331447 202929
rect 356437 202827 356471 211089
rect 358921 208403 358955 212585
rect 381093 212551 381127 215373
rect 397653 212551 397687 215305
rect 408693 202895 408727 212449
rect 236285 189091 236319 198645
rect 270785 193171 270819 196061
rect 266461 183379 266495 191777
rect 232145 162911 232179 180761
rect 236377 161483 236411 179333
rect 252845 172567 252879 182121
rect 292773 180863 292807 198645
rect 309333 193239 309367 195993
rect 298293 191879 298327 193205
rect 324421 191879 324455 196061
rect 397653 193239 397687 195993
rect 295625 183583 295659 188445
rect 298385 183583 298419 186473
rect 334449 183583 334483 186405
rect 357541 183583 357575 186405
rect 254133 172567 254167 177293
rect 243093 161483 243127 171037
rect 232145 151827 232179 161381
rect 259653 154615 259687 164169
rect 265265 151827 265299 161381
rect 267013 153187 267047 157437
rect 283113 154955 283147 164169
rect 288633 154955 288667 164169
rect 295533 161483 295567 171037
rect 298293 166991 298327 172465
rect 309333 164203 309367 172465
rect 324513 161483 324547 171037
rect 334357 169779 334391 175865
rect 386613 171139 386647 180761
rect 392133 171139 392167 180761
rect 427921 173927 427955 176681
rect 433625 173927 433659 176613
rect 451657 173927 451691 183481
rect 270693 147611 270727 154513
rect 292773 142171 292807 151725
rect 294061 149107 294095 158661
rect 231961 124219 231995 142069
rect 236469 132515 236503 142069
rect 240149 132515 240183 142069
rect 243093 124219 243127 133841
rect 266461 132515 266495 142069
rect 295625 140811 295659 150365
rect 321753 143599 321787 153153
rect 331413 151827 331447 161381
rect 347973 155771 348007 164169
rect 352021 154547 352055 162809
rect 353493 153255 353527 162809
rect 356437 153255 356471 162809
rect 357633 154615 357667 164169
rect 359013 154615 359047 157301
rect 364533 154615 364567 167637
rect 324605 142171 324639 151725
rect 265357 124627 265391 132413
rect 270693 128299 270727 135201
rect 281641 129047 281675 135201
rect 236377 113203 236411 122757
rect 283113 115991 283147 125545
rect 294061 121499 294095 139349
rect 295533 121499 295567 131053
rect 298385 124219 298419 133773
rect 327181 132515 327215 135269
rect 334357 135167 334391 144857
rect 347973 144823 348007 153153
rect 353493 144823 353527 153085
rect 370053 147611 370087 154513
rect 381001 147611 381035 162809
rect 387993 158015 388027 162809
rect 422401 157335 422435 164169
rect 427921 157335 427955 164169
rect 392133 135303 392167 148325
rect 400505 147611 400539 153153
rect 408693 147611 408727 154513
rect 451657 147611 451691 154513
rect 466561 147611 466595 154445
rect 393237 135303 393271 144857
rect 397745 137955 397779 143497
rect 422401 137955 422435 144857
rect 427921 135303 427955 138057
rect 309333 122859 309367 132413
rect 294153 116603 294187 121329
rect 254133 108987 254167 115889
rect 298385 114563 298419 119357
rect 305193 115991 305227 120717
rect 310713 115991 310747 125545
rect 321753 122859 321787 132413
rect 324421 122859 324455 132413
rect 370053 128299 370087 135201
rect 408693 128299 408727 135201
rect 472081 128299 472115 143497
rect 230857 89675 230891 96577
rect 232145 95251 232179 104805
rect 243185 96747 243219 106165
rect 252753 96679 252787 106165
rect 267013 104975 267047 114461
rect 267013 95251 267047 104805
rect 230949 77299 230983 80121
rect 231961 75939 231995 85493
rect 236285 75939 236319 85493
rect 241805 77299 241839 86921
rect 252753 77299 252787 86853
rect 254133 77299 254167 86853
rect 259653 77299 259687 86853
rect 265173 85595 265207 95149
rect 270877 92531 270911 102085
rect 283113 96679 283147 106233
rect 292773 103615 292807 113101
rect 292681 93891 292715 103445
rect 295625 102187 295659 111741
rect 298201 104907 298235 114393
rect 298385 95251 298419 99433
rect 305193 96679 305227 106233
rect 310713 96679 310747 106233
rect 318993 104907 319027 118745
rect 346593 115991 346627 125545
rect 364533 115991 364567 125545
rect 376953 115991 376987 125545
rect 393237 115991 393271 125545
rect 327181 104907 327215 114461
rect 334357 113203 334391 114529
rect 342453 108987 342487 115889
rect 353585 114563 353619 115957
rect 400321 114563 400355 124117
rect 422401 118643 422435 125545
rect 427921 118643 427955 125545
rect 433625 118643 433659 125545
rect 451473 114563 451507 124117
rect 466653 114563 466687 124117
rect 298385 85595 298419 89709
rect 230949 66283 230983 75837
rect 236285 67643 236319 70329
rect 236377 47039 236411 66181
rect 270693 64923 270727 82773
rect 243001 55267 243035 64821
rect 244381 46971 244415 56525
rect 249993 46971 250027 56525
rect 255421 46971 255455 56525
rect 259653 48331 259687 59721
rect 260849 55267 260883 64821
rect 271981 63563 272015 73117
rect 277409 70363 277443 77197
rect 298293 67643 298327 80733
rect 305193 77299 305227 86921
rect 308045 77299 308079 86921
rect 309333 77299 309367 86921
rect 310713 77299 310747 86921
rect 324513 85595 324547 95149
rect 327273 85595 327307 95149
rect 334357 93891 334391 103445
rect 346593 96679 346627 106233
rect 356437 104975 356471 114461
rect 370145 106335 370179 109021
rect 353493 95251 353527 104805
rect 356437 95251 356471 104805
rect 376953 96679 376987 106233
rect 387993 104907 388027 114461
rect 408693 95251 408727 104805
rect 422401 99331 422435 106233
rect 427921 99331 427955 106233
rect 451565 95251 451599 104805
rect 331413 77299 331447 86853
rect 334357 77299 334391 86853
rect 342453 77299 342487 86921
rect 346593 80767 346627 86921
rect 270601 46971 270635 57545
rect 271981 45611 272015 58565
rect 281733 56627 281767 66181
rect 308045 57987 308079 67541
rect 319085 66283 319119 67609
rect 327181 66283 327215 75837
rect 353585 66283 353619 75837
rect 282929 47039 282963 56525
rect 288541 48331 288575 57885
rect 292773 45611 292807 55165
rect 298293 46971 298327 56525
rect 309425 48399 309459 66045
rect 330033 64991 330067 66249
rect 243001 35955 243035 45509
rect 252753 29019 252787 37349
rect 255513 27591 255547 44829
rect 267013 35955 267047 45509
rect 272073 37247 272107 38709
rect 277593 35955 277627 45509
rect 282929 27659 282963 45509
rect 292773 35955 292807 37145
rect 294153 29087 294187 38573
rect 298385 32419 298419 42041
rect 308137 38675 308171 48229
rect 318993 46971 319027 59993
rect 324421 55335 324455 57885
rect 309333 29019 309367 42041
rect 310529 41395 310563 46869
rect 324513 45611 324547 55165
rect 329941 53839 329975 63461
rect 331413 48331 331447 55641
rect 332885 55199 332919 63461
rect 334357 48331 334391 55641
rect 336933 46971 336967 56525
rect 352021 53839 352055 58089
rect 356437 57987 356471 67541
rect 357541 64923 357575 74477
rect 359013 73219 359047 82773
rect 364533 77299 364567 86853
rect 370053 77299 370087 86853
rect 386613 77299 386647 86853
rect 387993 85595 388027 95149
rect 392133 77299 392167 86853
rect 393237 85595 393271 95149
rect 397653 77299 397687 86921
rect 400321 77299 400355 86921
rect 408785 77299 408819 82093
rect 422401 77299 422435 86921
rect 427921 77299 427955 86921
rect 433441 77299 433475 86921
rect 408785 67643 408819 70397
rect 416881 67643 416915 77197
rect 451473 67643 451507 85493
rect 466561 75939 466595 85493
rect 472081 67643 472115 80733
rect 359105 53839 359139 63461
rect 370053 48331 370087 61081
rect 371433 56695 371467 60605
rect 371433 47039 371467 56525
rect 375573 48331 375607 61081
rect 382381 48331 382415 57885
rect 387993 56627 388027 66181
rect 393237 57987 393271 67541
rect 397653 57987 397687 67541
rect 408785 57987 408819 62781
rect 451473 60707 451507 66181
rect 392133 47039 392167 56525
rect 400413 48399 400447 51153
rect 408785 48399 408819 51153
rect 416881 48399 416915 57885
rect 433625 48331 433659 57885
rect 466469 56627 466503 66181
rect 451657 46971 451691 56525
rect 472081 48331 472115 57885
rect 332701 35955 332735 45509
rect 342453 37315 342487 46869
rect 359013 35955 359047 45509
rect 369961 38607 369995 41429
rect 375481 37315 375515 41565
rect 387901 37315 387935 46869
rect 408785 38539 408819 46869
rect 230673 8347 230707 26197
rect 252845 18003 252879 27557
rect 259837 18003 259871 27557
rect 270693 14739 270727 22593
rect 271981 18003 272015 27557
rect 277501 16643 277535 26197
rect 293969 18003 294003 27557
rect 305101 19363 305135 22185
rect 308045 19363 308079 28917
rect 321661 18003 321695 27557
rect 334357 26299 334391 35853
rect 400689 29087 400723 31773
rect 416881 29019 416915 38573
rect 387809 27659 387843 27761
rect 336841 18003 336875 27557
rect 346409 22763 346443 27557
rect 232789 11747 232823 12461
rect 260941 11747 260975 12529
rect 293969 11883 294003 12461
rect 347881 12427 347915 22729
rect 353677 19295 353711 27557
rect 359013 18003 359047 27557
rect 393237 19363 393271 28917
rect 422493 27659 422527 38573
rect 433625 37383 433659 41293
rect 433625 27659 433659 37213
rect 472081 29019 472115 38573
rect 400597 18003 400631 27557
rect 451749 19363 451783 28917
rect 346501 8483 346535 9605
rect 381001 8347 381035 17901
rect 382381 8347 382415 17901
rect 315221 5899 315255 6749
rect 322213 5831 322247 6001
rect 277961 3655 277995 3961
rect 278053 3723 278087 3961
rect 278145 3655 278179 3689
rect 277961 3621 278179 3655
rect 238217 3519 238251 3621
rect 278053 3383 278087 3553
rect 280169 3315 280203 4097
rect 384313 3723 384347 3961
rect 391213 3927 391247 4097
rect 392961 3859 392995 4029
rect 292589 3315 292623 3553
rect 302157 3315 302191 3485
rect 374653 3451 374687 3689
rect 335185 3179 335219 3281
rect 82921 2975 82955 3145
rect 363245 3111 363279 3281
rect 98653 2839 98687 2941
rect 369869 2907 369903 3145
rect 374745 2975 374779 3417
rect 121503 2873 121653 2907
rect 393053 595 393087 9605
rect 400413 8347 400447 17833
rect 416973 12291 417007 19261
rect 393881 3247 393915 4097
rect 393973 3383 394007 4029
rect 400045 3859 400079 4029
rect 403265 3723 403299 4301
rect 403357 3859 403391 4165
rect 403449 3961 403725 3995
rect 402437 3247 402471 3417
rect 403449 3315 403483 3961
rect 408233 3723 408267 4233
rect 408325 3995 408359 4165
rect 408417 3995 408451 4301
rect 408543 4029 409245 4063
rect 403541 3689 403725 3723
rect 403541 3451 403575 3689
rect 408417 3451 408451 3621
rect 409245 3417 409889 3451
rect 403541 3281 403817 3315
rect 403541 3247 403575 3281
rect 403391 3213 403575 3247
rect 403299 3145 403541 3179
rect 403633 2975 403667 3213
rect 409245 2907 409279 3417
rect 409521 3111 409555 3349
rect 412557 3315 412591 3417
rect 413385 3383 413419 4029
rect 413661 3451 413695 4097
rect 413477 3349 413569 3383
rect 413477 3315 413511 3349
rect 412557 3281 413511 3315
rect 414397 595 414431 3213
rect 416145 2839 416179 4097
rect 419089 3995 419123 4097
rect 418077 3451 418111 3689
rect 418997 3519 419031 3961
rect 421297 3519 421331 3961
rect 423045 3655 423079 3893
rect 416789 3111 416823 3213
rect 418169 2839 418203 3349
rect 418261 3111 418295 3349
rect 418905 2975 418939 3485
rect 422861 3179 422895 3621
rect 425069 3519 425103 4097
rect 432613 3927 432647 3961
rect 432613 3893 432797 3927
rect 447701 3587 447735 3689
rect 427737 2839 427771 3417
rect 509709 3383 509743 3825
rect 523049 3655 523083 3825
rect 540161 2975 540195 3213
<< viali >>
rect 429485 684437 429519 684471
rect 559297 684437 559331 684471
rect 429485 666553 429519 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559297 666553 559331 666587
rect 429209 656829 429243 656863
rect 429209 647241 429243 647275
rect 559205 656829 559239 656863
rect 559205 647241 559239 647275
rect 325801 641665 325835 641699
rect 307125 640237 307159 640271
rect 287161 640101 287195 640135
rect 267841 640033 267875 640067
rect 229661 639829 229695 639863
rect 37381 639557 37415 639591
rect 37473 639557 37507 639591
rect 193229 639557 193263 639591
rect 193413 639557 193447 639591
rect 212641 639557 212675 639591
rect 212733 639557 212767 639591
rect 24777 639489 24811 639523
rect 15209 639421 15243 639455
rect 15209 639285 15243 639319
rect 24777 639285 24811 639319
rect 27629 639489 27663 639523
rect 27629 639285 27663 639319
rect 37197 639489 37231 639523
rect 37197 639285 37231 639319
rect 37289 639489 37323 639523
rect 37289 639285 37323 639319
rect 46949 639489 46983 639523
rect 60657 639489 60691 639523
rect 67649 639489 67683 639523
rect 60841 639421 60875 639455
rect 67649 639353 67683 639387
rect 75929 639489 75963 639523
rect 46949 639285 46983 639319
rect 86969 639489 87003 639523
rect 75929 639285 75963 639319
rect 85497 639421 85531 639455
rect 99297 639489 99331 639523
rect 106289 639489 106323 639523
rect 99481 639421 99515 639455
rect 86969 639353 87003 639387
rect 118617 639489 118651 639523
rect 125609 639489 125643 639523
rect 153209 639489 153243 639523
rect 118801 639421 118835 639455
rect 106289 639353 106323 639387
rect 153577 639421 153611 639455
rect 164249 639489 164283 639523
rect 176577 639489 176611 639523
rect 183569 639489 183603 639523
rect 195897 639489 195931 639523
rect 176761 639421 176795 639455
rect 125609 639353 125643 639387
rect 143549 639353 143583 639387
rect 143641 639353 143675 639387
rect 164249 639353 164283 639387
rect 212549 639489 212583 639523
rect 239321 639829 239355 639863
rect 229753 639761 229787 639795
rect 229753 639557 229787 639591
rect 251833 639829 251867 639863
rect 239321 639557 239355 639591
rect 239413 639761 239447 639795
rect 239413 639557 239447 639591
rect 247601 639761 247635 639795
rect 247601 639557 247635 639591
rect 251833 639557 251867 639591
rect 257905 639829 257939 639863
rect 267749 639829 267783 639863
rect 257905 639557 257939 639591
rect 257997 639761 258031 639795
rect 257997 639557 258031 639591
rect 267749 639557 267783 639591
rect 267841 639557 267875 639591
rect 277225 640033 277259 640067
rect 287069 640033 287103 640067
rect 277225 639557 277259 639591
rect 277317 639829 277351 639863
rect 277317 639557 277351 639591
rect 287069 639557 287103 639591
rect 287161 639557 287195 639591
rect 290565 640101 290599 640135
rect 290565 639557 290599 639591
rect 292589 640033 292623 640067
rect 292589 639557 292623 639591
rect 307033 640033 307067 640067
rect 307033 639557 307067 639591
rect 307125 639557 307159 639591
rect 311817 640237 311851 640271
rect 335185 641665 335219 641699
rect 311817 639557 311851 639591
rect 311909 640033 311943 640067
rect 311909 639557 311943 639591
rect 325801 640033 325835 640067
rect 325801 639557 325835 639591
rect 325893 639557 325927 639591
rect 345029 641665 345063 641699
rect 335185 639557 335219 639591
rect 336013 640033 336047 640067
rect 336013 639557 336047 639591
rect 345029 639557 345063 639591
rect 354597 641665 354631 641699
rect 354597 639557 354631 639591
rect 364349 641665 364383 641699
rect 364349 639557 364383 639591
rect 373917 641665 373951 641699
rect 373917 639557 373951 639591
rect 383669 641665 383703 641699
rect 383669 639557 383703 639591
rect 393237 641665 393271 641699
rect 393237 639557 393271 639591
rect 402989 641665 403023 641699
rect 412557 641665 412591 641699
rect 408325 639625 408359 639659
rect 408509 639625 408543 639659
rect 402989 639557 403023 639591
rect 441721 640645 441755 640679
rect 412557 639557 412591 639591
rect 441629 639693 441663 639727
rect 441629 639557 441663 639591
rect 441721 639557 441755 639591
rect 445217 640645 445251 640679
rect 445217 639557 445251 639591
rect 463709 639693 463743 639727
rect 463709 639557 463743 639591
rect 473277 639693 473311 639727
rect 473277 639557 473311 639591
rect 195989 639421 196023 639455
rect 202889 639421 202923 639455
rect 183569 639353 183603 639387
rect 85497 639285 85531 639319
rect 202889 639285 202923 639319
rect 212457 639421 212491 639455
rect 212641 639421 212675 639455
rect 229661 639421 229695 639455
rect 212457 639285 212491 639319
rect 385049 338113 385083 338147
rect 295625 338045 295659 338079
rect 234629 337705 234663 337739
rect 237481 337705 237515 337739
rect 237481 337569 237515 337603
rect 239413 337637 239447 337671
rect 228097 337501 228131 337535
rect 234997 337501 235031 337535
rect 239413 337501 239447 337535
rect 267473 337501 267507 337535
rect 228281 337365 228315 337399
rect 267473 337365 267507 337399
rect 267565 337501 267599 337535
rect 267565 328457 267599 328491
rect 294061 333897 294095 333931
rect 252661 328389 252695 328423
rect 230673 325533 230707 325567
rect 230673 318801 230707 318835
rect 249993 321657 250027 321691
rect 292773 327029 292807 327063
rect 252661 320093 252695 320127
rect 259653 321589 259687 321623
rect 259653 318801 259687 318835
rect 249993 317441 250027 317475
rect 288633 318733 288667 318767
rect 231961 315945 231995 315979
rect 230673 304249 230707 304283
rect 230673 299489 230707 299523
rect 277593 311865 277627 311899
rect 267105 309145 267139 309179
rect 267105 307785 267139 307819
rect 270693 309077 270727 309111
rect 243001 307717 243035 307751
rect 231961 298129 231995 298163
rect 241805 299421 241839 299455
rect 236285 298061 236319 298095
rect 292773 317441 292807 317475
rect 326353 337909 326387 337943
rect 384313 337909 384347 337943
rect 384221 337773 384255 337807
rect 363245 337705 363279 337739
rect 363337 337705 363371 337739
rect 384313 337569 384347 337603
rect 384405 337705 384439 337739
rect 384405 337501 384439 337535
rect 363337 337433 363371 337467
rect 363429 337433 363463 337467
rect 374561 337433 374595 337467
rect 326353 337161 326387 337195
rect 355977 337297 356011 337331
rect 355977 337093 356011 337127
rect 374561 336753 374595 336787
rect 381461 337433 381495 337467
rect 384221 337433 384255 337467
rect 395445 338113 395479 338147
rect 421021 338045 421055 338079
rect 385049 337297 385083 337331
rect 393881 337909 393915 337943
rect 395445 337909 395479 337943
rect 398757 337909 398791 337943
rect 398757 337297 398791 337331
rect 412925 337433 412959 337467
rect 408509 337229 408543 337263
rect 408509 336957 408543 336991
rect 427553 338045 427587 338079
rect 421021 337161 421055 337195
rect 422953 337841 422987 337875
rect 412925 336889 412959 336923
rect 393881 336821 393915 336855
rect 423045 337433 423079 337467
rect 423045 337229 423079 337263
rect 422953 336821 422987 336855
rect 451473 338045 451507 338079
rect 442181 337841 442215 337875
rect 432153 337569 432187 337603
rect 433441 337501 433475 337535
rect 432153 337365 432187 337399
rect 432613 337365 432647 337399
rect 430497 337161 430531 337195
rect 433349 337297 433383 337331
rect 433441 337297 433475 337331
rect 444021 337841 444055 337875
rect 444021 337501 444055 337535
rect 442181 337297 442215 337331
rect 433349 337161 433383 337195
rect 432613 337093 432647 337127
rect 430497 337025 430531 337059
rect 432889 337025 432923 337059
rect 435833 337025 435867 337059
rect 432521 336957 432555 336991
rect 427553 336821 427587 336855
rect 381461 336753 381495 336787
rect 435833 336753 435867 336787
rect 356529 336685 356563 336719
rect 295625 328457 295659 328491
rect 309425 331245 309459 331279
rect 309425 328457 309459 328491
rect 342637 331245 342671 331279
rect 342637 328457 342671 328491
rect 318993 326145 319027 326179
rect 370053 336685 370087 336719
rect 357633 335257 357667 335291
rect 370053 327097 370087 327131
rect 375573 336685 375607 336719
rect 375573 327097 375607 327131
rect 393145 331245 393179 331279
rect 498945 338045 498979 338079
rect 486341 337773 486375 337807
rect 498945 337637 498979 337671
rect 499773 337637 499807 337671
rect 486341 337365 486375 337399
rect 526729 337569 526763 337603
rect 499773 337297 499807 337331
rect 523601 337501 523635 337535
rect 514033 336957 514067 336991
rect 524061 337433 524095 337467
rect 523693 337161 523727 337195
rect 524061 337161 524095 337195
rect 526729 337161 526763 337195
rect 528661 337161 528695 337195
rect 529857 337161 529891 337195
rect 523693 336957 523727 336991
rect 523601 336821 523635 336855
rect 514033 336753 514067 336787
rect 451473 330497 451507 330531
rect 393145 327097 393179 327131
rect 416881 328389 416915 328423
rect 357633 325805 357667 325839
rect 356529 325669 356563 325703
rect 393237 324173 393271 324207
rect 359013 321589 359047 321623
rect 359013 318801 359047 318835
rect 392133 321589 392167 321623
rect 392133 318801 392167 318835
rect 318993 317441 319027 317475
rect 327273 318733 327307 318767
rect 294061 316013 294095 316047
rect 288633 309145 288667 309179
rect 327273 309145 327307 309179
rect 332793 318733 332827 318767
rect 371341 318733 371375 318767
rect 356529 315945 356563 315979
rect 346593 311797 346627 311831
rect 332793 309145 332827 309179
rect 334449 309145 334483 309179
rect 346593 309145 346627 309179
rect 309333 309077 309367 309111
rect 277593 306357 277627 306391
rect 292773 307717 292807 307751
rect 270693 299489 270727 299523
rect 243001 298129 243035 298163
rect 281641 299421 281675 299455
rect 241805 289833 241839 289867
rect 249901 298061 249935 298095
rect 236285 289697 236319 289731
rect 249901 288405 249935 288439
rect 255513 298061 255547 298095
rect 265265 298061 265299 298095
rect 255513 288405 255547 288439
rect 259653 289765 259687 289799
rect 249901 285821 249935 285855
rect 230857 280109 230891 280143
rect 230857 273241 230891 273275
rect 241805 280109 241839 280143
rect 265265 288405 265299 288439
rect 267013 298061 267047 298095
rect 259653 282761 259687 282795
rect 267013 280177 267047 280211
rect 277593 298061 277627 298095
rect 334449 307785 334483 307819
rect 342453 309009 342487 309043
rect 342453 299557 342487 299591
rect 309333 299489 309367 299523
rect 292773 298197 292807 298231
rect 305193 299421 305227 299455
rect 281641 289833 281675 289867
rect 292681 298061 292715 298095
rect 277593 280177 277627 280211
rect 287253 289765 287287 289799
rect 295717 298061 295751 298095
rect 295717 293233 295751 293267
rect 298385 296633 298419 296667
rect 292681 288405 292715 288439
rect 305193 289833 305227 289867
rect 310713 299421 310747 299455
rect 346593 299421 346627 299455
rect 310713 289833 310747 289867
rect 324513 299353 324547 299387
rect 324513 289833 324547 289867
rect 331413 298061 331447 298095
rect 298385 287045 298419 287079
rect 309333 289697 309367 289731
rect 287253 280177 287287 280211
rect 331413 288405 331447 288439
rect 334265 298061 334299 298095
rect 376861 318733 376895 318767
rect 371341 309281 371375 309315
rect 375757 317373 375791 317407
rect 376861 309281 376895 309315
rect 381277 317373 381311 317407
rect 375757 309077 375791 309111
rect 376861 309077 376895 309111
rect 381277 307785 381311 307819
rect 382289 317373 382323 317407
rect 387901 317373 387935 317407
rect 416881 318801 416915 318835
rect 422401 328389 422435 328423
rect 422401 318801 422435 318835
rect 427921 328389 427955 328423
rect 427921 318801 427955 318835
rect 433717 328389 433751 328423
rect 472081 328389 472115 328423
rect 433717 318801 433751 318835
rect 466561 321589 466595 321623
rect 466561 318801 466595 318835
rect 472081 318801 472115 318835
rect 397745 318733 397779 318767
rect 397745 312137 397779 312171
rect 451565 315945 451599 315979
rect 393237 309145 393271 309179
rect 387901 307785 387935 307819
rect 416881 309077 416915 309111
rect 382289 302073 382323 302107
rect 387901 304861 387935 304895
rect 376861 299489 376895 299523
rect 356529 298129 356563 298163
rect 382473 299421 382507 299455
rect 346593 289833 346627 289867
rect 353493 298061 353527 298095
rect 370145 298061 370179 298095
rect 387901 298129 387935 298163
rect 408785 302209 408819 302243
rect 422493 309077 422527 309111
rect 422493 299897 422527 299931
rect 428013 309077 428047 309111
rect 416881 299489 416915 299523
rect 428013 299489 428047 299523
rect 433441 309077 433475 309111
rect 451565 302073 451599 302107
rect 466561 309077 466595 309111
rect 433441 299489 433475 299523
rect 466561 299489 466595 299523
rect 472081 309077 472115 309111
rect 472081 299489 472115 299523
rect 408785 298129 408819 298163
rect 382473 289833 382507 289867
rect 408785 293029 408819 293063
rect 370145 289697 370179 289731
rect 353493 288405 353527 288439
rect 334265 282761 334299 282795
rect 342545 282897 342579 282931
rect 408785 282761 408819 282795
rect 342545 280245 342579 280279
rect 309333 280177 309367 280211
rect 249901 278749 249935 278783
rect 283113 280109 283147 280143
rect 241805 270521 241839 270555
rect 270601 278681 270635 278715
rect 252753 270453 252787 270487
rect 231869 263585 231903 263619
rect 270601 269093 270635 269127
rect 277685 275077 277719 275111
rect 305193 280109 305227 280143
rect 283113 270521 283147 270555
rect 295441 278681 295475 278715
rect 277685 269093 277719 269127
rect 287253 270453 287287 270487
rect 252753 260865 252787 260899
rect 267013 263585 267047 263619
rect 231869 259437 231903 259471
rect 241805 260797 241839 260831
rect 230949 254405 230983 254439
rect 305193 270521 305227 270555
rect 310713 280109 310747 280143
rect 327273 280109 327307 280143
rect 327273 272153 327307 272187
rect 334357 280109 334391 280143
rect 334357 270589 334391 270623
rect 346593 280109 346627 280143
rect 310713 270521 310747 270555
rect 364533 280109 364567 280143
rect 364533 273173 364567 273207
rect 371433 280109 371467 280143
rect 346593 270521 346627 270555
rect 376953 280109 376987 280143
rect 371433 270521 371467 270555
rect 375481 278681 375515 278715
rect 295441 269093 295475 269127
rect 309333 270385 309367 270419
rect 287253 260865 287287 260899
rect 309333 260865 309367 260899
rect 324421 263585 324455 263619
rect 324421 260865 324455 260899
rect 342545 263585 342579 263619
rect 376953 270521 376987 270555
rect 393237 280109 393271 280143
rect 393237 270521 393271 270555
rect 400505 280109 400539 280143
rect 416881 280109 416915 280143
rect 400505 270521 400539 270555
rect 408785 278681 408819 278715
rect 392133 270453 392167 270487
rect 375481 263449 375515 263483
rect 381093 270385 381127 270419
rect 342545 260865 342579 260899
rect 392133 264265 392167 264299
rect 416881 270521 416915 270555
rect 433625 280109 433659 280143
rect 466561 280109 466595 280143
rect 433625 270521 433659 270555
rect 451565 273717 451599 273751
rect 408785 263449 408819 263483
rect 466561 270521 466595 270555
rect 472081 280109 472115 280143
rect 472081 270521 472115 270555
rect 451565 263449 451599 263483
rect 381093 260865 381127 260899
rect 267013 259437 267047 259471
rect 283113 260797 283147 260831
rect 241805 251209 241839 251243
rect 281917 259369 281951 259403
rect 252753 251141 252787 251175
rect 230949 244137 230983 244171
rect 236285 244273 236319 244307
rect 305193 260797 305227 260831
rect 295441 259369 295475 259403
rect 283113 251209 283147 251243
rect 292957 258009 292991 258043
rect 281917 241553 281951 241587
rect 287253 251141 287287 251175
rect 252753 241485 252787 241519
rect 292957 249713 292991 249747
rect 287253 241485 287287 241519
rect 236285 240193 236319 240227
rect 281917 241417 281951 241451
rect 236285 240057 236319 240091
rect 310713 260797 310747 260831
rect 305193 251209 305227 251243
rect 309333 260729 309367 260763
rect 309333 251209 309367 251243
rect 310713 251209 310747 251243
rect 327273 260797 327307 260831
rect 334357 260797 334391 260831
rect 346593 260797 346627 260831
rect 334357 251277 334391 251311
rect 342453 260729 342487 260763
rect 327273 251209 327307 251243
rect 342453 251209 342487 251243
rect 359013 260797 359047 260831
rect 346593 251209 346627 251243
rect 348065 254609 348099 254643
rect 298201 251141 298235 251175
rect 334357 251141 334391 251175
rect 334357 244137 334391 244171
rect 298201 242641 298235 242675
rect 348065 241485 348099 241519
rect 353585 254609 353619 254643
rect 356437 253997 356471 254031
rect 359013 251277 359047 251311
rect 371433 260797 371467 260831
rect 371433 251209 371467 251243
rect 375573 260797 375607 260831
rect 375573 251209 375607 251243
rect 376953 260797 376987 260831
rect 376953 251209 376987 251243
rect 400505 260797 400539 260831
rect 400505 251209 400539 251243
rect 416881 260797 416915 260831
rect 416881 251209 416915 251243
rect 433625 260797 433659 260831
rect 466561 260797 466595 260831
rect 433625 251209 433659 251243
rect 451565 259369 451599 259403
rect 356437 251073 356471 251107
rect 359013 251141 359047 251175
rect 359013 244137 359047 244171
rect 369961 251141 369995 251175
rect 353585 241485 353619 241519
rect 369961 241485 369995 241519
rect 381093 251073 381127 251107
rect 466561 251209 466595 251243
rect 472081 260797 472115 260831
rect 472081 251209 472115 251243
rect 451565 244137 451599 244171
rect 381093 241485 381127 241519
rect 295441 240057 295475 240091
rect 348065 238697 348099 238731
rect 281917 234549 281951 234583
rect 295533 237337 295567 237371
rect 259653 231761 259687 231795
rect 236285 230537 236319 230571
rect 243185 231693 243219 231727
rect 243185 224213 243219 224247
rect 392133 236725 392167 236759
rect 364441 235909 364475 235943
rect 356437 234685 356471 234719
rect 348065 230333 348099 230367
rect 352021 234617 352055 234651
rect 352021 230333 352055 230367
rect 356437 229177 356471 229211
rect 295533 227749 295567 227783
rect 356437 229041 356471 229075
rect 259653 222173 259687 222207
rect 267105 224961 267139 224995
rect 324421 224961 324455 224995
rect 356437 224893 356471 224927
rect 324421 222241 324455 222275
rect 267105 220813 267139 220847
rect 281917 222173 281951 222207
rect 281917 220813 281951 220847
rect 324421 222105 324455 222139
rect 324421 219521 324455 219555
rect 267013 219385 267047 219419
rect 243093 217957 243127 217991
rect 236285 205581 236319 205615
rect 236285 202861 236319 202895
rect 381093 234685 381127 234719
rect 381093 231829 381127 231863
rect 381185 224961 381219 224995
rect 381185 222173 381219 222207
rect 392133 222173 392167 222207
rect 408693 231761 408727 231795
rect 408693 222173 408727 222207
rect 364441 218025 364475 218059
rect 298293 215441 298327 215475
rect 295441 215373 295475 215407
rect 381093 215373 381127 215407
rect 309333 215305 309367 215339
rect 309333 212517 309367 212551
rect 358921 212585 358955 212619
rect 298293 211225 298327 211259
rect 267013 209797 267047 209831
rect 281733 211089 281767 211123
rect 295441 211089 295475 211123
rect 298293 211089 298327 211123
rect 265173 209729 265207 209763
rect 265173 202793 265207 202827
rect 356437 211089 356471 211123
rect 298293 205581 298327 205615
rect 309425 205649 309459 205683
rect 309425 202861 309459 202895
rect 324421 205649 324455 205683
rect 324421 202861 324455 202895
rect 331413 202929 331447 202963
rect 281733 202793 281767 202827
rect 381093 212517 381127 212551
rect 397653 215305 397687 215339
rect 397653 212517 397687 212551
rect 358921 208369 358955 208403
rect 408693 212449 408727 212483
rect 408693 202861 408727 202895
rect 356437 202793 356471 202827
rect 331413 201501 331447 201535
rect 243093 201433 243127 201467
rect 236285 198645 236319 198679
rect 292773 198645 292807 198679
rect 270785 196061 270819 196095
rect 270785 193137 270819 193171
rect 236285 189057 236319 189091
rect 266461 191777 266495 191811
rect 266461 183345 266495 183379
rect 252845 182121 252879 182155
rect 232145 180761 232179 180795
rect 232145 162877 232179 162911
rect 236377 179333 236411 179367
rect 324421 196061 324455 196095
rect 309333 195993 309367 196027
rect 298293 193205 298327 193239
rect 309333 193205 309367 193239
rect 298293 191845 298327 191879
rect 397653 195993 397687 196027
rect 397653 193205 397687 193239
rect 324421 191845 324455 191879
rect 295625 188445 295659 188479
rect 295625 183549 295659 183583
rect 298385 186473 298419 186507
rect 298385 183549 298419 183583
rect 334449 186405 334483 186439
rect 334449 183549 334483 183583
rect 357541 186405 357575 186439
rect 357541 183549 357575 183583
rect 292773 180829 292807 180863
rect 451657 183481 451691 183515
rect 386613 180761 386647 180795
rect 252845 172533 252879 172567
rect 254133 177293 254167 177327
rect 254133 172533 254167 172567
rect 334357 175865 334391 175899
rect 298293 172465 298327 172499
rect 236377 161449 236411 161483
rect 243093 171037 243127 171071
rect 295533 171037 295567 171071
rect 243093 161449 243127 161483
rect 259653 164169 259687 164203
rect 232145 161381 232179 161415
rect 283113 164169 283147 164203
rect 259653 154581 259687 154615
rect 265265 161381 265299 161415
rect 232145 151793 232179 151827
rect 267013 157437 267047 157471
rect 283113 154921 283147 154955
rect 288633 164169 288667 164203
rect 298293 166957 298327 166991
rect 309333 172465 309367 172499
rect 309333 164169 309367 164203
rect 324513 171037 324547 171071
rect 295533 161449 295567 161483
rect 386613 171105 386647 171139
rect 392133 180761 392167 180795
rect 427921 176681 427955 176715
rect 427921 173893 427955 173927
rect 433625 176613 433659 176647
rect 433625 173893 433659 173927
rect 451657 173893 451691 173927
rect 392133 171105 392167 171139
rect 334357 169745 334391 169779
rect 364533 167637 364567 167671
rect 324513 161449 324547 161483
rect 347973 164169 348007 164203
rect 331413 161381 331447 161415
rect 288633 154921 288667 154955
rect 294061 158661 294095 158695
rect 267013 153153 267047 153187
rect 270693 154513 270727 154547
rect 265265 151793 265299 151827
rect 270693 147577 270727 147611
rect 292773 151725 292807 151759
rect 321753 153153 321787 153187
rect 294061 149073 294095 149107
rect 295625 150365 295659 150399
rect 292773 142137 292807 142171
rect 231961 142069 231995 142103
rect 236469 142069 236503 142103
rect 236469 132481 236503 132515
rect 240149 142069 240183 142103
rect 266461 142069 266495 142103
rect 240149 132481 240183 132515
rect 243093 133841 243127 133875
rect 231961 124185 231995 124219
rect 357633 164169 357667 164203
rect 347973 155737 348007 155771
rect 352021 162809 352055 162843
rect 352021 154513 352055 154547
rect 353493 162809 353527 162843
rect 353493 153221 353527 153255
rect 356437 162809 356471 162843
rect 357633 154581 357667 154615
rect 359013 157301 359047 157335
rect 359013 154581 359047 154615
rect 422401 164169 422435 164203
rect 364533 154581 364567 154615
rect 381001 162809 381035 162843
rect 356437 153221 356471 153255
rect 370053 154513 370087 154547
rect 331413 151793 331447 151827
rect 347973 153153 348007 153187
rect 321753 143565 321787 143599
rect 324605 151725 324639 151759
rect 324605 142137 324639 142171
rect 334357 144857 334391 144891
rect 295625 140777 295659 140811
rect 294061 139349 294095 139383
rect 266461 132481 266495 132515
rect 270693 135201 270727 135235
rect 265357 132413 265391 132447
rect 281641 135201 281675 135235
rect 281641 129013 281675 129047
rect 270693 128265 270727 128299
rect 265357 124593 265391 124627
rect 283113 125545 283147 125579
rect 243093 124185 243127 124219
rect 236377 122757 236411 122791
rect 327181 135269 327215 135303
rect 298385 133773 298419 133807
rect 294061 121465 294095 121499
rect 295533 131053 295567 131087
rect 347973 144789 348007 144823
rect 353493 153085 353527 153119
rect 370053 147577 370087 147611
rect 387993 162809 388027 162843
rect 387993 157981 388027 158015
rect 422401 157301 422435 157335
rect 427921 164169 427955 164203
rect 427921 157301 427955 157335
rect 408693 154513 408727 154547
rect 400505 153153 400539 153187
rect 381001 147577 381035 147611
rect 392133 148325 392167 148359
rect 353493 144789 353527 144823
rect 400505 147577 400539 147611
rect 408693 147577 408727 147611
rect 451657 154513 451691 154547
rect 451657 147577 451691 147611
rect 466561 154445 466595 154479
rect 466561 147577 466595 147611
rect 392133 135269 392167 135303
rect 393237 144857 393271 144891
rect 422401 144857 422435 144891
rect 397745 143497 397779 143531
rect 397745 137921 397779 137955
rect 472081 143497 472115 143531
rect 422401 137921 422435 137955
rect 427921 138057 427955 138091
rect 393237 135269 393271 135303
rect 427921 135269 427955 135303
rect 334357 135133 334391 135167
rect 370053 135201 370087 135235
rect 327181 132481 327215 132515
rect 298385 124185 298419 124219
rect 309333 132413 309367 132447
rect 321753 132413 321787 132447
rect 309333 122825 309367 122859
rect 310713 125545 310747 125579
rect 295533 121465 295567 121499
rect 294153 121329 294187 121363
rect 305193 120717 305227 120751
rect 294153 116569 294187 116603
rect 298385 119357 298419 119391
rect 283113 115957 283147 115991
rect 236377 113169 236411 113203
rect 254133 115889 254167 115923
rect 305193 115957 305227 115991
rect 321753 122825 321787 122859
rect 324421 132413 324455 132447
rect 370053 128265 370087 128299
rect 408693 135201 408727 135235
rect 408693 128265 408727 128299
rect 472081 128265 472115 128299
rect 324421 122825 324455 122859
rect 346593 125545 346627 125579
rect 310713 115957 310747 115991
rect 318993 118745 319027 118779
rect 298385 114529 298419 114563
rect 254133 108953 254167 108987
rect 267013 114461 267047 114495
rect 243185 106165 243219 106199
rect 232145 104805 232179 104839
rect 230857 96577 230891 96611
rect 243185 96713 243219 96747
rect 252753 106165 252787 106199
rect 298201 114393 298235 114427
rect 292773 113101 292807 113135
rect 267013 104941 267047 104975
rect 283113 106233 283147 106267
rect 252753 96645 252787 96679
rect 267013 104805 267047 104839
rect 232145 95217 232179 95251
rect 267013 95217 267047 95251
rect 270877 102085 270911 102119
rect 230857 89641 230891 89675
rect 265173 95149 265207 95183
rect 241805 86921 241839 86955
rect 231961 85493 231995 85527
rect 230949 80121 230983 80155
rect 230949 77265 230983 77299
rect 231961 75905 231995 75939
rect 236285 85493 236319 85527
rect 241805 77265 241839 77299
rect 252753 86853 252787 86887
rect 252753 77265 252787 77299
rect 254133 86853 254167 86887
rect 254133 77265 254167 77299
rect 259653 86853 259687 86887
rect 292773 103581 292807 103615
rect 295625 111741 295659 111775
rect 283113 96645 283147 96679
rect 292681 103445 292715 103479
rect 298201 104873 298235 104907
rect 305193 106233 305227 106267
rect 295625 102153 295659 102187
rect 298385 99433 298419 99467
rect 305193 96645 305227 96679
rect 310713 106233 310747 106267
rect 364533 125545 364567 125579
rect 346593 115957 346627 115991
rect 353585 115957 353619 115991
rect 364533 115957 364567 115991
rect 376953 125545 376987 125579
rect 376953 115957 376987 115991
rect 393237 125545 393271 125579
rect 422401 125545 422435 125579
rect 393237 115957 393271 115991
rect 400321 124117 400355 124151
rect 342453 115889 342487 115923
rect 334357 114529 334391 114563
rect 318993 104873 319027 104907
rect 327181 114461 327215 114495
rect 334357 113169 334391 113203
rect 353585 114529 353619 114563
rect 422401 118609 422435 118643
rect 427921 125545 427955 125579
rect 427921 118609 427955 118643
rect 433625 125545 433659 125579
rect 433625 118609 433659 118643
rect 451473 124117 451507 124151
rect 400321 114529 400355 114563
rect 451473 114529 451507 114563
rect 466653 124117 466687 124151
rect 466653 114529 466687 114563
rect 342453 108953 342487 108987
rect 356437 114461 356471 114495
rect 327181 104873 327215 104907
rect 346593 106233 346627 106267
rect 310713 96645 310747 96679
rect 334357 103445 334391 103479
rect 298385 95217 298419 95251
rect 292681 93857 292715 93891
rect 324513 95149 324547 95183
rect 270877 92497 270911 92531
rect 265173 85561 265207 85595
rect 298385 89709 298419 89743
rect 298385 85561 298419 85595
rect 305193 86921 305227 86955
rect 259653 77265 259687 77299
rect 270693 82773 270727 82807
rect 236285 75905 236319 75939
rect 230949 75837 230983 75871
rect 236285 70329 236319 70363
rect 236285 67609 236319 67643
rect 230949 66249 230983 66283
rect 236377 66181 236411 66215
rect 298293 80733 298327 80767
rect 277409 77197 277443 77231
rect 270693 64889 270727 64923
rect 271981 73117 272015 73151
rect 243001 64821 243035 64855
rect 260849 64821 260883 64855
rect 259653 59721 259687 59755
rect 243001 55233 243035 55267
rect 244381 56525 244415 56559
rect 236377 47005 236411 47039
rect 244381 46937 244415 46971
rect 249993 56525 250027 56559
rect 249993 46937 250027 46971
rect 255421 56525 255455 56559
rect 277409 70329 277443 70363
rect 305193 77265 305227 77299
rect 308045 86921 308079 86955
rect 308045 77265 308079 77299
rect 309333 86921 309367 86955
rect 309333 77265 309367 77299
rect 310713 86921 310747 86955
rect 324513 85561 324547 85595
rect 327273 95149 327307 95183
rect 387993 114461 388027 114495
rect 370145 109021 370179 109055
rect 370145 106301 370179 106335
rect 356437 104941 356471 104975
rect 376953 106233 376987 106267
rect 346593 96645 346627 96679
rect 353493 104805 353527 104839
rect 353493 95217 353527 95251
rect 356437 104805 356471 104839
rect 387993 104873 388027 104907
rect 422401 106233 422435 106267
rect 376953 96645 376987 96679
rect 408693 104805 408727 104839
rect 356437 95217 356471 95251
rect 422401 99297 422435 99331
rect 427921 106233 427955 106267
rect 427921 99297 427955 99331
rect 451565 104805 451599 104839
rect 408693 95217 408727 95251
rect 451565 95217 451599 95251
rect 334357 93857 334391 93891
rect 387993 95149 388027 95183
rect 342453 86921 342487 86955
rect 327273 85561 327307 85595
rect 331413 86853 331447 86887
rect 310713 77265 310747 77299
rect 331413 77265 331447 77299
rect 334357 86853 334391 86887
rect 334357 77265 334391 77299
rect 346593 86921 346627 86955
rect 364533 86853 364567 86887
rect 346593 80733 346627 80767
rect 359013 82773 359047 82807
rect 342453 77265 342487 77299
rect 327181 75837 327215 75871
rect 298293 67609 298327 67643
rect 319085 67609 319119 67643
rect 308045 67541 308079 67575
rect 271981 63529 272015 63563
rect 281733 66181 281767 66215
rect 271981 58565 272015 58599
rect 260849 55233 260883 55267
rect 270601 57545 270635 57579
rect 259653 48297 259687 48331
rect 255421 46937 255455 46971
rect 270601 46937 270635 46971
rect 319085 66249 319119 66283
rect 353585 75837 353619 75871
rect 357541 74477 357575 74511
rect 327181 66249 327215 66283
rect 330033 66249 330067 66283
rect 353585 66249 353619 66283
rect 356437 67541 356471 67575
rect 308045 57953 308079 57987
rect 309425 66045 309459 66079
rect 281733 56593 281767 56627
rect 288541 57885 288575 57919
rect 282929 56525 282963 56559
rect 298293 56525 298327 56559
rect 288541 48297 288575 48331
rect 292773 55165 292807 55199
rect 282929 47005 282963 47039
rect 271981 45577 272015 45611
rect 330033 64957 330067 64991
rect 329941 63461 329975 63495
rect 309425 48365 309459 48399
rect 318993 59993 319027 60027
rect 298293 46937 298327 46971
rect 308137 48229 308171 48263
rect 292773 45577 292807 45611
rect 243001 45509 243035 45543
rect 267013 45509 267047 45543
rect 255513 44829 255547 44863
rect 243001 35921 243035 35955
rect 252753 37349 252787 37383
rect 252753 28985 252787 29019
rect 277593 45509 277627 45543
rect 272073 38709 272107 38743
rect 272073 37213 272107 37247
rect 267013 35921 267047 35955
rect 277593 35921 277627 35955
rect 282929 45509 282963 45543
rect 298385 42041 298419 42075
rect 294153 38573 294187 38607
rect 292773 37145 292807 37179
rect 292773 35921 292807 35955
rect 324421 57885 324455 57919
rect 324421 55301 324455 55335
rect 318993 46937 319027 46971
rect 324513 55165 324547 55199
rect 310529 46869 310563 46903
rect 308137 38641 308171 38675
rect 309333 42041 309367 42075
rect 298385 32385 298419 32419
rect 294153 29053 294187 29087
rect 332885 63461 332919 63495
rect 329941 53805 329975 53839
rect 331413 55641 331447 55675
rect 352021 58089 352055 58123
rect 336933 56525 336967 56559
rect 332885 55165 332919 55199
rect 334357 55641 334391 55675
rect 331413 48297 331447 48331
rect 334357 48297 334391 48331
rect 364533 77265 364567 77299
rect 370053 86853 370087 86887
rect 370053 77265 370087 77299
rect 386613 86853 386647 86887
rect 393237 95149 393271 95183
rect 387993 85561 388027 85595
rect 392133 86853 392167 86887
rect 386613 77265 386647 77299
rect 393237 85561 393271 85595
rect 397653 86921 397687 86955
rect 392133 77265 392167 77299
rect 397653 77265 397687 77299
rect 400321 86921 400355 86955
rect 422401 86921 422435 86955
rect 400321 77265 400355 77299
rect 408785 82093 408819 82127
rect 408785 77265 408819 77299
rect 422401 77265 422435 77299
rect 427921 86921 427955 86955
rect 427921 77265 427955 77299
rect 433441 86921 433475 86955
rect 433441 77265 433475 77299
rect 451473 85493 451507 85527
rect 359013 73185 359047 73219
rect 416881 77197 416915 77231
rect 408785 70397 408819 70431
rect 408785 67609 408819 67643
rect 416881 67609 416915 67643
rect 466561 85493 466595 85527
rect 466561 75905 466595 75939
rect 472081 80733 472115 80767
rect 451473 67609 451507 67643
rect 472081 67609 472115 67643
rect 393237 67541 393271 67575
rect 357541 64889 357575 64923
rect 387993 66181 388027 66215
rect 356437 57953 356471 57987
rect 359105 63461 359139 63495
rect 352021 53805 352055 53839
rect 359105 53805 359139 53839
rect 370053 61081 370087 61115
rect 375573 61081 375607 61115
rect 371433 60605 371467 60639
rect 371433 56661 371467 56695
rect 370053 48297 370087 48331
rect 371433 56525 371467 56559
rect 375573 48297 375607 48331
rect 382381 57885 382415 57919
rect 393237 57953 393271 57987
rect 397653 67541 397687 67575
rect 451473 66181 451507 66215
rect 397653 57953 397687 57987
rect 408785 62781 408819 62815
rect 451473 60673 451507 60707
rect 466469 66181 466503 66215
rect 408785 57953 408819 57987
rect 387993 56593 388027 56627
rect 416881 57885 416915 57919
rect 382381 48297 382415 48331
rect 392133 56525 392167 56559
rect 371433 47005 371467 47039
rect 400413 51153 400447 51187
rect 400413 48365 400447 48399
rect 408785 51153 408819 51187
rect 408785 48365 408819 48399
rect 416881 48365 416915 48399
rect 433625 57885 433659 57919
rect 466469 56593 466503 56627
rect 472081 57885 472115 57919
rect 433625 48297 433659 48331
rect 451657 56525 451691 56559
rect 392133 47005 392167 47039
rect 336933 46937 336967 46971
rect 472081 48297 472115 48331
rect 451657 46937 451691 46971
rect 324513 45577 324547 45611
rect 342453 46869 342487 46903
rect 310529 41361 310563 41395
rect 332701 45509 332735 45543
rect 387901 46869 387935 46903
rect 342453 37281 342487 37315
rect 359013 45509 359047 45543
rect 332701 35921 332735 35955
rect 375481 41565 375515 41599
rect 369961 41429 369995 41463
rect 369961 38573 369995 38607
rect 375481 37281 375515 37315
rect 408785 46869 408819 46903
rect 433625 41293 433659 41327
rect 408785 38505 408819 38539
rect 416881 38573 416915 38607
rect 387901 37281 387935 37315
rect 359013 35921 359047 35955
rect 309333 28985 309367 29019
rect 334357 35853 334391 35887
rect 282929 27625 282963 27659
rect 308045 28917 308079 28951
rect 252845 27557 252879 27591
rect 255513 27557 255547 27591
rect 259837 27557 259871 27591
rect 230673 26197 230707 26231
rect 252845 17969 252879 18003
rect 271981 27557 272015 27591
rect 259837 17969 259871 18003
rect 270693 22593 270727 22627
rect 293969 27557 294003 27591
rect 271981 17969 272015 18003
rect 277501 26197 277535 26231
rect 305101 22185 305135 22219
rect 305101 19329 305135 19363
rect 308045 19329 308079 19363
rect 321661 27557 321695 27591
rect 293969 17969 294003 18003
rect 400689 31773 400723 31807
rect 400689 29053 400723 29087
rect 416881 28985 416915 29019
rect 422493 38573 422527 38607
rect 393237 28917 393271 28951
rect 387809 27761 387843 27795
rect 387809 27625 387843 27659
rect 334357 26265 334391 26299
rect 336841 27557 336875 27591
rect 321661 17969 321695 18003
rect 346409 27557 346443 27591
rect 353677 27557 353711 27591
rect 346409 22729 346443 22763
rect 347881 22729 347915 22763
rect 336841 17969 336875 18003
rect 277501 16609 277535 16643
rect 270693 14705 270727 14739
rect 260941 12529 260975 12563
rect 232789 12461 232823 12495
rect 232789 11713 232823 11747
rect 293969 12461 294003 12495
rect 353677 19261 353711 19295
rect 359013 27557 359047 27591
rect 433625 37349 433659 37383
rect 472081 38573 472115 38607
rect 422493 27625 422527 27659
rect 433625 37213 433659 37247
rect 472081 28985 472115 29019
rect 433625 27625 433659 27659
rect 451749 28917 451783 28951
rect 393237 19329 393271 19363
rect 400597 27557 400631 27591
rect 359013 17969 359047 18003
rect 451749 19329 451783 19363
rect 400597 17969 400631 18003
rect 416973 19261 417007 19295
rect 347881 12393 347915 12427
rect 381001 17901 381035 17935
rect 293969 11849 294003 11883
rect 260941 11713 260975 11747
rect 346501 9605 346535 9639
rect 346501 8449 346535 8483
rect 230673 8313 230707 8347
rect 381001 8313 381035 8347
rect 382381 17901 382415 17935
rect 400413 17833 400447 17867
rect 382381 8313 382415 8347
rect 393053 9605 393087 9639
rect 315221 6749 315255 6783
rect 315221 5865 315255 5899
rect 322213 6001 322247 6035
rect 322213 5797 322247 5831
rect 280169 4097 280203 4131
rect 277961 3961 277995 3995
rect 278053 3961 278087 3995
rect 278053 3689 278087 3723
rect 278145 3689 278179 3723
rect 238217 3621 238251 3655
rect 238217 3485 238251 3519
rect 278053 3553 278087 3587
rect 278053 3349 278087 3383
rect 391213 4097 391247 4131
rect 384313 3961 384347 3995
rect 391213 3893 391247 3927
rect 392961 4029 392995 4063
rect 392961 3825 392995 3859
rect 374653 3689 374687 3723
rect 384313 3689 384347 3723
rect 280169 3281 280203 3315
rect 292589 3553 292623 3587
rect 292589 3281 292623 3315
rect 302157 3485 302191 3519
rect 374653 3417 374687 3451
rect 374745 3417 374779 3451
rect 302157 3281 302191 3315
rect 335185 3281 335219 3315
rect 82921 3145 82955 3179
rect 335185 3145 335219 3179
rect 363245 3281 363279 3315
rect 363245 3077 363279 3111
rect 369869 3145 369903 3179
rect 82921 2941 82955 2975
rect 98653 2941 98687 2975
rect 374745 2941 374779 2975
rect 121469 2873 121503 2907
rect 121653 2873 121687 2907
rect 369869 2873 369903 2907
rect 98653 2805 98687 2839
rect 416973 12257 417007 12291
rect 400413 8313 400447 8347
rect 403265 4301 403299 4335
rect 393881 4097 393915 4131
rect 393973 4029 394007 4063
rect 400045 4029 400079 4063
rect 400045 3825 400079 3859
rect 408417 4301 408451 4335
rect 408233 4233 408267 4267
rect 403357 4165 403391 4199
rect 403357 3825 403391 3859
rect 403725 3961 403759 3995
rect 403265 3689 403299 3723
rect 393973 3349 394007 3383
rect 402437 3417 402471 3451
rect 393881 3213 393915 3247
rect 408325 4165 408359 4199
rect 408325 3961 408359 3995
rect 413661 4097 413695 4131
rect 408509 4029 408543 4063
rect 409245 4029 409279 4063
rect 413385 4029 413419 4063
rect 408417 3961 408451 3995
rect 403725 3689 403759 3723
rect 408233 3689 408267 3723
rect 403541 3417 403575 3451
rect 408417 3621 408451 3655
rect 408417 3417 408451 3451
rect 409889 3417 409923 3451
rect 412557 3417 412591 3451
rect 403449 3281 403483 3315
rect 403817 3281 403851 3315
rect 402437 3213 402471 3247
rect 403357 3213 403391 3247
rect 403633 3213 403667 3247
rect 403265 3145 403299 3179
rect 403541 3145 403575 3179
rect 403633 2941 403667 2975
rect 409521 3349 409555 3383
rect 413661 3417 413695 3451
rect 416145 4097 416179 4131
rect 413385 3349 413419 3383
rect 413569 3349 413603 3383
rect 409521 3077 409555 3111
rect 414397 3213 414431 3247
rect 409245 2873 409279 2907
rect 393053 561 393087 595
rect 419089 4097 419123 4131
rect 425069 4097 425103 4131
rect 418997 3961 419031 3995
rect 419089 3961 419123 3995
rect 421297 3961 421331 3995
rect 418077 3689 418111 3723
rect 418077 3417 418111 3451
rect 418905 3485 418939 3519
rect 418997 3485 419031 3519
rect 423045 3893 423079 3927
rect 421297 3485 421331 3519
rect 422861 3621 422895 3655
rect 423045 3621 423079 3655
rect 418169 3349 418203 3383
rect 416789 3213 416823 3247
rect 416789 3077 416823 3111
rect 416145 2805 416179 2839
rect 418261 3349 418295 3383
rect 418261 3077 418295 3111
rect 432613 3961 432647 3995
rect 432797 3893 432831 3927
rect 509709 3825 509743 3859
rect 447701 3689 447735 3723
rect 447701 3553 447735 3587
rect 425069 3485 425103 3519
rect 422861 3145 422895 3179
rect 427737 3417 427771 3451
rect 418905 2941 418939 2975
rect 418169 2805 418203 2839
rect 523049 3825 523083 3859
rect 523049 3621 523083 3655
rect 509709 3349 509743 3383
rect 540161 3213 540195 3247
rect 540161 2941 540195 2975
rect 427737 2805 427771 2839
rect 414397 561 414431 595
<< metal1 >>
rect 218974 700952 218980 701004
rect 219032 700992 219038 701004
rect 393314 700992 393320 701004
rect 219032 700964 393320 700992
rect 219032 700952 219038 700964
rect 393314 700952 393320 700964
rect 393372 700952 393378 701004
rect 355962 700884 355968 700936
rect 356020 700924 356026 700936
rect 543458 700924 543464 700936
rect 356020 700896 543464 700924
rect 356020 700884 356026 700896
rect 543458 700884 543464 700896
rect 543516 700884 543522 700936
rect 202782 700816 202788 700868
rect 202840 700856 202846 700868
rect 390554 700856 390560 700868
rect 202840 700828 390560 700856
rect 202840 700816 202846 700828
rect 390554 700816 390560 700828
rect 390612 700816 390618 700868
rect 170306 700748 170312 700800
rect 170364 700788 170370 700800
rect 396074 700788 396080 700800
rect 170364 700760 396080 700788
rect 170364 700748 170370 700760
rect 396074 700748 396080 700760
rect 396132 700748 396138 700800
rect 154114 700680 154120 700732
rect 154172 700720 154178 700732
rect 401594 700720 401600 700732
rect 154172 700692 401600 700720
rect 154172 700680 154178 700692
rect 401594 700680 401600 700692
rect 401652 700680 401658 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 398834 700652 398840 700664
rect 137888 700624 398840 700652
rect 137888 700612 137894 700624
rect 398834 700612 398840 700624
rect 398892 700612 398898 700664
rect 105446 700544 105452 700596
rect 105504 700584 105510 700596
rect 404354 700584 404360 700596
rect 105504 700556 404360 700584
rect 105504 700544 105510 700556
rect 404354 700544 404360 700556
rect 404412 700544 404418 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 409874 700516 409880 700528
rect 89220 700488 409880 700516
rect 89220 700476 89226 700488
rect 409874 700476 409880 700488
rect 409932 700476 409938 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 407114 700448 407120 700460
rect 73028 700420 407120 700448
rect 73028 700408 73034 700420
rect 407114 700408 407120 700420
rect 407172 700408 407178 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 411254 700380 411260 700392
rect 40552 700352 411260 700380
rect 40552 700340 40558 700352
rect 411254 700340 411260 700352
rect 411312 700340 411318 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 416774 700312 416780 700324
rect 24360 700284 416780 700312
rect 24360 700272 24366 700284
rect 416774 700272 416780 700284
rect 416832 700272 416838 700324
rect 353202 700204 353208 700256
rect 353260 700244 353266 700256
rect 527174 700244 527180 700256
rect 353260 700216 527180 700244
rect 353260 700204 353266 700216
rect 527174 700204 527180 700216
rect 527232 700204 527238 700256
rect 267642 700136 267648 700188
rect 267700 700176 267706 700188
rect 383654 700176 383660 700188
rect 267700 700148 383660 700176
rect 267700 700136 267706 700148
rect 383654 700136 383660 700148
rect 383712 700136 383718 700188
rect 362862 700068 362868 700120
rect 362920 700108 362926 700120
rect 478506 700108 478512 700120
rect 362920 700080 478512 700108
rect 362920 700068 362926 700080
rect 478506 700068 478512 700080
rect 478564 700068 478570 700120
rect 360102 700000 360108 700052
rect 360160 700040 360166 700052
rect 462314 700040 462320 700052
rect 360160 700012 462320 700040
rect 360160 700000 360166 700012
rect 462314 700000 462320 700012
rect 462372 700000 462378 700052
rect 283834 699932 283840 699984
rect 283892 699972 283898 699984
rect 385034 699972 385040 699984
rect 283892 699944 385040 699972
rect 283892 699932 283898 699944
rect 385034 699932 385040 699944
rect 385092 699932 385098 699984
rect 332502 699864 332508 699916
rect 332560 699904 332566 699916
rect 375374 699904 375380 699916
rect 332560 699876 375380 699904
rect 332560 699864 332566 699876
rect 375374 699864 375380 699876
rect 375432 699864 375438 699916
rect 371142 699796 371148 699848
rect 371200 699836 371206 699848
rect 413646 699836 413652 699848
rect 371200 699808 413652 699836
rect 371200 699796 371206 699808
rect 413646 699796 413652 699808
rect 413704 699796 413710 699848
rect 348786 699728 348792 699780
rect 348844 699768 348850 699780
rect 378134 699768 378140 699780
rect 348844 699740 378140 699768
rect 348844 699728 348850 699740
rect 378134 699728 378140 699740
rect 378192 699728 378198 699780
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 364978 699660 364984 699712
rect 365036 699700 365042 699712
rect 365622 699700 365628 699712
rect 365036 699672 365628 699700
rect 365036 699660 365042 699672
rect 365622 699660 365628 699672
rect 365680 699660 365686 699712
rect 368382 699660 368388 699712
rect 368440 699700 368446 699712
rect 397454 699700 397460 699712
rect 368440 699672 397460 699700
rect 368440 699660 368446 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 344922 696940 344928 696992
rect 344980 696980 344986 696992
rect 580166 696980 580172 696992
rect 344980 696952 580172 696980
rect 344980 696940 344986 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 429212 685936 429976 685964
rect 347682 685856 347688 685908
rect 347740 685896 347746 685908
rect 429212 685896 429240 685936
rect 347740 685868 429240 685896
rect 429948 685896 429976 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 429948 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 347740 685856 347746 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429473 684471 429531 684477
rect 429473 684468 429485 684471
rect 429344 684440 429485 684468
rect 429344 684428 429350 684440
rect 429473 684437 429485 684440
rect 429519 684437 429531 684471
rect 429473 684431 429531 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 419534 681748 419540 681760
rect 3568 681720 419540 681748
rect 3568 681708 3574 681720
rect 419534 681708 419540 681720
rect 419592 681708 419598 681760
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 342162 673480 342168 673532
rect 342220 673520 342226 673532
rect 580166 673520 580172 673532
rect 342220 673492 580172 673520
rect 342220 673480 342226 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 269022 670692 269028 670744
rect 269080 670732 269086 670744
rect 577498 670732 577504 670744
rect 269080 670704 577504 670732
rect 269080 670692 269086 670704
rect 577498 670692 577504 670704
rect 577556 670692 577562 670744
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 425054 667944 425060 667956
rect 3476 667916 425060 667944
rect 3476 667904 3482 667916
rect 425054 667904 425060 667916
rect 425112 667904 425118 667956
rect 429470 666584 429476 666596
rect 429431 666556 429476 666584
rect 429470 666544 429476 666556
rect 429528 666544 429534 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 429197 656863 429255 656869
rect 429197 656829 429209 656863
rect 429243 656860 429255 656863
rect 429286 656860 429292 656872
rect 429243 656832 429292 656860
rect 429243 656829 429255 656832
rect 429197 656823 429255 656829
rect 429286 656820 429292 656832
rect 429344 656820 429350 656872
rect 559190 656860 559196 656872
rect 559151 656832 559196 656860
rect 559190 656820 559196 656832
rect 559248 656820 559254 656872
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 422294 652780 422300 652792
rect 3108 652752 422300 652780
rect 3108 652740 3114 652752
rect 422294 652740 422300 652752
rect 422352 652740 422358 652792
rect 336642 650020 336648 650072
rect 336700 650060 336706 650072
rect 580166 650060 580172 650072
rect 336700 650032 580172 650060
rect 336700 650020 336706 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 429194 647272 429200 647284
rect 429155 647244 429200 647272
rect 429194 647232 429200 647244
rect 429252 647232 429258 647284
rect 559193 647275 559251 647281
rect 559193 647241 559205 647275
rect 559239 647272 559251 647275
rect 559282 647272 559288 647284
rect 559239 647244 559288 647272
rect 559239 647241 559251 647244
rect 559193 647235 559251 647241
rect 559282 647232 559288 647244
rect 559340 647232 559346 647284
rect 411254 645124 411260 645176
rect 411312 645164 411318 645176
rect 412542 645164 412548 645176
rect 411312 645136 412548 645164
rect 411312 645124 411318 645136
rect 412542 645124 412548 645136
rect 412600 645124 412606 645176
rect 365162 643968 365168 644020
rect 365220 644008 365226 644020
rect 429194 644008 429200 644020
rect 365220 643980 429200 644008
rect 365220 643968 365226 643980
rect 429194 643968 429200 643980
rect 429252 643968 429258 644020
rect 300762 643900 300768 643952
rect 300820 643940 300826 643952
rect 380986 643940 380992 643952
rect 300820 643912 380992 643940
rect 300820 643900 300826 643912
rect 380986 643900 380992 643912
rect 381044 643900 381050 643952
rect 357342 643832 357348 643884
rect 357400 643872 357406 643884
rect 494054 643872 494060 643884
rect 357400 643844 494060 643872
rect 357400 643832 357406 643844
rect 494054 643832 494060 643844
rect 494112 643832 494118 643884
rect 235902 643764 235908 643816
rect 235960 643804 235966 643816
rect 388898 643804 388904 643816
rect 235960 643776 388904 643804
rect 235960 643764 235966 643776
rect 388898 643764 388904 643776
rect 388956 643764 388962 643816
rect 349430 643696 349436 643748
rect 349488 643736 349494 643748
rect 559282 643736 559288 643748
rect 349488 643708 559288 643736
rect 349488 643696 349494 643708
rect 559282 643696 559288 643708
rect 559340 643696 559346 643748
rect 365622 643084 365628 643136
rect 365680 643124 365686 643136
rect 373074 643124 373080 643136
rect 365680 643096 373080 643124
rect 365680 643084 365686 643096
rect 373074 643084 373080 643096
rect 373132 643084 373138 643136
rect 427740 643096 427860 643124
rect 283650 643016 283656 643068
rect 283708 643056 283714 643068
rect 427740 643056 427768 643096
rect 427832 643068 427860 643096
rect 283708 643028 427768 643056
rect 283708 643016 283714 643028
rect 427814 643016 427820 643068
rect 427872 643016 427878 643068
rect 429010 643016 429016 643068
rect 429068 643056 429074 643068
rect 523126 643056 523132 643068
rect 429068 643028 523132 643056
rect 429068 643016 429074 643028
rect 523126 643016 523132 643028
rect 523184 643016 523190 643068
rect 307294 642948 307300 643000
rect 307352 642988 307358 643000
rect 473354 642988 473360 643000
rect 307352 642960 473360 642988
rect 307352 642948 307358 642960
rect 473354 642948 473360 642960
rect 473412 642948 473418 643000
rect 331030 642880 331036 642932
rect 331088 642920 331094 642932
rect 532326 642920 532332 642932
rect 331088 642892 532332 642920
rect 331088 642880 331094 642892
rect 532326 642880 532332 642892
rect 532384 642880 532390 642932
rect 265158 642812 265164 642864
rect 265216 642852 265222 642864
rect 320818 642852 320824 642864
rect 265216 642824 320824 642852
rect 265216 642812 265222 642824
rect 320818 642812 320824 642824
rect 320876 642812 320882 642864
rect 323118 642812 323124 642864
rect 323176 642852 323182 642864
rect 532234 642852 532240 642864
rect 323176 642824 532240 642852
rect 323176 642812 323182 642824
rect 532234 642812 532240 642824
rect 532292 642812 532298 642864
rect 320450 642744 320456 642796
rect 320508 642784 320514 642796
rect 530394 642784 530400 642796
rect 320508 642756 530400 642784
rect 320508 642744 320514 642756
rect 530394 642744 530400 642756
rect 530452 642744 530458 642796
rect 288894 642676 288900 642728
rect 288952 642716 288958 642728
rect 307662 642716 307668 642728
rect 288952 642688 307668 642716
rect 288952 642676 288958 642688
rect 307662 642676 307668 642688
rect 307720 642676 307726 642728
rect 315206 642676 315212 642728
rect 315264 642716 315270 642728
rect 532142 642716 532148 642728
rect 315264 642688 532148 642716
rect 315264 642676 315270 642688
rect 532142 642676 532148 642688
rect 532200 642676 532206 642728
rect 267826 642608 267832 642660
rect 267884 642648 267890 642660
rect 269022 642648 269028 642660
rect 267884 642620 269028 642648
rect 267884 642608 267890 642620
rect 269022 642608 269028 642620
rect 269080 642608 269086 642660
rect 304626 642608 304632 642660
rect 304684 642648 304690 642660
rect 532050 642648 532056 642660
rect 304684 642620 532056 642648
rect 304684 642608 304690 642620
rect 532050 642608 532056 642620
rect 532108 642608 532114 642660
rect 236270 642540 236276 642592
rect 236328 642580 236334 642592
rect 289998 642580 290004 642592
rect 236328 642552 290004 642580
rect 236328 642540 236334 642552
rect 289998 642540 290004 642552
rect 290056 642540 290062 642592
rect 294138 642540 294144 642592
rect 294196 642580 294202 642592
rect 531038 642580 531044 642592
rect 294196 642552 531044 642580
rect 294196 642540 294202 642552
rect 531038 642540 531044 642552
rect 531096 642540 531102 642592
rect 270494 642472 270500 642524
rect 270552 642512 270558 642524
rect 530670 642512 530676 642524
rect 270552 642484 530676 642512
rect 270552 642472 270558 642484
rect 530670 642472 530676 642484
rect 530728 642472 530734 642524
rect 252002 642404 252008 642456
rect 252060 642444 252066 642456
rect 263594 642444 263600 642456
rect 252060 642416 263600 642444
rect 252060 642404 252066 642416
rect 263594 642404 263600 642416
rect 263652 642404 263658 642456
rect 278314 642404 278320 642456
rect 278372 642444 278378 642456
rect 580902 642444 580908 642456
rect 278372 642416 580908 642444
rect 278372 642404 278378 642416
rect 580902 642404 580908 642416
rect 580960 642404 580966 642456
rect 257338 642336 257344 642388
rect 257396 642376 257402 642388
rect 580626 642376 580632 642388
rect 257396 642348 580632 642376
rect 257396 642336 257402 642348
rect 580626 642336 580632 642348
rect 580684 642336 580690 642388
rect 86218 642268 86224 642320
rect 86276 642308 86282 642320
rect 438854 642308 438860 642320
rect 86276 642280 438860 642308
rect 86276 642268 86282 642280
rect 438854 642268 438860 642280
rect 438912 642268 438918 642320
rect 438946 642268 438952 642320
rect 439004 642308 439010 642320
rect 454678 642308 454684 642320
rect 439004 642280 454684 642308
rect 439004 642268 439010 642280
rect 454678 642268 454684 642280
rect 454736 642268 454742 642320
rect 5442 642200 5448 642252
rect 5500 642240 5506 642252
rect 433610 642240 433616 642252
rect 5500 642212 433616 642240
rect 5500 642200 5506 642212
rect 433610 642200 433616 642212
rect 433668 642200 433674 642252
rect 5350 642132 5356 642184
rect 5408 642172 5414 642184
rect 441522 642172 441528 642184
rect 5408 642144 441528 642172
rect 5408 642132 5414 642144
rect 441522 642132 441528 642144
rect 441580 642132 441586 642184
rect 7926 642064 7932 642116
rect 7984 642104 7990 642116
rect 446766 642104 446772 642116
rect 7984 642076 446772 642104
rect 7984 642064 7990 642076
rect 446766 642064 446772 642076
rect 446824 642064 446830 642116
rect 446858 642064 446864 642116
rect 446916 642104 446922 642116
rect 486234 642104 486240 642116
rect 446916 642076 486240 642104
rect 446916 642064 446922 642076
rect 486234 642064 486240 642076
rect 486292 642064 486298 642116
rect 5258 641996 5264 642048
rect 5316 642036 5322 642048
rect 449434 642036 449440 642048
rect 5316 642008 449440 642036
rect 5316 641996 5322 642008
rect 449434 641996 449440 642008
rect 449492 641996 449498 642048
rect 7650 641928 7656 641980
rect 7708 641968 7714 641980
rect 462590 641968 462596 641980
rect 7708 641940 462596 641968
rect 7708 641928 7714 641940
rect 462590 641928 462596 641940
rect 462648 641928 462654 641980
rect 462958 641928 462964 641980
rect 463016 641968 463022 641980
rect 502058 641968 502064 641980
rect 463016 641940 502064 641968
rect 463016 641928 463022 641940
rect 502058 641928 502064 641940
rect 502116 641928 502122 641980
rect 5166 641860 5172 641912
rect 5224 641900 5230 641912
rect 465166 641900 465172 641912
rect 5224 641872 465172 641900
rect 5224 641860 5230 641872
rect 465166 641860 465172 641872
rect 465224 641860 465230 641912
rect 5074 641792 5080 641844
rect 5132 641832 5138 641844
rect 473078 641832 473084 641844
rect 5132 641804 473084 641832
rect 5132 641792 5138 641804
rect 473078 641792 473084 641804
rect 473136 641792 473142 641844
rect 485130 641792 485136 641844
rect 485188 641832 485194 641844
rect 517790 641832 517796 641844
rect 485188 641804 517796 641832
rect 485188 641792 485194 641804
rect 517790 641792 517796 641804
rect 517848 641792 517854 641844
rect 4982 641724 4988 641776
rect 5040 641764 5046 641776
rect 488902 641764 488908 641776
rect 5040 641736 488908 641764
rect 5040 641724 5046 641736
rect 488902 641724 488908 641736
rect 488960 641724 488966 641776
rect 325789 641699 325847 641705
rect 325789 641665 325801 641699
rect 325835 641696 325847 641699
rect 335173 641699 335231 641705
rect 335173 641696 335185 641699
rect 325835 641668 335185 641696
rect 325835 641665 325847 641668
rect 325789 641659 325847 641665
rect 335173 641665 335185 641668
rect 335219 641665 335231 641699
rect 335173 641659 335231 641665
rect 345017 641699 345075 641705
rect 345017 641665 345029 641699
rect 345063 641696 345075 641699
rect 354585 641699 354643 641705
rect 354585 641696 354597 641699
rect 345063 641668 354597 641696
rect 345063 641665 345075 641668
rect 345017 641659 345075 641665
rect 354585 641665 354597 641668
rect 354631 641665 354643 641699
rect 354585 641659 354643 641665
rect 364337 641699 364395 641705
rect 364337 641665 364349 641699
rect 364383 641696 364395 641699
rect 373905 641699 373963 641705
rect 373905 641696 373917 641699
rect 364383 641668 373917 641696
rect 364383 641665 364395 641668
rect 364337 641659 364395 641665
rect 373905 641665 373917 641668
rect 373951 641665 373963 641699
rect 373905 641659 373963 641665
rect 383657 641699 383715 641705
rect 383657 641665 383669 641699
rect 383703 641696 383715 641699
rect 393225 641699 393283 641705
rect 393225 641696 393237 641699
rect 383703 641668 393237 641696
rect 383703 641665 383715 641668
rect 383657 641659 383715 641665
rect 393225 641665 393237 641668
rect 393271 641665 393283 641699
rect 393225 641659 393283 641665
rect 402977 641699 403035 641705
rect 402977 641665 402989 641699
rect 403023 641696 403035 641699
rect 412545 641699 412603 641705
rect 412545 641696 412557 641699
rect 403023 641668 412557 641696
rect 403023 641665 403035 641668
rect 402977 641659 403035 641665
rect 412545 641665 412557 641668
rect 412591 641665 412603 641699
rect 412545 641659 412603 641665
rect 427814 641656 427820 641708
rect 427872 641696 427878 641708
rect 580350 641696 580356 641708
rect 427872 641668 580356 641696
rect 427872 641656 427878 641668
rect 580350 641656 580356 641668
rect 580408 641656 580414 641708
rect 333606 641588 333612 641640
rect 333664 641628 333670 641640
rect 530210 641628 530216 641640
rect 333664 641600 530216 641628
rect 333664 641588 333670 641600
rect 530210 641588 530216 641600
rect 530268 641588 530274 641640
rect 317782 641520 317788 641572
rect 317840 641560 317846 641572
rect 529842 641560 529848 641572
rect 317840 641532 529848 641560
rect 317840 641520 317846 641532
rect 529842 641520 529848 641532
rect 529900 641520 529906 641572
rect 312538 641452 312544 641504
rect 312596 641492 312602 641504
rect 530486 641492 530492 641504
rect 312596 641464 530492 641492
rect 312596 641452 312602 641464
rect 530486 641452 530492 641464
rect 530544 641452 530550 641504
rect 309962 641384 309968 641436
rect 310020 641424 310026 641436
rect 529750 641424 529756 641436
rect 310020 641396 529756 641424
rect 310020 641384 310026 641396
rect 529750 641384 529756 641396
rect 529808 641384 529814 641436
rect 299382 641316 299388 641368
rect 299440 641356 299446 641368
rect 531958 641356 531964 641368
rect 299440 641328 531964 641356
rect 299440 641316 299446 641328
rect 531958 641316 531964 641328
rect 532016 641316 532022 641368
rect 286226 641248 286232 641300
rect 286284 641288 286290 641300
rect 530946 641288 530952 641300
rect 286284 641260 530952 641288
rect 286284 641248 286290 641260
rect 530946 641248 530952 641260
rect 531004 641248 531010 641300
rect 275738 641180 275744 641232
rect 275796 641220 275802 641232
rect 530762 641220 530768 641232
rect 275796 641192 530768 641220
rect 275796 641180 275802 641192
rect 530762 641180 530768 641192
rect 530820 641180 530826 641232
rect 262582 641112 262588 641164
rect 262640 641152 262646 641164
rect 530578 641152 530584 641164
rect 262640 641124 530584 641152
rect 262640 641112 262646 641124
rect 530578 641112 530584 641124
rect 530636 641112 530642 641164
rect 246758 641044 246764 641096
rect 246816 641084 246822 641096
rect 529566 641084 529572 641096
rect 246816 641056 529572 641084
rect 246816 641044 246822 641056
rect 529566 641044 529572 641056
rect 529624 641044 529630 641096
rect 3970 640976 3976 641028
rect 4028 641016 4034 641028
rect 258718 641016 258724 641028
rect 4028 640988 258724 641016
rect 4028 640976 4034 640988
rect 258718 640976 258724 640988
rect 258776 640976 258782 641028
rect 291470 640976 291476 641028
rect 291528 641016 291534 641028
rect 580074 641016 580080 641028
rect 291528 640988 580080 641016
rect 291528 640976 291534 640988
rect 580074 640976 580080 640988
rect 580132 640976 580138 641028
rect 238846 640908 238852 640960
rect 238904 640948 238910 640960
rect 529474 640948 529480 640960
rect 238904 640920 529480 640948
rect 238904 640908 238910 640920
rect 529474 640908 529480 640920
rect 529532 640908 529538 640960
rect 8202 640840 8208 640892
rect 8260 640880 8266 640892
rect 428366 640880 428372 640892
rect 8260 640852 428372 640880
rect 8260 640840 8266 640852
rect 428366 640840 428372 640852
rect 428424 640840 428430 640892
rect 473354 640840 473360 640892
rect 473412 640880 473418 640892
rect 579890 640880 579896 640892
rect 473412 640852 579896 640880
rect 473412 640840 473418 640852
rect 579890 640840 579896 640852
rect 579948 640840 579954 640892
rect 8110 640772 8116 640824
rect 8168 640812 8174 640824
rect 431034 640812 431040 640824
rect 8168 640784 431040 640812
rect 8168 640772 8174 640784
rect 431034 640772 431040 640784
rect 431092 640772 431098 640824
rect 444190 640812 444196 640824
rect 440804 640784 444196 640812
rect 8018 640704 8024 640756
rect 8076 640744 8082 640756
rect 436278 640744 436284 640756
rect 8076 640716 436284 640744
rect 8076 640704 8082 640716
rect 436278 640704 436284 640716
rect 436336 640704 436342 640756
rect 6546 640636 6552 640688
rect 6604 640676 6610 640688
rect 440804 640676 440832 640784
rect 444190 640772 444196 640784
rect 444248 640772 444254 640824
rect 6604 640648 440832 640676
rect 441709 640679 441767 640685
rect 6604 640636 6610 640648
rect 441709 640645 441721 640679
rect 441755 640676 441767 640679
rect 445205 640679 445263 640685
rect 445205 640676 445217 640679
rect 441755 640648 445217 640676
rect 441755 640645 441767 640648
rect 441709 640639 441767 640645
rect 445205 640645 445217 640648
rect 445251 640645 445263 640679
rect 445205 640639 445263 640645
rect 6454 640568 6460 640620
rect 6512 640608 6518 640620
rect 452010 640608 452016 640620
rect 6512 640580 452016 640608
rect 6512 640568 6518 640580
rect 452010 640568 452016 640580
rect 452068 640568 452074 640620
rect 7742 640500 7748 640552
rect 7800 640540 7806 640552
rect 459922 640540 459928 640552
rect 7800 640512 459928 640540
rect 7800 640500 7806 640512
rect 459922 640500 459928 640512
rect 459980 640500 459986 640552
rect 6362 640432 6368 640484
rect 6420 640472 6426 640484
rect 467834 640472 467840 640484
rect 6420 640444 467840 640472
rect 6420 640432 6426 640444
rect 467834 640432 467840 640444
rect 467892 640432 467898 640484
rect 7558 640364 7564 640416
rect 7616 640404 7622 640416
rect 475746 640404 475752 640416
rect 7616 640376 475752 640404
rect 7616 640364 7622 640376
rect 475746 640364 475752 640376
rect 475804 640364 475810 640416
rect 4798 640296 4804 640348
rect 4856 640336 4862 640348
rect 515214 640336 515220 640348
rect 4856 640308 515220 640336
rect 4856 640296 4862 640308
rect 515214 640296 515220 640308
rect 515272 640296 515278 640348
rect 307113 640271 307171 640277
rect 307113 640237 307125 640271
rect 307159 640268 307171 640271
rect 311805 640271 311863 640277
rect 311805 640268 311817 640271
rect 307159 640240 311817 640268
rect 307159 640237 307171 640240
rect 307113 640231 307171 640237
rect 311805 640237 311817 640240
rect 311851 640237 311863 640271
rect 311805 640231 311863 640237
rect 320818 640228 320824 640280
rect 320876 640268 320882 640280
rect 580718 640268 580724 640280
rect 320876 640240 580724 640268
rect 320876 640228 320882 640240
rect 580718 640228 580724 640240
rect 580776 640228 580782 640280
rect 307662 640160 307668 640212
rect 307720 640200 307726 640212
rect 579982 640200 579988 640212
rect 307720 640172 579988 640200
rect 307720 640160 307726 640172
rect 579982 640160 579988 640172
rect 580040 640160 580046 640212
rect 287149 640135 287207 640141
rect 287149 640101 287161 640135
rect 287195 640132 287207 640135
rect 290553 640135 290611 640141
rect 290553 640132 290565 640135
rect 287195 640104 290565 640132
rect 287195 640101 287207 640104
rect 287149 640095 287207 640101
rect 290553 640101 290565 640104
rect 290599 640101 290611 640135
rect 290553 640095 290611 640101
rect 296806 640092 296812 640144
rect 296864 640132 296870 640144
rect 531130 640132 531136 640144
rect 296864 640104 531136 640132
rect 296864 640092 296870 640104
rect 531130 640092 531136 640104
rect 531188 640092 531194 640144
rect 267829 640067 267887 640073
rect 267829 640033 267841 640067
rect 267875 640064 267887 640067
rect 277213 640067 277271 640073
rect 277213 640064 277225 640067
rect 267875 640036 277225 640064
rect 267875 640033 267887 640036
rect 267829 640027 267887 640033
rect 277213 640033 277225 640036
rect 277259 640033 277271 640067
rect 277213 640027 277271 640033
rect 287057 640067 287115 640073
rect 287057 640033 287069 640067
rect 287103 640064 287115 640067
rect 292577 640067 292635 640073
rect 292577 640064 292589 640067
rect 287103 640036 292589 640064
rect 287103 640033 287115 640036
rect 287057 640027 287115 640033
rect 292577 640033 292589 640036
rect 292623 640033 292635 640067
rect 292577 640027 292635 640033
rect 307021 640067 307079 640073
rect 307021 640033 307033 640067
rect 307067 640064 307079 640067
rect 311897 640067 311955 640073
rect 311897 640064 311909 640067
rect 307067 640036 311909 640064
rect 307067 640033 307079 640036
rect 307021 640027 307079 640033
rect 311897 640033 311909 640036
rect 311943 640033 311955 640067
rect 311897 640027 311955 640033
rect 325789 640067 325847 640073
rect 325789 640033 325801 640067
rect 325835 640064 325847 640067
rect 336001 640067 336059 640073
rect 336001 640064 336013 640067
rect 325835 640036 336013 640064
rect 325835 640033 325847 640036
rect 325789 640027 325847 640033
rect 336001 640033 336013 640036
rect 336047 640033 336059 640067
rect 336001 640027 336059 640033
rect 339218 640024 339224 640076
rect 339276 640064 339282 640076
rect 580166 640064 580172 640076
rect 339276 640036 580172 640064
rect 339276 640024 339282 640036
rect 580166 640024 580172 640036
rect 580224 640024 580230 640076
rect 229738 639956 229744 640008
rect 229796 639996 229802 640008
rect 478046 639996 478052 640008
rect 229796 639968 478052 639996
rect 229796 639956 229802 639968
rect 478046 639956 478052 639968
rect 478104 639956 478110 640008
rect 220906 639888 220912 639940
rect 220964 639928 220970 639940
rect 235258 639928 235264 639940
rect 220964 639900 235264 639928
rect 220964 639888 220970 639900
rect 235258 639888 235264 639900
rect 235316 639888 235322 639940
rect 263594 639888 263600 639940
rect 263652 639928 263658 639940
rect 580534 639928 580540 639940
rect 263652 639900 580540 639928
rect 263652 639888 263658 639900
rect 580534 639888 580540 639900
rect 580592 639888 580598 639940
rect 229649 639863 229707 639869
rect 229649 639829 229661 639863
rect 229695 639860 229707 639863
rect 239309 639863 239367 639869
rect 239309 639860 239321 639863
rect 229695 639832 239321 639860
rect 229695 639829 229707 639832
rect 229649 639823 229707 639829
rect 239309 639829 239321 639832
rect 239355 639829 239367 639863
rect 239309 639823 239367 639829
rect 251821 639863 251879 639869
rect 251821 639829 251833 639863
rect 251867 639860 251879 639863
rect 257893 639863 257951 639869
rect 257893 639860 257905 639863
rect 251867 639832 257905 639860
rect 251867 639829 251879 639832
rect 251821 639823 251879 639829
rect 257893 639829 257905 639832
rect 257939 639829 257951 639863
rect 257893 639823 257951 639829
rect 267737 639863 267795 639869
rect 267737 639829 267749 639863
rect 267783 639860 267795 639863
rect 277305 639863 277363 639869
rect 277305 639860 277317 639863
rect 267783 639832 277317 639860
rect 267783 639829 267795 639832
rect 267737 639823 267795 639829
rect 277305 639829 277317 639832
rect 277351 639829 277363 639863
rect 277305 639823 277363 639829
rect 281258 639820 281264 639872
rect 281316 639860 281322 639872
rect 530854 639860 530860 639872
rect 281316 639832 530860 639860
rect 281316 639820 281322 639832
rect 530854 639820 530860 639832
rect 530912 639820 530918 639872
rect 229741 639795 229799 639801
rect 229741 639761 229753 639795
rect 229787 639792 229799 639795
rect 239401 639795 239459 639801
rect 239401 639792 239413 639795
rect 229787 639764 239413 639792
rect 229787 639761 229799 639764
rect 229741 639755 229799 639761
rect 239401 639761 239413 639764
rect 239447 639761 239459 639795
rect 239401 639755 239459 639761
rect 247589 639795 247647 639801
rect 247589 639761 247601 639795
rect 247635 639792 247647 639795
rect 257985 639795 258043 639801
rect 257985 639792 257997 639795
rect 247635 639764 257997 639792
rect 247635 639761 247647 639764
rect 247589 639755 247647 639761
rect 257985 639761 257997 639764
rect 258031 639761 258043 639795
rect 257985 639755 258043 639761
rect 273162 639752 273168 639804
rect 273220 639792 273226 639804
rect 580810 639792 580816 639804
rect 273220 639764 580816 639792
rect 273220 639752 273226 639764
rect 580810 639752 580816 639764
rect 580868 639752 580874 639804
rect 3326 639684 3332 639736
rect 3384 639724 3390 639736
rect 438946 639724 438952 639736
rect 3384 639696 438952 639724
rect 3384 639684 3390 639696
rect 438946 639684 438952 639696
rect 439004 639684 439010 639736
rect 441617 639727 441675 639733
rect 441617 639693 441629 639727
rect 441663 639724 441675 639727
rect 457070 639724 457076 639736
rect 441663 639696 457076 639724
rect 441663 639693 441675 639696
rect 441617 639687 441675 639693
rect 457070 639684 457076 639696
rect 457128 639684 457134 639736
rect 463697 639727 463755 639733
rect 463697 639693 463709 639727
rect 463743 639724 463755 639727
rect 473265 639727 473323 639733
rect 473265 639724 473277 639727
rect 463743 639696 473277 639724
rect 463743 639693 463755 639696
rect 463697 639687 463755 639693
rect 473265 639693 473277 639696
rect 473311 639693 473323 639727
rect 473265 639687 473323 639693
rect 4062 639616 4068 639668
rect 4120 639656 4126 639668
rect 408313 639659 408371 639665
rect 408313 639656 408325 639659
rect 4120 639628 408325 639656
rect 4120 639616 4126 639628
rect 408313 639625 408325 639628
rect 408359 639625 408371 639659
rect 408313 639619 408371 639625
rect 408497 639659 408555 639665
rect 408497 639625 408509 639659
rect 408543 639656 408555 639659
rect 446858 639656 446864 639668
rect 408543 639628 446864 639656
rect 408543 639625 408555 639628
rect 408497 639619 408555 639625
rect 446858 639616 446864 639628
rect 446916 639616 446922 639668
rect 480622 639656 480628 639668
rect 476040 639628 480628 639656
rect 7834 639548 7840 639600
rect 7892 639588 7898 639600
rect 37369 639591 37427 639597
rect 37369 639588 37381 639591
rect 7892 639560 37381 639588
rect 7892 639548 7898 639560
rect 37369 639557 37381 639560
rect 37415 639557 37427 639591
rect 37369 639551 37427 639557
rect 37461 639591 37519 639597
rect 37461 639557 37473 639591
rect 37507 639588 37519 639591
rect 193217 639591 193275 639597
rect 193217 639588 193229 639591
rect 37507 639560 193229 639588
rect 37507 639557 37519 639560
rect 37461 639551 37519 639557
rect 193217 639557 193229 639560
rect 193263 639557 193275 639591
rect 193217 639551 193275 639557
rect 193401 639591 193459 639597
rect 193401 639557 193413 639591
rect 193447 639588 193459 639591
rect 212629 639591 212687 639597
rect 212629 639588 212641 639591
rect 193447 639560 212641 639588
rect 193447 639557 193459 639560
rect 193401 639551 193459 639557
rect 212629 639557 212641 639560
rect 212675 639557 212687 639591
rect 212629 639551 212687 639557
rect 212721 639591 212779 639597
rect 212721 639557 212733 639591
rect 212767 639588 212779 639591
rect 229741 639591 229799 639597
rect 229741 639588 229753 639591
rect 212767 639560 229753 639588
rect 212767 639557 212779 639560
rect 212721 639551 212779 639557
rect 229741 639557 229753 639560
rect 229787 639557 229799 639591
rect 229741 639551 229799 639557
rect 239309 639591 239367 639597
rect 239309 639557 239321 639591
rect 239355 639557 239367 639591
rect 239309 639551 239367 639557
rect 239401 639591 239459 639597
rect 239401 639557 239413 639591
rect 239447 639588 239459 639591
rect 247589 639591 247647 639597
rect 247589 639588 247601 639591
rect 239447 639560 247601 639588
rect 239447 639557 239459 639560
rect 239401 639551 239459 639557
rect 247589 639557 247601 639560
rect 247635 639557 247647 639591
rect 247589 639551 247647 639557
rect 251821 639591 251879 639597
rect 251821 639557 251833 639591
rect 251867 639557 251879 639591
rect 251821 639551 251879 639557
rect 257893 639591 257951 639597
rect 257893 639557 257905 639591
rect 257939 639557 257951 639591
rect 257893 639551 257951 639557
rect 257985 639591 258043 639597
rect 257985 639557 257997 639591
rect 258031 639588 258043 639591
rect 267737 639591 267795 639597
rect 267737 639588 267749 639591
rect 258031 639560 267749 639588
rect 258031 639557 258043 639560
rect 257985 639551 258043 639557
rect 267737 639557 267749 639560
rect 267783 639557 267795 639591
rect 267737 639551 267795 639557
rect 267829 639591 267887 639597
rect 267829 639557 267841 639591
rect 267875 639557 267887 639591
rect 267829 639551 267887 639557
rect 277213 639591 277271 639597
rect 277213 639557 277225 639591
rect 277259 639557 277271 639591
rect 277213 639551 277271 639557
rect 277305 639591 277363 639597
rect 277305 639557 277317 639591
rect 277351 639588 277363 639591
rect 287057 639591 287115 639597
rect 287057 639588 287069 639591
rect 277351 639560 287069 639588
rect 277351 639557 277363 639560
rect 277305 639551 277363 639557
rect 287057 639557 287069 639560
rect 287103 639557 287115 639591
rect 287057 639551 287115 639557
rect 287149 639591 287207 639597
rect 287149 639557 287161 639591
rect 287195 639557 287207 639591
rect 287149 639551 287207 639557
rect 290553 639591 290611 639597
rect 290553 639557 290565 639591
rect 290599 639557 290611 639591
rect 290553 639551 290611 639557
rect 292577 639591 292635 639597
rect 292577 639557 292589 639591
rect 292623 639588 292635 639591
rect 307021 639591 307079 639597
rect 307021 639588 307033 639591
rect 292623 639560 307033 639588
rect 292623 639557 292635 639560
rect 292577 639551 292635 639557
rect 307021 639557 307033 639560
rect 307067 639557 307079 639591
rect 307021 639551 307079 639557
rect 307113 639591 307171 639597
rect 307113 639557 307125 639591
rect 307159 639557 307171 639591
rect 307113 639551 307171 639557
rect 311805 639591 311863 639597
rect 311805 639557 311817 639591
rect 311851 639557 311863 639591
rect 311805 639551 311863 639557
rect 311897 639591 311955 639597
rect 311897 639557 311909 639591
rect 311943 639588 311955 639591
rect 325789 639591 325847 639597
rect 325789 639588 325801 639591
rect 311943 639560 325801 639588
rect 311943 639557 311955 639560
rect 311897 639551 311955 639557
rect 325789 639557 325801 639560
rect 325835 639557 325847 639591
rect 325789 639551 325847 639557
rect 325881 639591 325939 639597
rect 325881 639557 325893 639591
rect 325927 639557 325939 639591
rect 325881 639551 325939 639557
rect 335173 639591 335231 639597
rect 335173 639557 335185 639591
rect 335219 639557 335231 639591
rect 335173 639551 335231 639557
rect 336001 639591 336059 639597
rect 336001 639557 336013 639591
rect 336047 639588 336059 639591
rect 345017 639591 345075 639597
rect 345017 639588 345029 639591
rect 336047 639560 345029 639588
rect 336047 639557 336059 639560
rect 336001 639551 336059 639557
rect 345017 639557 345029 639560
rect 345063 639557 345075 639591
rect 354585 639591 354643 639597
rect 345017 639551 345075 639557
rect 345124 639560 354536 639588
rect 5534 639480 5540 639532
rect 5592 639520 5598 639532
rect 23290 639520 23296 639532
rect 5592 639492 23296 639520
rect 5592 639480 5598 639492
rect 23290 639480 23296 639492
rect 23348 639480 23354 639532
rect 24765 639523 24823 639529
rect 24765 639489 24777 639523
rect 24811 639520 24823 639523
rect 27617 639523 27675 639529
rect 27617 639520 27629 639523
rect 24811 639492 27629 639520
rect 24811 639489 24823 639492
rect 24765 639483 24823 639489
rect 27617 639489 27629 639492
rect 27663 639489 27675 639523
rect 27617 639483 27675 639489
rect 37185 639523 37243 639529
rect 37185 639489 37197 639523
rect 37231 639520 37243 639523
rect 37277 639523 37335 639529
rect 37277 639520 37289 639523
rect 37231 639492 37289 639520
rect 37231 639489 37243 639492
rect 37185 639483 37243 639489
rect 37277 639489 37289 639492
rect 37323 639489 37335 639523
rect 37277 639483 37335 639489
rect 46937 639523 46995 639529
rect 46937 639489 46949 639523
rect 46983 639520 46995 639523
rect 60645 639523 60703 639529
rect 60645 639520 60657 639523
rect 46983 639492 60657 639520
rect 46983 639489 46995 639492
rect 46937 639483 46995 639489
rect 60645 639489 60657 639492
rect 60691 639489 60703 639523
rect 60645 639483 60703 639489
rect 67637 639523 67695 639529
rect 67637 639489 67649 639523
rect 67683 639520 67695 639523
rect 75917 639523 75975 639529
rect 75917 639520 75929 639523
rect 67683 639492 75929 639520
rect 67683 639489 67695 639492
rect 67637 639483 67695 639489
rect 75917 639489 75929 639492
rect 75963 639489 75975 639523
rect 75917 639483 75975 639489
rect 86957 639523 87015 639529
rect 86957 639489 86969 639523
rect 87003 639520 87015 639523
rect 99285 639523 99343 639529
rect 99285 639520 99297 639523
rect 87003 639492 99297 639520
rect 87003 639489 87015 639492
rect 86957 639483 87015 639489
rect 99285 639489 99297 639492
rect 99331 639489 99343 639523
rect 99285 639483 99343 639489
rect 106277 639523 106335 639529
rect 106277 639489 106289 639523
rect 106323 639520 106335 639523
rect 118605 639523 118663 639529
rect 118605 639520 118617 639523
rect 106323 639492 118617 639520
rect 106323 639489 106335 639492
rect 106277 639483 106335 639489
rect 118605 639489 118617 639492
rect 118651 639489 118663 639523
rect 118605 639483 118663 639489
rect 125597 639523 125655 639529
rect 125597 639489 125609 639523
rect 125643 639520 125655 639523
rect 153197 639523 153255 639529
rect 153197 639520 153209 639523
rect 125643 639492 143488 639520
rect 125643 639489 125655 639492
rect 125597 639483 125655 639489
rect 6270 639412 6276 639464
rect 6328 639452 6334 639464
rect 15197 639455 15255 639461
rect 15197 639452 15209 639455
rect 6328 639424 15209 639452
rect 6328 639412 6334 639424
rect 15197 639421 15209 639424
rect 15243 639421 15255 639455
rect 15197 639415 15255 639421
rect 60829 639455 60887 639461
rect 60829 639421 60841 639455
rect 60875 639452 60887 639455
rect 85485 639455 85543 639461
rect 60875 639424 67680 639452
rect 60875 639421 60887 639424
rect 60829 639415 60887 639421
rect 67652 639393 67680 639424
rect 85485 639421 85497 639455
rect 85531 639452 85543 639455
rect 99469 639455 99527 639461
rect 85531 639424 87000 639452
rect 85531 639421 85543 639424
rect 85485 639415 85543 639421
rect 86972 639393 87000 639424
rect 99469 639421 99481 639455
rect 99515 639452 99527 639455
rect 118789 639455 118847 639461
rect 99515 639424 106320 639452
rect 99515 639421 99527 639424
rect 99469 639415 99527 639421
rect 106292 639393 106320 639424
rect 118789 639421 118801 639455
rect 118835 639452 118847 639455
rect 143460 639452 143488 639492
rect 148244 639492 153209 639520
rect 118835 639424 125640 639452
rect 143460 639424 143580 639452
rect 118835 639421 118847 639424
rect 118789 639415 118847 639421
rect 125612 639393 125640 639424
rect 143552 639393 143580 639424
rect 67637 639387 67695 639393
rect 67637 639353 67649 639387
rect 67683 639353 67695 639387
rect 67637 639347 67695 639353
rect 86957 639387 87015 639393
rect 86957 639353 86969 639387
rect 87003 639353 87015 639387
rect 86957 639347 87015 639353
rect 106277 639387 106335 639393
rect 106277 639353 106289 639387
rect 106323 639353 106335 639387
rect 106277 639347 106335 639353
rect 125597 639387 125655 639393
rect 125597 639353 125609 639387
rect 125643 639353 125655 639387
rect 125597 639347 125655 639353
rect 143537 639387 143595 639393
rect 143537 639353 143549 639387
rect 143583 639353 143595 639387
rect 143537 639347 143595 639353
rect 143629 639387 143687 639393
rect 143629 639353 143641 639387
rect 143675 639384 143687 639387
rect 148244 639384 148272 639492
rect 153197 639489 153209 639492
rect 153243 639489 153255 639523
rect 153197 639483 153255 639489
rect 156322 639480 156328 639532
rect 156380 639520 156386 639532
rect 162670 639520 162676 639532
rect 156380 639492 162676 639520
rect 156380 639480 156386 639492
rect 162670 639480 162676 639492
rect 162728 639480 162734 639532
rect 164237 639523 164295 639529
rect 164237 639489 164249 639523
rect 164283 639520 164295 639523
rect 176565 639523 176623 639529
rect 176565 639520 176577 639523
rect 164283 639492 176577 639520
rect 164283 639489 164295 639492
rect 164237 639483 164295 639489
rect 176565 639489 176577 639492
rect 176611 639489 176623 639523
rect 176565 639483 176623 639489
rect 183557 639523 183615 639529
rect 183557 639489 183569 639523
rect 183603 639520 183615 639523
rect 195885 639523 195943 639529
rect 195885 639520 195897 639523
rect 183603 639492 195897 639520
rect 183603 639489 183615 639492
rect 183557 639483 183615 639489
rect 195885 639489 195897 639492
rect 195931 639489 195943 639523
rect 195885 639483 195943 639489
rect 201494 639480 201500 639532
rect 201552 639520 201558 639532
rect 211062 639520 211068 639532
rect 201552 639492 211068 639520
rect 201552 639480 201558 639492
rect 211062 639480 211068 639492
rect 211120 639480 211126 639532
rect 212537 639523 212595 639529
rect 212537 639520 212549 639523
rect 212460 639492 212549 639520
rect 212460 639461 212488 639492
rect 212537 639489 212549 639492
rect 212583 639489 212595 639523
rect 239324 639520 239352 639551
rect 251836 639520 251864 639551
rect 239324 639492 251864 639520
rect 257908 639520 257936 639551
rect 267844 639520 267872 639551
rect 257908 639492 267872 639520
rect 277228 639520 277256 639551
rect 287164 639520 287192 639551
rect 277228 639492 287192 639520
rect 290568 639520 290596 639551
rect 307128 639520 307156 639551
rect 290568 639492 307156 639520
rect 311820 639520 311848 639551
rect 325896 639520 325924 639551
rect 311820 639492 325924 639520
rect 335188 639520 335216 639551
rect 345124 639520 345152 639560
rect 335188 639492 345152 639520
rect 354508 639520 354536 639560
rect 354585 639557 354597 639591
rect 354631 639588 354643 639591
rect 364337 639591 364395 639597
rect 364337 639588 364349 639591
rect 354631 639560 364349 639588
rect 354631 639557 354643 639560
rect 354585 639551 354643 639557
rect 364337 639557 364349 639560
rect 364383 639557 364395 639591
rect 373905 639591 373963 639597
rect 364337 639551 364395 639557
rect 364996 639560 373856 639588
rect 364996 639520 365024 639560
rect 354508 639492 365024 639520
rect 373828 639520 373856 639560
rect 373905 639557 373917 639591
rect 373951 639588 373963 639591
rect 383657 639591 383715 639597
rect 383657 639588 383669 639591
rect 373951 639560 383669 639588
rect 373951 639557 373963 639560
rect 373905 639551 373963 639557
rect 383657 639557 383669 639560
rect 383703 639557 383715 639591
rect 393225 639591 393283 639597
rect 383657 639551 383715 639557
rect 384316 639560 393176 639588
rect 384316 639520 384344 639560
rect 373828 639492 384344 639520
rect 393148 639520 393176 639560
rect 393225 639557 393237 639591
rect 393271 639588 393283 639591
rect 402977 639591 403035 639597
rect 402977 639588 402989 639591
rect 393271 639560 402989 639588
rect 393271 639557 393283 639560
rect 393225 639551 393283 639557
rect 402977 639557 402989 639560
rect 403023 639557 403035 639591
rect 402977 639551 403035 639557
rect 412545 639591 412603 639597
rect 412545 639557 412557 639591
rect 412591 639588 412603 639591
rect 441617 639591 441675 639597
rect 441617 639588 441629 639591
rect 412591 639560 441629 639588
rect 412591 639557 412603 639560
rect 412545 639551 412603 639557
rect 441617 639557 441629 639560
rect 441663 639557 441675 639591
rect 441617 639551 441675 639557
rect 441709 639591 441767 639597
rect 441709 639557 441721 639591
rect 441755 639557 441767 639591
rect 441709 639551 441767 639557
rect 445205 639591 445263 639597
rect 445205 639557 445217 639591
rect 445251 639557 445263 639591
rect 445205 639551 445263 639557
rect 463697 639591 463755 639597
rect 463697 639557 463709 639591
rect 463743 639557 463755 639591
rect 463697 639551 463755 639557
rect 473265 639591 473323 639597
rect 473265 639557 473277 639591
rect 473311 639588 473323 639591
rect 476040 639588 476068 639628
rect 480622 639616 480628 639628
rect 480680 639616 480686 639668
rect 473311 639560 476068 639588
rect 473311 639557 473323 639560
rect 473265 639551 473323 639557
rect 441724 639520 441752 639551
rect 393148 639492 441752 639520
rect 445220 639520 445248 639551
rect 463712 639520 463740 639551
rect 445220 639492 463740 639520
rect 212537 639483 212595 639489
rect 153565 639455 153623 639461
rect 153565 639421 153577 639455
rect 153611 639452 153623 639455
rect 176749 639455 176807 639461
rect 153611 639424 164280 639452
rect 153611 639421 153623 639424
rect 153565 639415 153623 639421
rect 164252 639393 164280 639424
rect 176749 639421 176761 639455
rect 176795 639452 176807 639455
rect 195977 639455 196035 639461
rect 176795 639424 183600 639452
rect 176795 639421 176807 639424
rect 176749 639415 176807 639421
rect 183572 639393 183600 639424
rect 195977 639421 195989 639455
rect 196023 639452 196035 639455
rect 202877 639455 202935 639461
rect 202877 639452 202889 639455
rect 196023 639424 202889 639452
rect 196023 639421 196035 639424
rect 195977 639415 196035 639421
rect 202877 639421 202889 639424
rect 202923 639421 202935 639455
rect 202877 639415 202935 639421
rect 212445 639455 212503 639461
rect 212445 639421 212457 639455
rect 212491 639421 212503 639455
rect 212445 639415 212503 639421
rect 212629 639455 212687 639461
rect 212629 639421 212641 639455
rect 212675 639452 212687 639455
rect 229649 639455 229707 639461
rect 229649 639452 229661 639455
rect 212675 639424 229661 639452
rect 212675 639421 212687 639424
rect 212629 639415 212687 639421
rect 229649 639421 229661 639424
rect 229695 639421 229707 639455
rect 229649 639415 229707 639421
rect 143675 639356 148272 639384
rect 164237 639387 164295 639393
rect 143675 639353 143687 639356
rect 143629 639347 143687 639353
rect 164237 639353 164249 639387
rect 164283 639353 164295 639387
rect 164237 639347 164295 639353
rect 183557 639387 183615 639393
rect 183557 639353 183569 639387
rect 183603 639353 183615 639387
rect 183557 639347 183615 639353
rect 15197 639319 15255 639325
rect 15197 639285 15209 639319
rect 15243 639316 15255 639319
rect 24765 639319 24823 639325
rect 24765 639316 24777 639319
rect 15243 639288 24777 639316
rect 15243 639285 15255 639288
rect 15197 639279 15255 639285
rect 24765 639285 24777 639288
rect 24811 639285 24823 639319
rect 24765 639279 24823 639285
rect 27617 639319 27675 639325
rect 27617 639285 27629 639319
rect 27663 639316 27675 639319
rect 37185 639319 37243 639325
rect 37185 639316 37197 639319
rect 27663 639288 37197 639316
rect 27663 639285 27675 639288
rect 27617 639279 27675 639285
rect 37185 639285 37197 639288
rect 37231 639285 37243 639319
rect 37185 639279 37243 639285
rect 37277 639319 37335 639325
rect 37277 639285 37289 639319
rect 37323 639316 37335 639319
rect 46937 639319 46995 639325
rect 46937 639316 46949 639319
rect 37323 639288 46949 639316
rect 37323 639285 37335 639288
rect 37277 639279 37335 639285
rect 46937 639285 46949 639288
rect 46983 639285 46995 639319
rect 46937 639279 46995 639285
rect 75917 639319 75975 639325
rect 75917 639285 75929 639319
rect 75963 639316 75975 639319
rect 85485 639319 85543 639325
rect 85485 639316 85497 639319
rect 75963 639288 85497 639316
rect 75963 639285 75975 639288
rect 75917 639279 75975 639285
rect 85485 639285 85497 639288
rect 85531 639285 85543 639319
rect 85485 639279 85543 639285
rect 202877 639319 202935 639325
rect 202877 639285 202889 639319
rect 202923 639316 202935 639319
rect 212445 639319 212503 639325
rect 212445 639316 212457 639319
rect 202923 639288 212457 639316
rect 202923 639285 202935 639288
rect 202877 639279 202935 639285
rect 212445 639285 212457 639288
rect 212491 639285 212503 639319
rect 212445 639279 212503 639285
rect 60642 639208 60648 639260
rect 60700 639248 60706 639260
rect 66162 639248 66168 639260
rect 60700 639220 66168 639248
rect 60700 639208 60706 639220
rect 66162 639208 66168 639220
rect 66220 639208 66226 639260
rect 579798 639140 579804 639192
rect 579856 639180 579862 639192
rect 580350 639180 580356 639192
rect 579856 639152 580356 639180
rect 579856 639140 579862 639152
rect 580350 639140 580356 639152
rect 580408 639140 580414 639192
rect 530210 627852 530216 627904
rect 530268 627892 530274 627904
rect 579798 627892 579804 627904
rect 530268 627864 579804 627892
rect 530268 627852 530274 627864
rect 579798 627852 579804 627864
rect 579856 627852 579862 627904
rect 3234 624860 3240 624912
rect 3292 624900 3298 624912
rect 8202 624900 8208 624912
rect 3292 624872 8208 624900
rect 3292 624860 3298 624872
rect 8202 624860 8208 624872
rect 8260 624860 8266 624912
rect 2774 610580 2780 610632
rect 2832 610620 2838 610632
rect 5442 610620 5448 610632
rect 2832 610592 5448 610620
rect 2832 610580 2838 610592
rect 5442 610580 5448 610592
rect 5500 610580 5506 610632
rect 530302 604392 530308 604444
rect 530360 604432 530366 604444
rect 579798 604432 579804 604444
rect 530360 604404 579804 604432
rect 530360 604392 530366 604404
rect 579798 604392 579804 604404
rect 579856 604392 579862 604444
rect 3234 596028 3240 596080
rect 3292 596068 3298 596080
rect 8110 596068 8116 596080
rect 3292 596040 8116 596068
rect 3292 596028 3298 596040
rect 8110 596028 8116 596040
rect 8168 596028 8174 596080
rect 532326 593308 532332 593360
rect 532384 593348 532390 593360
rect 579798 593348 579804 593360
rect 532384 593320 579804 593348
rect 532384 593308 532390 593320
rect 579798 593308 579804 593320
rect 579856 593308 579862 593360
rect 3234 567740 3240 567792
rect 3292 567780 3298 567792
rect 8018 567780 8024 567792
rect 3292 567752 8024 567780
rect 3292 567740 3298 567752
rect 8018 567740 8024 567752
rect 8076 567740 8082 567792
rect 530394 557472 530400 557524
rect 530452 557512 530458 557524
rect 579798 557512 579804 557524
rect 530452 557484 579804 557512
rect 530452 557472 530458 557484
rect 579798 557472 579804 557484
rect 579856 557472 579862 557524
rect 2774 553052 2780 553104
rect 2832 553092 2838 553104
rect 5350 553092 5356 553104
rect 2832 553064 5356 553092
rect 2832 553052 2838 553064
rect 5350 553052 5356 553064
rect 5408 553052 5414 553104
rect 532234 546388 532240 546440
rect 532292 546428 532298 546440
rect 579798 546428 579804 546440
rect 532292 546400 579804 546428
rect 532292 546388 532298 546400
rect 579798 546388 579804 546400
rect 579856 546388 579862 546440
rect 3234 539520 3240 539572
rect 3292 539560 3298 539572
rect 86218 539560 86224 539572
rect 3292 539532 86224 539560
rect 3292 539520 3298 539532
rect 86218 539520 86224 539532
rect 86276 539520 86282 539572
rect 529842 534012 529848 534064
rect 529900 534052 529906 534064
rect 579798 534052 579804 534064
rect 529900 534024 579804 534052
rect 529900 534012 529906 534024
rect 579798 534012 579804 534024
rect 579856 534012 579862 534064
rect 530486 510552 530492 510604
rect 530544 510592 530550 510604
rect 579798 510592 579804 510604
rect 530544 510564 579804 510592
rect 530544 510552 530550 510564
rect 579798 510552 579804 510564
rect 579856 510552 579862 510604
rect 3234 510348 3240 510400
rect 3292 510388 3298 510400
rect 6546 510388 6552 510400
rect 3292 510360 6552 510388
rect 3292 510348 3298 510360
rect 6546 510348 6552 510360
rect 6604 510348 6610 510400
rect 532142 499468 532148 499520
rect 532200 499508 532206 499520
rect 579798 499508 579804 499520
rect 532200 499480 579804 499508
rect 532200 499468 532206 499480
rect 579798 499468 579804 499480
rect 579856 499468 579862 499520
rect 2774 496680 2780 496732
rect 2832 496720 2838 496732
rect 5258 496720 5264 496732
rect 2832 496692 5264 496720
rect 2832 496680 2838 496692
rect 5258 496680 5264 496692
rect 5316 496680 5322 496732
rect 529750 487092 529756 487144
rect 529808 487132 529814 487144
rect 579798 487132 579804 487144
rect 529808 487104 579804 487132
rect 529808 487092 529814 487104
rect 579798 487092 579804 487104
rect 579856 487092 579862 487144
rect 3234 481108 3240 481160
rect 3292 481148 3298 481160
rect 7926 481148 7932 481160
rect 3292 481120 7932 481148
rect 3292 481108 3298 481120
rect 7926 481108 7932 481120
rect 7984 481108 7990 481160
rect 532050 463632 532056 463684
rect 532108 463672 532114 463684
rect 579798 463672 579804 463684
rect 532108 463644 579804 463672
rect 532108 463632 532114 463644
rect 579798 463632 579804 463644
rect 579856 463632 579862 463684
rect 3142 452412 3148 452464
rect 3200 452452 3206 452464
rect 6454 452452 6460 452464
rect 3200 452424 6460 452452
rect 3200 452412 3206 452424
rect 6454 452412 6460 452424
rect 6512 452412 6518 452464
rect 531222 440172 531228 440224
rect 531280 440212 531286 440224
rect 579890 440212 579896 440224
rect 531280 440184 579896 440212
rect 531280 440172 531286 440184
rect 579890 440172 579896 440184
rect 579948 440172 579954 440224
rect 3142 438744 3148 438796
rect 3200 438784 3206 438796
rect 7834 438784 7840 438796
rect 3200 438756 7840 438784
rect 3200 438744 3206 438756
rect 7834 438744 7840 438756
rect 7892 438744 7898 438796
rect 531130 416712 531136 416764
rect 531188 416752 531194 416764
rect 579890 416752 579896 416764
rect 531188 416724 579896 416752
rect 531188 416712 531194 416724
rect 579890 416712 579896 416724
rect 579948 416712 579954 416764
rect 531958 405628 531964 405680
rect 532016 405668 532022 405680
rect 579890 405668 579896 405680
rect 532016 405640 579896 405668
rect 532016 405628 532022 405640
rect 579890 405628 579896 405640
rect 579948 405628 579954 405680
rect 3142 395428 3148 395480
rect 3200 395468 3206 395480
rect 7742 395468 7748 395480
rect 3200 395440 7748 395468
rect 3200 395428 3206 395440
rect 7742 395428 7748 395440
rect 7800 395428 7806 395480
rect 531038 393252 531044 393304
rect 531096 393292 531102 393304
rect 579890 393292 579896 393304
rect 531096 393264 579896 393292
rect 531096 393252 531102 393264
rect 579890 393252 579896 393264
rect 579948 393252 579954 393304
rect 2774 380604 2780 380656
rect 2832 380644 2838 380656
rect 5166 380644 5172 380656
rect 2832 380616 5172 380644
rect 2832 380604 2838 380616
rect 5166 380604 5172 380616
rect 5224 380604 5230 380656
rect 3326 366460 3332 366512
rect 3384 366500 3390 366512
rect 7650 366500 7656 366512
rect 3384 366472 7656 366500
rect 3384 366460 3390 366472
rect 7650 366460 7656 366472
rect 7708 366460 7714 366512
rect 530946 346332 530952 346384
rect 531004 346372 531010 346384
rect 579798 346372 579804 346384
rect 531004 346344 579804 346372
rect 531004 346332 531010 346344
rect 579798 346332 579804 346344
rect 579856 346332 579862 346384
rect 385037 338147 385095 338153
rect 385037 338113 385049 338147
rect 385083 338144 385095 338147
rect 395433 338147 395491 338153
rect 395433 338144 395445 338147
rect 385083 338116 395445 338144
rect 385083 338113 385095 338116
rect 385037 338107 385095 338113
rect 395433 338113 395445 338116
rect 395479 338113 395491 338147
rect 395433 338107 395491 338113
rect 71038 338036 71044 338088
rect 71096 338076 71102 338088
rect 264882 338076 264888 338088
rect 71096 338048 264888 338076
rect 71096 338036 71102 338048
rect 264882 338036 264888 338048
rect 264940 338036 264946 338088
rect 295613 338079 295671 338085
rect 295613 338045 295625 338079
rect 295659 338076 295671 338079
rect 295794 338076 295800 338088
rect 295659 338048 295800 338076
rect 295659 338045 295671 338048
rect 295613 338039 295671 338045
rect 295794 338036 295800 338048
rect 295852 338036 295858 338088
rect 332502 338036 332508 338088
rect 332560 338076 332566 338088
rect 400214 338076 400220 338088
rect 332560 338048 400220 338076
rect 332560 338036 332566 338048
rect 400214 338036 400220 338048
rect 400272 338036 400278 338088
rect 404998 338036 405004 338088
rect 405056 338076 405062 338088
rect 411806 338076 411812 338088
rect 405056 338048 411812 338076
rect 405056 338036 405062 338048
rect 411806 338036 411812 338048
rect 411864 338036 411870 338088
rect 412082 338036 412088 338088
rect 412140 338076 412146 338088
rect 419166 338076 419172 338088
rect 412140 338048 419172 338076
rect 412140 338036 412146 338048
rect 419166 338036 419172 338048
rect 419224 338036 419230 338088
rect 421009 338079 421067 338085
rect 421009 338045 421021 338079
rect 421055 338076 421067 338079
rect 427446 338076 427452 338088
rect 421055 338048 427452 338076
rect 421055 338045 421067 338048
rect 421009 338039 421067 338045
rect 427446 338036 427452 338048
rect 427504 338036 427510 338088
rect 427541 338079 427599 338085
rect 427541 338045 427553 338079
rect 427587 338076 427599 338079
rect 445478 338076 445484 338088
rect 427587 338048 445484 338076
rect 427587 338045 427599 338048
rect 427541 338039 427599 338045
rect 445478 338036 445484 338048
rect 445536 338036 445542 338088
rect 451461 338079 451519 338085
rect 451461 338045 451473 338079
rect 451507 338076 451519 338079
rect 451734 338076 451740 338088
rect 451507 338048 451740 338076
rect 451507 338045 451519 338048
rect 451461 338039 451519 338045
rect 451734 338036 451740 338048
rect 451792 338036 451798 338088
rect 490834 338036 490840 338088
rect 490892 338076 490898 338088
rect 498933 338079 498991 338085
rect 498933 338076 498945 338079
rect 490892 338048 498945 338076
rect 490892 338036 490898 338048
rect 498933 338045 498945 338048
rect 498979 338045 498991 338079
rect 498933 338039 498991 338045
rect 509142 338036 509148 338088
rect 509200 338076 509206 338088
rect 542354 338076 542360 338088
rect 509200 338048 542360 338076
rect 509200 338036 509206 338048
rect 542354 338036 542360 338048
rect 542412 338036 542418 338088
rect 66898 337968 66904 338020
rect 66956 338008 66962 338020
rect 261202 338008 261208 338020
rect 66956 337980 261208 338008
rect 66956 337968 66962 337980
rect 261202 337968 261208 337980
rect 261260 337968 261266 338020
rect 322750 337968 322756 338020
rect 322808 338008 322814 338020
rect 395246 338008 395252 338020
rect 322808 337980 395252 338008
rect 322808 337968 322814 337980
rect 395246 337968 395252 337980
rect 395304 337968 395310 338020
rect 402606 338008 402612 338020
rect 395356 337980 402612 338008
rect 3234 337900 3240 337952
rect 3292 337940 3298 337952
rect 6362 337940 6368 337952
rect 3292 337912 6368 337940
rect 3292 337900 3298 337912
rect 6362 337900 6368 337912
rect 6420 337900 6426 337952
rect 57238 337900 57244 337952
rect 57296 337940 57302 337952
rect 257522 337940 257528 337952
rect 57296 337912 257528 337940
rect 57296 337900 57302 337912
rect 257522 337900 257528 337912
rect 257580 337900 257586 337952
rect 309778 337900 309784 337952
rect 309836 337940 309842 337952
rect 309836 337912 315528 337940
rect 309836 337900 309842 337912
rect 50338 337832 50344 337884
rect 50396 337872 50402 337884
rect 251358 337872 251364 337884
rect 50396 337844 251364 337872
rect 50396 337832 50402 337844
rect 251358 337832 251364 337844
rect 251416 337832 251422 337884
rect 268378 337832 268384 337884
rect 268436 337872 268442 337884
rect 288710 337872 288716 337884
rect 268436 337844 288716 337872
rect 268436 337832 268442 337844
rect 288710 337832 288716 337844
rect 288768 337832 288774 337884
rect 311894 337832 311900 337884
rect 311952 337872 311958 337884
rect 312262 337872 312268 337884
rect 311952 337844 312268 337872
rect 311952 337832 311958 337844
rect 312262 337832 312268 337844
rect 312320 337832 312326 337884
rect 313458 337832 313464 337884
rect 313516 337872 313522 337884
rect 314102 337872 314108 337884
rect 313516 337844 314108 337872
rect 313516 337832 313522 337844
rect 314102 337832 314108 337844
rect 314160 337832 314166 337884
rect 314654 337832 314660 337884
rect 314712 337872 314718 337884
rect 315390 337872 315396 337884
rect 314712 337844 315396 337872
rect 314712 337832 314718 337844
rect 315390 337832 315396 337844
rect 315448 337832 315454 337884
rect 315500 337872 315528 337912
rect 316034 337900 316040 337952
rect 316092 337940 316098 337952
rect 316678 337940 316684 337952
rect 316092 337912 316684 337940
rect 316092 337900 316098 337912
rect 316678 337900 316684 337912
rect 316736 337900 316742 337952
rect 317598 337900 317604 337952
rect 317656 337940 317662 337952
rect 318334 337940 318340 337952
rect 317656 337912 318340 337940
rect 317656 337900 317662 337912
rect 318334 337900 318340 337912
rect 318392 337900 318398 337952
rect 320174 337900 320180 337952
rect 320232 337940 320238 337952
rect 320910 337940 320916 337952
rect 320232 337912 320916 337940
rect 320232 337900 320238 337912
rect 320910 337900 320916 337912
rect 320968 337900 320974 337952
rect 326341 337943 326399 337949
rect 326341 337909 326353 337943
rect 326387 337940 326399 337943
rect 384301 337943 384359 337949
rect 384301 337940 384313 337943
rect 326387 337912 384313 337940
rect 326387 337909 326399 337912
rect 326341 337903 326399 337909
rect 384301 337909 384313 337912
rect 384347 337909 384359 337943
rect 384301 337903 384359 337909
rect 385678 337900 385684 337952
rect 385736 337940 385742 337952
rect 389726 337940 389732 337952
rect 385736 337912 389732 337940
rect 385736 337900 385742 337912
rect 389726 337900 389732 337912
rect 389784 337900 389790 337952
rect 393869 337943 393927 337949
rect 393869 337909 393881 337943
rect 393915 337940 393927 337943
rect 395356 337940 395384 337980
rect 402606 337968 402612 337980
rect 402664 337968 402670 338020
rect 416682 337968 416688 338020
rect 416740 338008 416746 338020
rect 443638 338008 443644 338020
rect 416740 337980 443644 338008
rect 416740 337968 416746 337980
rect 443638 337968 443644 337980
rect 443696 337968 443702 338020
rect 450354 338008 450360 338020
rect 443748 337980 450360 338008
rect 393915 337912 395384 337940
rect 395433 337943 395491 337949
rect 393915 337909 393927 337912
rect 393869 337903 393927 337909
rect 395433 337909 395445 337943
rect 395479 337940 395491 337943
rect 398745 337943 398803 337949
rect 398745 337940 398757 337943
rect 395479 337912 398757 337940
rect 395479 337909 395491 337912
rect 395433 337903 395491 337909
rect 398745 337909 398757 337912
rect 398791 337909 398803 337943
rect 398745 337903 398803 337909
rect 407758 337900 407764 337952
rect 407816 337940 407822 337952
rect 415486 337940 415492 337952
rect 407816 337912 415492 337940
rect 407816 337900 407822 337912
rect 415486 337900 415492 337912
rect 415544 337900 415550 337952
rect 416038 337900 416044 337952
rect 416096 337940 416102 337952
rect 442994 337940 443000 337952
rect 416096 337912 443000 337940
rect 416096 337900 416102 337912
rect 442994 337900 443000 337912
rect 443052 337900 443058 337952
rect 387978 337872 387984 337884
rect 315500 337844 387984 337872
rect 387978 337832 387984 337844
rect 388036 337832 388042 337884
rect 391198 337832 391204 337884
rect 391256 337872 391262 337884
rect 397086 337872 397092 337884
rect 391256 337844 397092 337872
rect 391256 337832 391262 337844
rect 397086 337832 397092 337844
rect 397144 337832 397150 337884
rect 422941 337875 422999 337881
rect 422941 337841 422953 337875
rect 422987 337872 422999 337875
rect 441246 337872 441252 337884
rect 422987 337844 441252 337872
rect 422987 337841 422999 337844
rect 422941 337835 422999 337841
rect 441246 337832 441252 337844
rect 441304 337832 441310 337884
rect 442169 337875 442227 337881
rect 442169 337841 442181 337875
rect 442215 337872 442227 337875
rect 443748 337872 443776 337980
rect 450354 337968 450360 337980
rect 450412 337968 450418 338020
rect 451918 337968 451924 338020
rect 451976 338008 451982 338020
rect 459002 338008 459008 338020
rect 451976 337980 459008 338008
rect 451976 337968 451982 337980
rect 459002 337968 459008 337980
rect 459060 337968 459066 338020
rect 477310 337968 477316 338020
rect 477368 338008 477374 338020
rect 480254 338008 480260 338020
rect 477368 337980 480260 338008
rect 477368 337968 477374 337980
rect 480254 337968 480260 337980
rect 480312 337968 480318 338020
rect 498746 337968 498752 338020
rect 498804 338008 498810 338020
rect 499482 338008 499488 338020
rect 498804 337980 499488 338008
rect 498804 337968 498810 337980
rect 499482 337968 499488 337980
rect 499540 337968 499546 338020
rect 512822 337968 512828 338020
rect 512880 338008 512886 338020
rect 547138 338008 547144 338020
rect 512880 337980 547144 338008
rect 512880 337968 512886 337980
rect 547138 337968 547144 337980
rect 547196 337968 547202 338020
rect 490190 337900 490196 337952
rect 490248 337940 490254 337952
rect 501598 337940 501604 337952
rect 490248 337912 501604 337940
rect 490248 337900 490254 337912
rect 501598 337900 501604 337912
rect 501656 337900 501662 337952
rect 503438 337900 503444 337952
rect 503496 337940 503502 337952
rect 503622 337940 503628 337952
rect 503496 337912 503628 337940
rect 503496 337900 503502 337912
rect 503622 337900 503628 337912
rect 503680 337900 503686 337952
rect 512270 337900 512276 337952
rect 512328 337940 512334 337952
rect 547230 337940 547236 337952
rect 512328 337912 547236 337940
rect 512328 337900 512334 337912
rect 547230 337900 547236 337912
rect 547288 337900 547294 337952
rect 442215 337844 443776 337872
rect 444009 337875 444067 337881
rect 442215 337841 442227 337844
rect 442169 337835 442227 337841
rect 444009 337841 444021 337875
rect 444055 337872 444067 337875
rect 450998 337872 451004 337884
rect 444055 337844 451004 337872
rect 444055 337841 444067 337844
rect 444009 337835 444067 337841
rect 450998 337832 451004 337844
rect 451056 337832 451062 337884
rect 453298 337832 453304 337884
rect 453356 337872 453362 337884
rect 462038 337872 462044 337884
rect 453356 337844 462044 337872
rect 453356 337832 453362 337844
rect 462038 337832 462044 337844
rect 462096 337832 462102 337884
rect 463602 337832 463608 337884
rect 463660 337872 463666 337884
rect 468110 337872 468116 337884
rect 463660 337844 468116 337872
rect 463660 337832 463666 337844
rect 468110 337832 468116 337844
rect 468168 337832 468174 337884
rect 487154 337832 487160 337884
rect 487212 337872 487218 337884
rect 499758 337872 499764 337884
rect 487212 337844 499764 337872
rect 487212 337832 487218 337844
rect 499758 337832 499764 337844
rect 499816 337832 499822 337884
rect 501230 337832 501236 337884
rect 501288 337872 501294 337884
rect 501288 337844 513052 337872
rect 501288 337832 501294 337844
rect 46198 337764 46204 337816
rect 46256 337804 46262 337816
rect 247678 337804 247684 337816
rect 46256 337776 247684 337804
rect 46256 337764 46262 337776
rect 247678 337764 247684 337776
rect 247736 337764 247742 337816
rect 269758 337764 269764 337816
rect 269816 337804 269822 337816
rect 292390 337804 292396 337816
rect 269816 337776 292396 337804
rect 269816 337764 269822 337776
rect 292390 337764 292396 337776
rect 292448 337764 292454 337816
rect 294598 337764 294604 337816
rect 294656 337804 294662 337816
rect 375098 337804 375104 337816
rect 294656 337776 375104 337804
rect 294656 337764 294662 337776
rect 375098 337764 375104 337776
rect 375156 337764 375162 337816
rect 375282 337764 375288 337816
rect 375340 337804 375346 337816
rect 384209 337807 384267 337813
rect 384209 337804 384221 337807
rect 375340 337776 384221 337804
rect 375340 337764 375346 337776
rect 384209 337773 384221 337776
rect 384255 337773 384267 337807
rect 406286 337804 406292 337816
rect 384209 337767 384267 337773
rect 384316 337776 406292 337804
rect 39298 337696 39304 337748
rect 39356 337736 39362 337748
rect 234617 337739 234675 337745
rect 234617 337736 234629 337739
rect 39356 337708 234629 337736
rect 39356 337696 39362 337708
rect 234617 337705 234629 337708
rect 234663 337705 234675 337739
rect 234617 337699 234675 337705
rect 237469 337739 237527 337745
rect 237469 337705 237481 337739
rect 237515 337736 237527 337739
rect 240410 337736 240416 337748
rect 237515 337708 240416 337736
rect 237515 337705 237527 337708
rect 237469 337699 237527 337705
rect 240410 337696 240416 337708
rect 240468 337696 240474 337748
rect 248414 337696 248420 337748
rect 248472 337736 248478 337748
rect 249518 337736 249524 337748
rect 248472 337708 249524 337736
rect 248472 337696 248478 337708
rect 249518 337696 249524 337708
rect 249576 337696 249582 337748
rect 249978 337696 249984 337748
rect 250036 337736 250042 337748
rect 250806 337736 250812 337748
rect 250036 337708 250812 337736
rect 250036 337696 250042 337708
rect 250806 337696 250812 337708
rect 250864 337696 250870 337748
rect 258718 337696 258724 337748
rect 258776 337736 258782 337748
rect 266722 337736 266728 337748
rect 258776 337708 266728 337736
rect 258776 337696 258782 337708
rect 266722 337696 266728 337708
rect 266780 337696 266786 337748
rect 287698 337696 287704 337748
rect 287756 337736 287762 337748
rect 363233 337739 363291 337745
rect 363233 337736 363245 337739
rect 287756 337708 363245 337736
rect 287756 337696 287762 337708
rect 363233 337705 363245 337708
rect 363279 337705 363291 337739
rect 363233 337699 363291 337705
rect 363325 337739 363383 337745
rect 363325 337705 363337 337739
rect 363371 337736 363383 337739
rect 373258 337736 373264 337748
rect 363371 337708 373264 337736
rect 363371 337705 363383 337708
rect 363325 337699 363383 337705
rect 373258 337696 373264 337708
rect 373316 337696 373322 337748
rect 376018 337696 376024 337748
rect 376076 337736 376082 337748
rect 384316 337736 384344 337776
rect 406286 337764 406292 337776
rect 406344 337764 406350 337816
rect 409782 337764 409788 337816
rect 409840 337804 409846 337816
rect 439958 337804 439964 337816
rect 409840 337776 439964 337804
rect 409840 337764 409846 337776
rect 439958 337764 439964 337776
rect 440016 337764 440022 337816
rect 445018 337764 445024 337816
rect 445076 337804 445082 337816
rect 456518 337804 456524 337816
rect 445076 337776 456524 337804
rect 445076 337764 445082 337776
rect 456518 337764 456524 337776
rect 456576 337764 456582 337816
rect 464982 337764 464988 337816
rect 465040 337804 465046 337816
rect 468754 337804 468760 337816
rect 465040 337776 468760 337804
rect 465040 337764 465046 337776
rect 468754 337764 468760 337776
rect 468812 337764 468818 337816
rect 482830 337764 482836 337816
rect 482888 337804 482894 337816
rect 486329 337807 486387 337813
rect 486329 337804 486341 337807
rect 482888 337776 486341 337804
rect 482888 337764 482894 337776
rect 486329 337773 486341 337776
rect 486375 337773 486387 337807
rect 486329 337767 486387 337773
rect 497550 337764 497556 337816
rect 497608 337804 497614 337816
rect 509878 337804 509884 337816
rect 497608 337776 509884 337804
rect 497608 337764 497614 337776
rect 509878 337764 509884 337776
rect 509936 337764 509942 337816
rect 376076 337708 384344 337736
rect 384393 337739 384451 337745
rect 376076 337696 376082 337708
rect 384393 337705 384405 337739
rect 384439 337736 384451 337739
rect 409966 337736 409972 337748
rect 384439 337708 409972 337736
rect 384439 337705 384451 337708
rect 384393 337699 384451 337705
rect 409966 337696 409972 337708
rect 410024 337696 410030 337748
rect 412542 337696 412548 337748
rect 412600 337736 412606 337748
rect 441798 337736 441804 337748
rect 412600 337708 441804 337736
rect 412600 337696 412606 337708
rect 441798 337696 441804 337708
rect 441856 337696 441862 337748
rect 442350 337696 442356 337748
rect 442408 337736 442414 337748
rect 454678 337736 454684 337748
rect 442408 337708 454684 337736
rect 442408 337696 442414 337708
rect 454678 337696 454684 337708
rect 454736 337696 454742 337748
rect 456058 337696 456064 337748
rect 456116 337736 456122 337748
rect 463878 337736 463884 337748
rect 456116 337708 463884 337736
rect 456116 337696 456122 337708
rect 463878 337696 463884 337708
rect 463936 337696 463942 337748
rect 477954 337696 477960 337748
rect 478012 337736 478018 337748
rect 478782 337736 478788 337748
rect 478012 337708 478788 337736
rect 478012 337696 478018 337708
rect 478782 337696 478788 337708
rect 478840 337696 478846 337748
rect 479150 337696 479156 337748
rect 479208 337736 479214 337748
rect 479208 337708 480300 337736
rect 479208 337696 479214 337708
rect 32398 337628 32404 337680
rect 32456 337668 32462 337680
rect 239401 337671 239459 337677
rect 239401 337668 239413 337671
rect 32456 337640 239413 337668
rect 32456 337628 32462 337640
rect 239401 337637 239413 337640
rect 239447 337637 239459 337671
rect 239401 337631 239459 337637
rect 264330 337628 264336 337680
rect 264388 337668 264394 337680
rect 281442 337668 281448 337680
rect 264388 337640 281448 337668
rect 264388 337628 264394 337640
rect 281442 337628 281448 337640
rect 281500 337628 281506 337680
rect 283558 337628 283564 337680
rect 283616 337668 283622 337680
rect 365898 337668 365904 337680
rect 283616 337640 365904 337668
rect 283616 337628 283622 337640
rect 365898 337628 365904 337640
rect 365956 337628 365962 337680
rect 366910 337628 366916 337680
rect 366968 337668 366974 337680
rect 418522 337668 418528 337680
rect 366968 337640 418528 337668
rect 366968 337628 366974 337640
rect 418522 337628 418528 337640
rect 418580 337628 418586 337680
rect 420822 337628 420828 337680
rect 420880 337668 420886 337680
rect 446122 337668 446128 337680
rect 420880 337640 446128 337668
rect 420880 337628 420886 337640
rect 446122 337628 446128 337640
rect 446180 337628 446186 337680
rect 449250 337628 449256 337680
rect 449308 337668 449314 337680
rect 457162 337668 457168 337680
rect 449308 337640 457168 337668
rect 449308 337628 449314 337640
rect 457162 337628 457168 337640
rect 457220 337628 457226 337680
rect 466362 337628 466368 337680
rect 466420 337668 466426 337680
rect 469398 337668 469404 337680
rect 466420 337640 469404 337668
rect 466420 337628 466426 337640
rect 469398 337628 469404 337640
rect 469456 337628 469462 337680
rect 475470 337628 475476 337680
rect 475528 337668 475534 337680
rect 477586 337668 477592 337680
rect 475528 337640 477592 337668
rect 475528 337628 475534 337640
rect 477586 337628 477592 337640
rect 477644 337628 477650 337680
rect 480272 337668 480300 337708
rect 480346 337696 480352 337748
rect 480404 337736 480410 337748
rect 481542 337736 481548 337748
rect 480404 337708 481548 337736
rect 480404 337696 480410 337708
rect 481542 337696 481548 337708
rect 481600 337696 481606 337748
rect 488994 337696 489000 337748
rect 489052 337736 489058 337748
rect 489052 337708 499896 337736
rect 489052 337696 489058 337708
rect 480272 337640 483336 337668
rect 28258 337560 28264 337612
rect 28316 337600 28322 337612
rect 237469 337603 237527 337609
rect 237469 337600 237481 337603
rect 28316 337572 237481 337600
rect 28316 337560 28322 337572
rect 237469 337569 237481 337572
rect 237515 337569 237527 337603
rect 248322 337600 248328 337612
rect 237469 337563 237527 337569
rect 237576 337572 248328 337600
rect 17218 337492 17224 337544
rect 17276 337532 17282 337544
rect 228085 337535 228143 337541
rect 228085 337532 228097 337535
rect 17276 337504 228097 337532
rect 17276 337492 17282 337504
rect 228085 337501 228097 337504
rect 228131 337501 228143 337535
rect 228085 337495 228143 337501
rect 228174 337492 228180 337544
rect 228232 337532 228238 337544
rect 234890 337532 234896 337544
rect 228232 337504 234896 337532
rect 228232 337492 228238 337504
rect 234890 337492 234896 337504
rect 234948 337492 234954 337544
rect 234985 337535 235043 337541
rect 234985 337501 234997 337535
rect 235031 337532 235043 337535
rect 237576 337532 237604 337572
rect 248322 337560 248328 337572
rect 248380 337560 248386 337612
rect 289998 337600 290004 337612
rect 248432 337572 290004 337600
rect 235031 337504 237604 337532
rect 239401 337535 239459 337541
rect 235031 337501 235043 337504
rect 234985 337495 235043 337501
rect 239401 337501 239413 337535
rect 239447 337532 239459 337535
rect 244642 337532 244648 337544
rect 239447 337504 244648 337532
rect 239447 337501 239459 337504
rect 239401 337495 239459 337501
rect 244642 337492 244648 337504
rect 244700 337492 244706 337544
rect 246298 337492 246304 337544
rect 246356 337532 246362 337544
rect 248432 337532 248460 337572
rect 289998 337560 290004 337572
rect 290056 337560 290062 337612
rect 293862 337560 293868 337612
rect 293920 337600 293926 337612
rect 380618 337600 380624 337612
rect 293920 337572 380624 337600
rect 293920 337560 293926 337572
rect 380618 337560 380624 337572
rect 380676 337560 380682 337612
rect 384301 337603 384359 337609
rect 384301 337569 384313 337603
rect 384347 337600 384359 337603
rect 391566 337600 391572 337612
rect 384347 337572 391572 337600
rect 384347 337569 384359 337572
rect 384301 337563 384359 337569
rect 391566 337560 391572 337572
rect 391624 337560 391630 337612
rect 393130 337560 393136 337612
rect 393188 337600 393194 337612
rect 432046 337600 432052 337612
rect 393188 337572 432052 337600
rect 393188 337560 393194 337572
rect 432046 337560 432052 337572
rect 432104 337560 432110 337612
rect 432141 337603 432199 337609
rect 432141 337569 432153 337603
rect 432187 337600 432199 337603
rect 432187 337572 433564 337600
rect 432187 337569 432199 337572
rect 432141 337563 432199 337569
rect 246356 337504 248460 337532
rect 246356 337492 246362 337504
rect 262858 337492 262864 337544
rect 262916 337532 262922 337544
rect 267461 337535 267519 337541
rect 267461 337532 267473 337535
rect 262916 337504 267473 337532
rect 262916 337492 262922 337504
rect 267461 337501 267473 337504
rect 267507 337501 267519 337535
rect 267461 337495 267519 337501
rect 267553 337535 267611 337541
rect 267553 337501 267565 337535
rect 267599 337532 267611 337535
rect 285030 337532 285036 337544
rect 267599 337504 285036 337532
rect 267599 337501 267611 337504
rect 267553 337495 267611 337501
rect 285030 337492 285036 337504
rect 285088 337492 285094 337544
rect 286962 337492 286968 337544
rect 287020 337532 287026 337544
rect 376938 337532 376944 337544
rect 287020 337504 376944 337532
rect 287020 337492 287026 337504
rect 376938 337492 376944 337504
rect 376996 337492 377002 337544
rect 384022 337532 384028 337544
rect 377048 337504 384028 337532
rect 24118 337424 24124 337476
rect 24176 337464 24182 337476
rect 24176 337436 237236 337464
rect 24176 337424 24182 337436
rect 15838 337356 15844 337408
rect 15896 337396 15902 337408
rect 228174 337396 228180 337408
rect 15896 337368 228180 337396
rect 15896 337356 15902 337368
rect 228174 337356 228180 337368
rect 228232 337356 228238 337408
rect 228269 337399 228327 337405
rect 228269 337365 228281 337399
rect 228315 337396 228327 337399
rect 235442 337396 235448 337408
rect 228315 337368 235448 337396
rect 228315 337365 228327 337368
rect 228269 337359 228327 337365
rect 235442 337356 235448 337368
rect 235500 337356 235506 337408
rect 237208 337396 237236 337436
rect 261478 337424 261484 337476
rect 261536 337464 261542 337476
rect 261536 337436 264192 337464
rect 261536 337424 261542 337436
rect 239766 337396 239772 337408
rect 237208 337368 239772 337396
rect 239766 337356 239772 337368
rect 239824 337356 239830 337408
rect 257338 337356 257344 337408
rect 257396 337396 257402 337408
rect 263042 337396 263048 337408
rect 257396 337368 263048 337396
rect 257396 337356 257402 337368
rect 263042 337356 263048 337368
rect 263100 337356 263106 337408
rect 61378 337288 61384 337340
rect 61436 337328 61442 337340
rect 252002 337328 252008 337340
rect 61436 337300 252008 337328
rect 61436 337288 61442 337300
rect 252002 337288 252008 337300
rect 252060 337288 252066 337340
rect 255958 337288 255964 337340
rect 256016 337328 256022 337340
rect 259362 337328 259368 337340
rect 256016 337300 259368 337328
rect 256016 337288 256022 337300
rect 259362 337288 259368 337300
rect 259420 337288 259426 337340
rect 264164 337328 264192 337436
rect 264238 337424 264244 337476
rect 264296 337464 264302 337476
rect 279602 337464 279608 337476
rect 264296 337436 279608 337464
rect 264296 337424 264302 337436
rect 279602 337424 279608 337436
rect 279660 337424 279666 337476
rect 280062 337424 280068 337476
rect 280120 337464 280126 337476
rect 363325 337467 363383 337473
rect 363325 337464 363337 337467
rect 280120 337436 363337 337464
rect 280120 337424 280126 337436
rect 363325 337433 363337 337436
rect 363371 337433 363383 337467
rect 363325 337427 363383 337433
rect 363417 337467 363475 337473
rect 363417 337433 363429 337467
rect 363463 337464 363475 337467
rect 369578 337464 369584 337476
rect 363463 337436 369584 337464
rect 363463 337433 363475 337436
rect 363417 337427 363475 337433
rect 369578 337424 369584 337436
rect 369636 337424 369642 337476
rect 374549 337467 374607 337473
rect 374549 337433 374561 337467
rect 374595 337464 374607 337467
rect 377048 337464 377076 337504
rect 384022 337492 384028 337504
rect 384080 337492 384086 337544
rect 384393 337535 384451 337541
rect 384393 337532 384405 337535
rect 384132 337504 384405 337532
rect 381449 337467 381507 337473
rect 374595 337436 377076 337464
rect 379348 337436 379652 337464
rect 374595 337433 374607 337436
rect 374549 337427 374607 337433
rect 267461 337399 267519 337405
rect 267461 337365 267473 337399
rect 267507 337396 267519 337399
rect 275922 337396 275928 337408
rect 267507 337368 275928 337396
rect 267507 337365 267519 337368
rect 267461 337359 267519 337365
rect 275922 337356 275928 337368
rect 275980 337356 275986 337408
rect 276658 337356 276664 337408
rect 276716 337396 276722 337408
rect 371418 337396 371424 337408
rect 276716 337368 371424 337396
rect 276716 337356 276722 337368
rect 371418 337356 371424 337368
rect 371476 337356 371482 337408
rect 372522 337356 372528 337408
rect 372580 337396 372586 337408
rect 379348 337396 379376 337436
rect 372580 337368 379376 337396
rect 379624 337396 379652 337436
rect 381449 337433 381461 337467
rect 381495 337464 381507 337467
rect 384132 337464 384160 337504
rect 384393 337501 384405 337504
rect 384439 337501 384451 337535
rect 384393 337495 384451 337501
rect 389082 337492 389088 337544
rect 389140 337532 389146 337544
rect 389140 337504 422984 337532
rect 389140 337492 389146 337504
rect 381495 337436 384160 337464
rect 384209 337467 384267 337473
rect 381495 337433 381507 337436
rect 381449 337427 381507 337433
rect 384209 337433 384221 337467
rect 384255 337464 384267 337467
rect 412913 337467 412971 337473
rect 412913 337464 412925 337467
rect 384255 337436 412925 337464
rect 384255 337433 384267 337436
rect 384209 337427 384267 337433
rect 412913 337433 412925 337436
rect 412959 337433 412971 337467
rect 412913 337427 412971 337433
rect 413462 337424 413468 337476
rect 413520 337464 413526 337476
rect 420362 337464 420368 337476
rect 413520 337436 420368 337464
rect 413520 337424 413526 337436
rect 420362 337424 420368 337436
rect 420420 337424 420426 337476
rect 421006 337396 421012 337408
rect 379624 337368 421012 337396
rect 372580 337356 372586 337368
rect 421006 337356 421012 337368
rect 421064 337356 421070 337408
rect 422956 337396 422984 337504
rect 429102 337492 429108 337544
rect 429160 337532 429166 337544
rect 433429 337535 433487 337541
rect 433429 337532 433441 337535
rect 429160 337504 433441 337532
rect 429160 337492 429166 337504
rect 433429 337501 433441 337504
rect 433475 337501 433487 337535
rect 433536 337532 433564 337572
rect 434622 337560 434628 337612
rect 434680 337600 434686 337612
rect 452838 337600 452844 337612
rect 434680 337572 452844 337600
rect 434680 337560 434686 337572
rect 452838 337560 452844 337572
rect 452896 337560 452902 337612
rect 453942 337560 453948 337612
rect 454000 337600 454006 337612
rect 463234 337600 463240 337612
rect 454000 337572 463240 337600
rect 454000 337560 454006 337572
rect 463234 337560 463240 337572
rect 463292 337560 463298 337612
rect 478506 337560 478512 337612
rect 478564 337600 478570 337612
rect 483198 337600 483204 337612
rect 478564 337572 483204 337600
rect 478564 337560 478570 337572
rect 483198 337560 483204 337572
rect 483256 337560 483262 337612
rect 483308 337600 483336 337640
rect 483474 337628 483480 337680
rect 483532 337668 483538 337680
rect 484210 337668 484216 337680
rect 483532 337640 484216 337668
rect 483532 337628 483538 337640
rect 484210 337628 484216 337640
rect 484268 337628 484274 337680
rect 485866 337628 485872 337680
rect 485924 337668 485930 337680
rect 489178 337668 489184 337680
rect 485924 337640 489184 337668
rect 485924 337628 485930 337640
rect 489178 337628 489184 337640
rect 489236 337628 489242 337680
rect 491386 337628 491392 337680
rect 491444 337668 491450 337680
rect 492582 337668 492588 337680
rect 491444 337640 492588 337668
rect 491444 337628 491450 337640
rect 492582 337628 492588 337640
rect 492640 337628 492646 337680
rect 493226 337628 493232 337680
rect 493284 337668 493290 337680
rect 493962 337668 493968 337680
rect 493284 337640 493968 337668
rect 493284 337628 493290 337640
rect 493962 337628 493968 337640
rect 494020 337628 494026 337680
rect 495636 337640 496860 337668
rect 484578 337600 484584 337612
rect 483308 337572 484584 337600
rect 484578 337560 484584 337572
rect 484636 337560 484642 337612
rect 492674 337560 492680 337612
rect 492732 337600 492738 337612
rect 495636 337600 495664 337640
rect 492732 337572 495664 337600
rect 492732 337560 492738 337572
rect 495710 337560 495716 337612
rect 495768 337600 495774 337612
rect 496722 337600 496728 337612
rect 495768 337572 496728 337600
rect 495768 337560 495774 337572
rect 496722 337560 496728 337572
rect 496780 337560 496786 337612
rect 496832 337600 496860 337640
rect 496906 337628 496912 337680
rect 496964 337668 496970 337680
rect 498838 337668 498844 337680
rect 496964 337640 498844 337668
rect 496964 337628 496970 337640
rect 498838 337628 498844 337640
rect 498896 337628 498902 337680
rect 498933 337671 498991 337677
rect 498933 337637 498945 337671
rect 498979 337668 498991 337671
rect 499761 337671 499819 337677
rect 499761 337668 499773 337671
rect 498979 337640 499773 337668
rect 498979 337637 498991 337640
rect 498933 337631 498991 337637
rect 499761 337637 499773 337640
rect 499807 337637 499819 337671
rect 499868 337668 499896 337708
rect 499942 337696 499948 337748
rect 500000 337736 500006 337748
rect 500770 337736 500776 337748
rect 500000 337708 500776 337736
rect 500000 337696 500006 337708
rect 500770 337696 500776 337708
rect 500828 337696 500834 337748
rect 502610 337736 502616 337748
rect 500880 337708 502616 337736
rect 500880 337668 500908 337708
rect 502610 337696 502616 337708
rect 502668 337696 502674 337748
rect 504266 337696 504272 337748
rect 504324 337736 504330 337748
rect 505002 337736 505008 337748
rect 504324 337708 505008 337736
rect 504324 337696 504330 337708
rect 505002 337696 505008 337708
rect 505060 337696 505066 337748
rect 505462 337696 505468 337748
rect 505520 337736 505526 337748
rect 506382 337736 506388 337748
rect 505520 337708 506388 337736
rect 505520 337696 505526 337708
rect 506382 337696 506388 337708
rect 506440 337696 506446 337748
rect 506750 337696 506756 337748
rect 506808 337736 506814 337748
rect 507762 337736 507768 337748
rect 506808 337708 507768 337736
rect 506808 337696 506814 337708
rect 507762 337696 507768 337708
rect 507820 337696 507826 337748
rect 507946 337696 507952 337748
rect 508004 337736 508010 337748
rect 509142 337736 509148 337748
rect 508004 337708 509148 337736
rect 508004 337696 508010 337708
rect 509142 337696 509148 337708
rect 509200 337696 509206 337748
rect 510982 337696 510988 337748
rect 511040 337736 511046 337748
rect 511902 337736 511908 337748
rect 511040 337708 511908 337736
rect 511040 337696 511046 337708
rect 511902 337696 511908 337708
rect 511960 337696 511966 337748
rect 499868 337640 500908 337668
rect 499761 337631 499819 337637
rect 502426 337628 502432 337680
rect 502484 337668 502490 337680
rect 503530 337668 503536 337680
rect 502484 337640 503536 337668
rect 502484 337628 502490 337640
rect 503530 337628 503536 337640
rect 503588 337628 503594 337680
rect 513024 337668 513052 337844
rect 514662 337832 514668 337884
rect 514720 337872 514726 337884
rect 514720 337844 518756 337872
rect 514720 337832 514726 337844
rect 515858 337764 515864 337816
rect 515916 337804 515922 337816
rect 518728 337804 518756 337844
rect 520826 337832 520832 337884
rect 520884 337872 520890 337884
rect 556798 337872 556804 337884
rect 520884 337844 556804 337872
rect 520884 337832 520890 337844
rect 556798 337832 556804 337844
rect 556856 337832 556862 337884
rect 553394 337804 553400 337816
rect 515916 337776 518664 337804
rect 518728 337776 553400 337804
rect 515916 337764 515922 337776
rect 516502 337696 516508 337748
rect 516560 337736 516566 337748
rect 517422 337736 517428 337748
rect 516560 337708 517428 337736
rect 516560 337696 516566 337708
rect 517422 337696 517428 337708
rect 517480 337696 517486 337748
rect 518636 337736 518664 337776
rect 553394 337764 553400 337776
rect 553452 337764 553458 337816
rect 554866 337736 554872 337748
rect 518636 337708 554872 337736
rect 554866 337696 554872 337708
rect 554924 337696 554930 337748
rect 516778 337668 516784 337680
rect 513024 337640 516784 337668
rect 516778 337628 516784 337640
rect 516836 337628 516842 337680
rect 518342 337628 518348 337680
rect 518400 337668 518406 337680
rect 560294 337668 560300 337680
rect 518400 337640 560300 337668
rect 518400 337628 518406 337640
rect 560294 337628 560300 337640
rect 560352 337628 560358 337680
rect 510798 337600 510804 337612
rect 496832 337572 510804 337600
rect 510798 337560 510804 337572
rect 510856 337560 510862 337612
rect 517698 337560 517704 337612
rect 517756 337600 517762 337612
rect 518802 337600 518808 337612
rect 517756 337572 518808 337600
rect 517756 337560 517762 337572
rect 518802 337560 518808 337572
rect 518860 337560 518866 337612
rect 518986 337560 518992 337612
rect 519044 337600 519050 337612
rect 520090 337600 520096 337612
rect 519044 337572 520096 337600
rect 519044 337560 519050 337572
rect 520090 337560 520096 337572
rect 520148 337560 520154 337612
rect 522022 337560 522028 337612
rect 522080 337600 522086 337612
rect 526717 337603 526775 337609
rect 522080 337572 526668 337600
rect 522080 337560 522086 337572
rect 444009 337535 444067 337541
rect 444009 337532 444021 337535
rect 433536 337504 444021 337532
rect 433429 337495 433487 337501
rect 444009 337501 444021 337504
rect 444055 337501 444067 337535
rect 446674 337532 446680 337544
rect 444009 337495 444067 337501
rect 444116 337504 446680 337532
rect 423033 337467 423091 337473
rect 423033 337433 423045 337467
rect 423079 337464 423091 337467
rect 444116 337464 444144 337504
rect 446674 337492 446680 337504
rect 446732 337492 446738 337544
rect 451182 337492 451188 337544
rect 451240 337532 451246 337544
rect 461394 337532 461400 337544
rect 451240 337504 461400 337532
rect 451240 337492 451246 337504
rect 461394 337492 461400 337504
rect 461452 337492 461458 337544
rect 479794 337492 479800 337544
rect 479852 337532 479858 337544
rect 479852 337504 480944 337532
rect 479852 337492 479858 337504
rect 423079 337436 444144 337464
rect 423079 337433 423091 337436
rect 423033 337427 423091 337433
rect 446398 337424 446404 337476
rect 446456 337464 446462 337476
rect 458358 337464 458364 337476
rect 446456 337436 458364 337464
rect 446456 337424 446462 337436
rect 458358 337424 458364 337436
rect 458416 337424 458422 337476
rect 429562 337396 429568 337408
rect 422956 337368 429568 337396
rect 429562 337356 429568 337368
rect 429620 337356 429626 337408
rect 430482 337356 430488 337408
rect 430540 337396 430546 337408
rect 432141 337399 432199 337405
rect 432141 337396 432153 337399
rect 430540 337368 432153 337396
rect 430540 337356 430546 337368
rect 432141 337365 432153 337368
rect 432187 337365 432199 337399
rect 432141 337359 432199 337365
rect 432601 337399 432659 337405
rect 432601 337365 432613 337399
rect 432647 337396 432659 337399
rect 447318 337396 447324 337408
rect 432647 337368 447324 337396
rect 432647 337365 432659 337368
rect 432601 337359 432659 337365
rect 447318 337356 447324 337368
rect 447376 337356 447382 337408
rect 448422 337356 448428 337408
rect 448480 337396 448486 337408
rect 460198 337396 460204 337408
rect 448480 337368 460204 337396
rect 448480 337356 448486 337368
rect 460198 337356 460204 337368
rect 460256 337356 460262 337408
rect 460842 337356 460848 337408
rect 460900 337396 460906 337408
rect 466914 337396 466920 337408
rect 460900 337368 466920 337396
rect 460900 337356 460906 337368
rect 466914 337356 466920 337368
rect 466972 337356 466978 337408
rect 270402 337328 270408 337340
rect 264164 337300 270408 337328
rect 270402 337288 270408 337300
rect 270460 337288 270466 337340
rect 284938 337288 284944 337340
rect 284996 337328 285002 337340
rect 338942 337328 338948 337340
rect 284996 337300 338948 337328
rect 284996 337288 285002 337300
rect 338942 337288 338948 337300
rect 339000 337288 339006 337340
rect 355965 337331 356023 337337
rect 355965 337297 355977 337331
rect 356011 337328 356023 337331
rect 365714 337328 365720 337340
rect 356011 337300 365720 337328
rect 356011 337297 356023 337300
rect 355965 337291 356023 337297
rect 365714 337288 365720 337300
rect 365772 337288 365778 337340
rect 378502 337288 378508 337340
rect 378560 337328 378566 337340
rect 385037 337331 385095 337337
rect 385037 337328 385049 337331
rect 378560 337300 385049 337328
rect 378560 337288 378566 337300
rect 385037 337297 385049 337300
rect 385083 337297 385095 337331
rect 385037 337291 385095 337297
rect 398745 337331 398803 337337
rect 398745 337297 398757 337331
rect 398791 337328 398803 337331
rect 403894 337328 403900 337340
rect 398791 337300 403900 337328
rect 398791 337297 398803 337300
rect 398745 337291 398803 337297
rect 403894 337288 403900 337300
rect 403952 337288 403958 337340
rect 409138 337288 409144 337340
rect 409196 337328 409202 337340
rect 428366 337328 428372 337340
rect 409196 337300 428372 337328
rect 409196 337288 409202 337300
rect 428366 337288 428372 337300
rect 428424 337288 428430 337340
rect 428550 337288 428556 337340
rect 428608 337328 428614 337340
rect 433337 337331 433395 337337
rect 433337 337328 433349 337331
rect 428608 337300 433349 337328
rect 428608 337288 428614 337300
rect 433337 337297 433349 337300
rect 433383 337297 433395 337331
rect 433337 337291 433395 337297
rect 433429 337331 433487 337337
rect 433429 337297 433441 337331
rect 433475 337328 433487 337331
rect 442169 337331 442227 337337
rect 442169 337328 442181 337331
rect 433475 337300 442181 337328
rect 433475 337297 433487 337300
rect 433429 337291 433487 337297
rect 442169 337297 442181 337300
rect 442215 337297 442227 337331
rect 442169 337291 442227 337297
rect 442258 337288 442264 337340
rect 442316 337328 442322 337340
rect 449802 337328 449808 337340
rect 442316 337300 449808 337328
rect 442316 337288 442322 337300
rect 449802 337288 449808 337300
rect 449860 337288 449866 337340
rect 480916 337328 480944 337504
rect 481634 337492 481640 337544
rect 481692 337532 481698 337544
rect 482830 337532 482836 337544
rect 481692 337504 482836 337532
rect 481692 337492 481698 337504
rect 482830 337492 482836 337504
rect 482888 337492 482894 337544
rect 494514 337492 494520 337544
rect 494572 337532 494578 337544
rect 513558 337532 513564 337544
rect 494572 337504 513564 337532
rect 494572 337492 494578 337504
rect 513558 337492 513564 337504
rect 513616 337492 513622 337544
rect 513834 337492 513840 337544
rect 513892 337532 513898 337544
rect 523589 337535 523647 337541
rect 523589 337532 523601 337535
rect 513892 337504 523601 337532
rect 513892 337492 513898 337504
rect 523589 337501 523601 337504
rect 523635 337501 523647 337535
rect 526640 337532 526668 337572
rect 526717 337569 526729 337603
rect 526763 337600 526775 337603
rect 563146 337600 563152 337612
rect 526763 337572 563152 337600
rect 526763 337569 526775 337572
rect 526717 337563 526775 337569
rect 563146 337560 563152 337572
rect 563204 337560 563210 337612
rect 567194 337532 567200 337544
rect 526640 337504 567200 337532
rect 523589 337495 523647 337501
rect 567194 337492 567200 337504
rect 567252 337492 567258 337544
rect 480990 337424 480996 337476
rect 481048 337464 481054 337476
rect 485038 337464 485044 337476
rect 481048 337436 485044 337464
rect 481048 337424 481054 337436
rect 485038 337424 485044 337436
rect 485096 337424 485102 337476
rect 485314 337424 485320 337476
rect 485372 337464 485378 337476
rect 493318 337464 493324 337476
rect 485372 337436 493324 337464
rect 485372 337424 485378 337436
rect 493318 337424 493324 337436
rect 493376 337424 493382 337476
rect 496262 337424 496268 337476
rect 496320 337464 496326 337476
rect 517606 337464 517612 337476
rect 496320 337436 517612 337464
rect 496320 337424 496326 337436
rect 517606 337424 517612 337436
rect 517664 337424 517670 337476
rect 519538 337424 519544 337476
rect 519596 337464 519602 337476
rect 524049 337467 524107 337473
rect 524049 337464 524061 337467
rect 519596 337436 524061 337464
rect 519596 337424 519602 337436
rect 524049 337433 524061 337436
rect 524095 337433 524107 337467
rect 569218 337464 569224 337476
rect 524049 337427 524107 337433
rect 526824 337436 569224 337464
rect 484670 337356 484676 337408
rect 484728 337396 484734 337408
rect 485682 337396 485688 337408
rect 484728 337368 485688 337396
rect 484728 337356 484734 337368
rect 485682 337356 485688 337368
rect 485740 337356 485746 337408
rect 486329 337399 486387 337405
rect 486329 337365 486341 337399
rect 486375 337396 486387 337399
rect 491478 337396 491484 337408
rect 486375 337368 491484 337396
rect 486375 337365 486387 337368
rect 486329 337359 486387 337365
rect 491478 337356 491484 337368
rect 491536 337356 491542 337408
rect 498102 337356 498108 337408
rect 498160 337396 498166 337408
rect 520366 337396 520372 337408
rect 498160 337368 520372 337396
rect 498160 337356 498166 337368
rect 520366 337356 520372 337368
rect 520424 337356 520430 337408
rect 523218 337356 523224 337408
rect 523276 337396 523282 337408
rect 526824 337396 526852 337436
rect 569218 337424 569224 337436
rect 569276 337424 569282 337476
rect 523276 337368 526852 337396
rect 523276 337356 523282 337368
rect 526898 337356 526904 337408
rect 526956 337396 526962 337408
rect 571978 337396 571984 337408
rect 526956 337368 571984 337396
rect 526956 337356 526962 337368
rect 571978 337356 571984 337368
rect 572036 337356 572042 337408
rect 485958 337328 485964 337340
rect 480916 337300 485964 337328
rect 485958 337288 485964 337300
rect 486016 337288 486022 337340
rect 499761 337331 499819 337337
rect 499761 337297 499773 337331
rect 499807 337328 499819 337331
rect 506658 337328 506664 337340
rect 499807 337300 506664 337328
rect 499807 337297 499819 337300
rect 499761 337291 499819 337297
rect 506658 337288 506664 337300
rect 506716 337288 506722 337340
rect 517146 337288 517152 337340
rect 517204 337328 517210 337340
rect 549898 337328 549904 337340
rect 517204 337300 549904 337328
rect 517204 337288 517210 337300
rect 549898 337288 549904 337300
rect 549956 337288 549962 337340
rect 84838 337220 84844 337272
rect 84896 337260 84902 337272
rect 272242 337260 272248 337272
rect 84896 337232 272248 337260
rect 84896 337220 84902 337232
rect 272242 337220 272248 337232
rect 272300 337220 272306 337272
rect 283650 337220 283656 337272
rect 283708 337260 283714 337272
rect 337102 337260 337108 337272
rect 283708 337232 337108 337260
rect 283708 337220 283714 337232
rect 337102 337220 337108 337232
rect 337160 337220 337166 337272
rect 339402 337220 339408 337272
rect 339460 337260 339466 337272
rect 339460 337232 345704 337260
rect 339460 337220 339466 337232
rect 97258 337152 97264 337204
rect 97316 337192 97322 337204
rect 277762 337192 277768 337204
rect 97316 337164 277768 337192
rect 97316 337152 97322 337164
rect 277762 337152 277768 337164
rect 277820 337152 277826 337204
rect 316678 337152 316684 337204
rect 316736 337192 316742 337204
rect 326341 337195 326399 337201
rect 326341 337192 326353 337195
rect 316736 337164 326353 337192
rect 316736 337152 316742 337164
rect 326341 337161 326353 337164
rect 326387 337161 326399 337195
rect 345676 337192 345704 337232
rect 346302 337220 346308 337272
rect 346360 337260 346366 337272
rect 407482 337260 407488 337272
rect 346360 337232 407488 337260
rect 346360 337220 346366 337232
rect 407482 337220 407488 337232
rect 407540 337220 407546 337272
rect 408497 337263 408555 337269
rect 408497 337229 408509 337263
rect 408543 337260 408555 337263
rect 408543 337232 411300 337260
rect 408543 337229 408555 337232
rect 408497 337223 408555 337229
rect 345676 337164 347912 337192
rect 326341 337155 326399 337161
rect 104802 337084 104808 337136
rect 104860 337124 104866 337136
rect 283190 337124 283196 337136
rect 104860 337096 283196 337124
rect 104860 337084 104866 337096
rect 283190 337084 283196 337096
rect 283248 337084 283254 337136
rect 347884 337124 347912 337164
rect 353202 337152 353208 337204
rect 353260 337192 353266 337204
rect 411162 337192 411168 337204
rect 353260 337164 411168 337192
rect 353260 337152 353266 337164
rect 411162 337152 411168 337164
rect 411220 337152 411226 337204
rect 411272 337192 411300 337232
rect 413370 337220 413376 337272
rect 413428 337260 413434 337272
rect 413428 337232 421144 337260
rect 413428 337220 413434 337232
rect 417326 337192 417332 337204
rect 411272 337164 417332 337192
rect 417326 337152 417332 337164
rect 417384 337152 417390 337204
rect 417602 337152 417608 337204
rect 417660 337192 417666 337204
rect 421009 337195 421067 337201
rect 421009 337192 421021 337195
rect 417660 337164 421021 337192
rect 417660 337152 417666 337164
rect 421009 337161 421021 337164
rect 421055 337161 421067 337195
rect 421116 337192 421144 337232
rect 422202 337220 422208 337272
rect 422260 337260 422266 337272
rect 423033 337263 423091 337269
rect 423033 337260 423045 337263
rect 422260 337232 423045 337260
rect 422260 337220 422266 337232
rect 423033 337229 423045 337232
rect 423079 337229 423091 337263
rect 423033 337223 423091 337229
rect 424962 337220 424968 337272
rect 425020 337260 425026 337272
rect 447962 337260 447968 337272
rect 425020 337232 447968 337260
rect 425020 337220 425026 337232
rect 447962 337220 447968 337232
rect 448020 337220 448026 337272
rect 508590 337220 508596 337272
rect 508648 337260 508654 337272
rect 540238 337260 540244 337272
rect 508648 337232 540244 337260
rect 508648 337220 508654 337232
rect 540238 337220 540244 337232
rect 540296 337220 540302 337272
rect 424042 337192 424048 337204
rect 421116 337164 424048 337192
rect 421009 337155 421067 337161
rect 424042 337152 424048 337164
rect 424100 337152 424106 337204
rect 430485 337195 430543 337201
rect 430485 337161 430497 337195
rect 430531 337192 430543 337195
rect 433242 337192 433248 337204
rect 430531 337164 433248 337192
rect 430531 337161 430543 337164
rect 430485 337155 430543 337161
rect 433242 337152 433248 337164
rect 433300 337152 433306 337204
rect 433337 337195 433395 337201
rect 433337 337161 433349 337195
rect 433383 337192 433395 337195
rect 449158 337192 449164 337204
rect 433383 337164 449164 337192
rect 433383 337161 433395 337164
rect 433337 337155 433395 337161
rect 449158 337152 449164 337164
rect 449216 337152 449222 337204
rect 453390 337152 453396 337204
rect 453448 337192 453454 337204
rect 460750 337192 460756 337204
rect 453448 337164 460756 337192
rect 453448 337152 453454 337164
rect 460750 337152 460756 337164
rect 460808 337152 460814 337204
rect 515306 337152 515312 337204
rect 515364 337192 515370 337204
rect 523681 337195 523739 337201
rect 523681 337192 523693 337195
rect 515364 337164 523693 337192
rect 515364 337152 515370 337164
rect 523681 337161 523693 337164
rect 523727 337161 523739 337195
rect 523681 337155 523739 337161
rect 524049 337195 524107 337201
rect 524049 337161 524061 337195
rect 524095 337192 524107 337195
rect 526717 337195 526775 337201
rect 526717 337192 526729 337195
rect 524095 337164 526729 337192
rect 524095 337161 524107 337164
rect 524049 337155 524107 337161
rect 526717 337161 526729 337164
rect 526763 337161 526775 337195
rect 526717 337155 526775 337161
rect 526806 337152 526812 337204
rect 526864 337192 526870 337204
rect 528649 337195 528707 337201
rect 528649 337192 528661 337195
rect 526864 337164 528661 337192
rect 526864 337152 526870 337164
rect 528649 337161 528661 337164
rect 528695 337161 528707 337195
rect 528649 337155 528707 337161
rect 528738 337152 528744 337204
rect 528796 337192 528802 337204
rect 529750 337192 529756 337204
rect 528796 337164 529756 337192
rect 528796 337152 528802 337164
rect 529750 337152 529756 337164
rect 529808 337152 529814 337204
rect 529845 337195 529903 337201
rect 529845 337161 529857 337195
rect 529891 337192 529903 337195
rect 558178 337192 558184 337204
rect 529891 337164 558184 337192
rect 529891 337161 529903 337164
rect 529845 337155 529903 337161
rect 558178 337152 558184 337164
rect 558236 337152 558242 337204
rect 355965 337127 356023 337133
rect 355965 337124 355977 337127
rect 347884 337096 355977 337124
rect 355965 337093 355977 337096
rect 356011 337093 356023 337127
rect 355965 337087 356023 337093
rect 357342 337084 357348 337136
rect 357400 337124 357406 337136
rect 413646 337124 413652 337136
rect 357400 337096 413652 337124
rect 357400 337084 357406 337096
rect 413646 337084 413652 337096
rect 413704 337084 413710 337136
rect 414658 337084 414664 337136
rect 414716 337124 414722 337136
rect 422846 337124 422852 337136
rect 414716 337096 422852 337124
rect 414716 337084 414722 337096
rect 422846 337084 422852 337096
rect 422904 337084 422910 337136
rect 423582 337084 423588 337136
rect 423640 337124 423646 337136
rect 432601 337127 432659 337133
rect 432601 337124 432613 337127
rect 423640 337096 432613 337124
rect 423640 337084 423646 337096
rect 432601 337093 432613 337096
rect 432647 337093 432659 337127
rect 451642 337124 451648 337136
rect 432601 337087 432659 337093
rect 432800 337096 451648 337124
rect 111702 337016 111708 337068
rect 111760 337056 111766 337068
rect 286870 337056 286876 337068
rect 111760 337028 286876 337056
rect 111760 337016 111766 337028
rect 286870 337016 286876 337028
rect 286928 337016 286934 337068
rect 360102 337016 360108 337068
rect 360160 337056 360166 337068
rect 414842 337056 414848 337068
rect 360160 337028 414848 337056
rect 360160 337016 360166 337028
rect 414842 337016 414848 337028
rect 414900 337016 414906 337068
rect 420270 337016 420276 337068
rect 420328 337056 420334 337068
rect 430485 337059 430543 337065
rect 430485 337056 430497 337059
rect 420328 337028 430497 337056
rect 420328 337016 420334 337028
rect 430485 337025 430497 337028
rect 430531 337025 430543 337059
rect 430485 337019 430543 337025
rect 431862 337016 431868 337068
rect 431920 337056 431926 337068
rect 432800 337056 432828 337096
rect 451642 337084 451648 337096
rect 451700 337084 451706 337136
rect 507302 337084 507308 337136
rect 507360 337124 507366 337136
rect 538214 337124 538220 337136
rect 507360 337096 538220 337124
rect 507360 337084 507366 337096
rect 538214 337084 538220 337096
rect 538272 337084 538278 337136
rect 431920 337028 432828 337056
rect 432877 337059 432935 337065
rect 431920 337016 431926 337028
rect 432877 337025 432889 337059
rect 432923 337056 432935 337059
rect 435821 337059 435879 337065
rect 435821 337056 435833 337059
rect 432923 337028 435833 337056
rect 432923 337025 432935 337028
rect 432877 337019 432935 337025
rect 435821 337025 435833 337028
rect 435867 337025 435879 337059
rect 435821 337019 435879 337025
rect 436002 337016 436008 337068
rect 436060 337056 436066 337068
rect 454034 337056 454040 337068
rect 436060 337028 454040 337056
rect 436060 337016 436066 337028
rect 454034 337016 454040 337028
rect 454092 337016 454098 337068
rect 487706 337016 487712 337068
rect 487764 337056 487770 337068
rect 488442 337056 488448 337068
rect 487764 337028 488448 337056
rect 487764 337016 487770 337028
rect 488442 337016 488448 337028
rect 488500 337016 488506 337068
rect 495066 337016 495072 337068
rect 495124 337056 495130 337068
rect 496078 337056 496084 337068
rect 495124 337028 496084 337056
rect 495124 337016 495130 337028
rect 496078 337016 496084 337028
rect 496136 337016 496142 337068
rect 509786 337016 509792 337068
rect 509844 337056 509850 337068
rect 540330 337056 540336 337068
rect 509844 337028 540336 337056
rect 509844 337016 509850 337028
rect 540330 337016 540336 337028
rect 540388 337016 540394 337068
rect 118602 336948 118608 337000
rect 118660 336988 118666 337000
rect 290550 336988 290556 337000
rect 118660 336960 290556 336988
rect 118660 336948 118666 336960
rect 290550 336948 290556 336960
rect 290608 336948 290614 337000
rect 366358 336948 366364 337000
rect 366416 336988 366422 337000
rect 408497 336991 408555 336997
rect 408497 336988 408509 336991
rect 366416 336960 408509 336988
rect 366416 336948 366422 336960
rect 408497 336957 408509 336960
rect 408543 336957 408555 336991
rect 408497 336951 408555 336957
rect 410518 336948 410524 337000
rect 410576 336988 410582 337000
rect 416406 336988 416412 337000
rect 410576 336960 416412 336988
rect 410576 336948 410582 336960
rect 416406 336948 416412 336960
rect 416464 336948 416470 337000
rect 420178 336948 420184 337000
rect 420236 336988 420242 337000
rect 420236 336960 422064 336988
rect 420236 336948 420242 336960
rect 125502 336880 125508 336932
rect 125560 336920 125566 336932
rect 294230 336920 294236 336932
rect 125560 336892 294236 336920
rect 125560 336880 125566 336892
rect 294230 336880 294236 336892
rect 294288 336880 294294 336932
rect 363690 336880 363696 336932
rect 363748 336920 363754 336932
rect 363748 336892 394004 336920
rect 363748 336880 363754 336892
rect 105538 336812 105544 336864
rect 105596 336852 105602 336864
rect 274082 336852 274088 336864
rect 105596 336824 274088 336852
rect 105596 336812 105602 336824
rect 274082 336812 274088 336824
rect 274140 336812 274146 336864
rect 366450 336812 366456 336864
rect 366508 336852 366514 336864
rect 393869 336855 393927 336861
rect 393869 336852 393881 336855
rect 366508 336824 393881 336852
rect 366508 336812 366514 336824
rect 393869 336821 393881 336824
rect 393915 336821 393927 336855
rect 393976 336852 394004 336892
rect 395430 336880 395436 336932
rect 395488 336920 395494 336932
rect 400766 336920 400772 336932
rect 395488 336892 400772 336920
rect 395488 336880 395494 336892
rect 400766 336880 400772 336892
rect 400824 336880 400830 336932
rect 412913 336923 412971 336929
rect 412913 336889 412925 336923
rect 412959 336920 412971 336923
rect 421926 336920 421932 336932
rect 412959 336892 421932 336920
rect 412959 336889 412971 336892
rect 412913 336883 412971 336889
rect 421926 336880 421932 336892
rect 421984 336880 421990 336932
rect 422036 336920 422064 336960
rect 424410 336948 424416 337000
rect 424468 336988 424474 337000
rect 432509 336991 432567 336997
rect 432509 336988 432521 336991
rect 424468 336960 432521 336988
rect 424468 336948 424474 336960
rect 432509 336957 432521 336960
rect 432555 336957 432567 336991
rect 438762 336988 438768 337000
rect 432509 336951 432567 336957
rect 432616 336960 438768 336988
rect 422036 336892 424824 336920
rect 398926 336852 398932 336864
rect 393976 336824 398932 336852
rect 393869 336815 393927 336821
rect 398926 336812 398932 336824
rect 398984 336812 398990 336864
rect 404446 336852 404452 336864
rect 400876 336824 404452 336852
rect 106918 336744 106924 336796
rect 106976 336784 106982 336796
rect 268562 336784 268568 336796
rect 106976 336756 267044 336784
rect 106976 336744 106982 336756
rect 267016 336716 267044 336756
rect 267660 336756 268568 336784
rect 267660 336716 267688 336756
rect 268562 336744 268568 336756
rect 268620 336744 268626 336796
rect 363598 336744 363604 336796
rect 363656 336784 363662 336796
rect 374549 336787 374607 336793
rect 374549 336784 374561 336787
rect 363656 336756 374561 336784
rect 363656 336744 363662 336756
rect 374549 336753 374561 336756
rect 374595 336753 374607 336787
rect 374549 336747 374607 336753
rect 374638 336744 374644 336796
rect 374696 336784 374702 336796
rect 381449 336787 381507 336793
rect 381449 336784 381461 336787
rect 374696 336756 381461 336784
rect 374696 336744 374702 336756
rect 381449 336753 381461 336756
rect 381495 336753 381507 336787
rect 381449 336747 381507 336753
rect 381538 336744 381544 336796
rect 381596 336784 381602 336796
rect 382458 336784 382464 336796
rect 381596 336756 382464 336784
rect 381596 336744 381602 336756
rect 382458 336744 382464 336756
rect 382516 336744 382522 336796
rect 382918 336744 382924 336796
rect 382976 336784 382982 336796
rect 386138 336784 386144 336796
rect 382976 336756 386144 336784
rect 382976 336744 382982 336756
rect 386138 336744 386144 336756
rect 386196 336744 386202 336796
rect 389910 336744 389916 336796
rect 389968 336784 389974 336796
rect 393406 336784 393412 336796
rect 389968 336756 393412 336784
rect 389968 336744 389974 336756
rect 393406 336744 393412 336756
rect 393464 336744 393470 336796
rect 396718 336744 396724 336796
rect 396776 336784 396782 336796
rect 400876 336784 400904 336824
rect 404446 336812 404452 336824
rect 404504 336812 404510 336864
rect 413278 336812 413284 336864
rect 413336 336852 413342 336864
rect 422941 336855 422999 336861
rect 422941 336852 422953 336855
rect 413336 336824 422953 336852
rect 413336 336812 413342 336824
rect 422941 336821 422953 336824
rect 422987 336821 422999 336855
rect 424686 336852 424692 336864
rect 422941 336815 422999 336821
rect 423048 336824 424692 336852
rect 396776 336756 400904 336784
rect 396776 336744 396782 336756
rect 401042 336744 401048 336796
rect 401100 336784 401106 336796
rect 408126 336784 408132 336796
rect 401100 336756 408132 336784
rect 401100 336744 401106 336756
rect 408126 336744 408132 336756
rect 408184 336744 408190 336796
rect 410610 336744 410616 336796
rect 410668 336784 410674 336796
rect 413002 336784 413008 336796
rect 410668 336756 413008 336784
rect 410668 336744 410674 336756
rect 413002 336744 413008 336756
rect 413060 336744 413066 336796
rect 416130 336744 416136 336796
rect 416188 336784 416194 336796
rect 423048 336784 423076 336824
rect 424686 336812 424692 336824
rect 424744 336812 424750 336864
rect 424796 336852 424824 336892
rect 427078 336880 427084 336932
rect 427136 336920 427142 336932
rect 432616 336920 432644 336960
rect 438762 336948 438768 336960
rect 438820 336948 438826 337000
rect 503438 336948 503444 337000
rect 503496 336988 503502 337000
rect 514021 336991 514079 336997
rect 514021 336988 514033 336991
rect 503496 336960 514033 336988
rect 503496 336948 503502 336960
rect 514021 336957 514033 336960
rect 514067 336957 514079 336991
rect 514021 336951 514079 336957
rect 523681 336991 523739 336997
rect 523681 336957 523693 336991
rect 523727 336988 523739 336991
rect 545758 336988 545764 337000
rect 523727 336960 545764 336988
rect 523727 336957 523739 336960
rect 523681 336951 523739 336957
rect 545758 336948 545764 336960
rect 545816 336948 545822 337000
rect 440602 336920 440608 336932
rect 427136 336892 432644 336920
rect 432708 336892 440608 336920
rect 427136 336880 427142 336892
rect 427541 336855 427599 336861
rect 427541 336852 427553 336855
rect 424796 336824 427553 336852
rect 427541 336821 427553 336824
rect 427587 336821 427599 336855
rect 427541 336815 427599 336821
rect 431218 336812 431224 336864
rect 431276 336852 431282 336864
rect 432708 336852 432736 336892
rect 440602 336880 440608 336892
rect 440660 336880 440666 336932
rect 453482 336920 453488 336932
rect 447152 336892 453488 336920
rect 431276 336824 432736 336852
rect 431276 336812 431282 336824
rect 435358 336812 435364 336864
rect 435416 336852 435422 336864
rect 442442 336852 442448 336864
rect 435416 336824 442448 336852
rect 435416 336812 435422 336824
rect 442442 336812 442448 336824
rect 442500 336812 442506 336864
rect 416188 336756 423076 336784
rect 416188 336744 416194 336756
rect 424318 336744 424324 336796
rect 424376 336784 424382 336796
rect 425882 336784 425888 336796
rect 424376 336756 425888 336784
rect 424376 336744 424382 336756
rect 425882 336744 425888 336756
rect 425940 336744 425946 336796
rect 432598 336744 432604 336796
rect 432656 336784 432662 336796
rect 435726 336784 435732 336796
rect 432656 336756 435732 336784
rect 432656 336744 432662 336756
rect 435726 336744 435732 336756
rect 435784 336744 435790 336796
rect 435821 336787 435879 336793
rect 435821 336753 435833 336787
rect 435867 336784 435879 336787
rect 436922 336784 436928 336796
rect 435867 336756 436928 336784
rect 435867 336753 435879 336756
rect 435821 336747 435879 336753
rect 436922 336744 436928 336756
rect 436980 336744 436986 336796
rect 438118 336744 438124 336796
rect 438176 336784 438182 336796
rect 444282 336784 444288 336796
rect 438176 336756 444288 336784
rect 438176 336744 438182 336756
rect 444282 336744 444288 336756
rect 444340 336744 444346 336796
rect 446490 336744 446496 336796
rect 446548 336784 446554 336796
rect 447152 336784 447180 336892
rect 453482 336880 453488 336892
rect 453540 336880 453546 336932
rect 460198 336880 460204 336932
rect 460256 336920 460262 336932
rect 464430 336920 464436 336932
rect 460256 336892 464436 336920
rect 460256 336880 460262 336892
rect 464430 336880 464436 336892
rect 464488 336880 464494 336932
rect 476114 336880 476120 336932
rect 476172 336920 476178 336932
rect 477770 336920 477776 336932
rect 476172 336892 477776 336920
rect 476172 336880 476178 336892
rect 477770 336880 477776 336892
rect 477828 336880 477834 336932
rect 504910 336880 504916 336932
rect 504968 336920 504974 336932
rect 534074 336920 534080 336932
rect 504968 336892 534080 336920
rect 504968 336880 504974 336892
rect 534074 336880 534080 336892
rect 534132 336880 534138 336932
rect 464338 336812 464344 336864
rect 464396 336852 464402 336864
rect 466270 336852 466276 336864
rect 464396 336824 466276 336852
rect 464396 336812 464402 336824
rect 466270 336812 466276 336824
rect 466328 336812 466334 336864
rect 467742 336812 467748 336864
rect 467800 336852 467806 336864
rect 469950 336852 469956 336864
rect 467800 336824 469956 336852
rect 467800 336812 467806 336824
rect 469950 336812 469956 336824
rect 470008 336812 470014 336864
rect 523589 336855 523647 336861
rect 523589 336821 523601 336855
rect 523635 336852 523647 336855
rect 542998 336852 543004 336864
rect 523635 336824 543004 336852
rect 523635 336821 523647 336824
rect 523589 336815 523647 336821
rect 542998 336812 543004 336824
rect 543056 336812 543062 336864
rect 446548 336756 447180 336784
rect 446548 336744 446554 336756
rect 447778 336744 447784 336796
rect 447836 336784 447842 336796
rect 455322 336784 455328 336796
rect 447836 336756 455328 336784
rect 447836 336744 447842 336756
rect 455322 336744 455328 336756
rect 455380 336744 455386 336796
rect 457438 336744 457444 336796
rect 457496 336784 457502 336796
rect 462590 336784 462596 336796
rect 457496 336756 462596 336784
rect 457496 336744 457502 336756
rect 462590 336744 462596 336756
rect 462648 336744 462654 336796
rect 464430 336744 464436 336796
rect 464488 336784 464494 336796
rect 465718 336784 465724 336796
rect 464488 336756 465724 336784
rect 464488 336744 464494 336756
rect 465718 336744 465724 336756
rect 465776 336744 465782 336796
rect 469858 336744 469864 336796
rect 469916 336784 469922 336796
rect 471238 336784 471244 336796
rect 469916 336756 471244 336784
rect 469916 336744 469922 336756
rect 471238 336744 471244 336756
rect 471296 336744 471302 336796
rect 474918 336744 474924 336796
rect 474976 336784 474982 336796
rect 476022 336784 476028 336796
rect 474976 336756 476028 336784
rect 474976 336744 474982 336756
rect 476022 336744 476028 336756
rect 476080 336744 476086 336796
rect 514021 336787 514079 336793
rect 514021 336753 514033 336787
rect 514067 336784 514079 336787
rect 514067 336756 524460 336784
rect 514067 336753 514079 336756
rect 514021 336747 514079 336753
rect 267016 336688 267688 336716
rect 356517 336719 356575 336725
rect 356517 336685 356529 336719
rect 356563 336716 356575 336719
rect 356790 336716 356796 336728
rect 356563 336688 356796 336716
rect 356563 336685 356575 336688
rect 356517 336679 356575 336685
rect 356790 336676 356796 336688
rect 356848 336676 356854 336728
rect 370041 336719 370099 336725
rect 370041 336685 370053 336719
rect 370087 336716 370099 336719
rect 370498 336716 370504 336728
rect 370087 336688 370504 336716
rect 370087 336685 370099 336688
rect 370041 336679 370099 336685
rect 370498 336676 370504 336688
rect 370556 336676 370562 336728
rect 375561 336719 375619 336725
rect 375561 336685 375573 336719
rect 375607 336716 375619 336719
rect 375742 336716 375748 336728
rect 375607 336688 375748 336716
rect 375607 336685 375619 336688
rect 375561 336679 375619 336685
rect 375742 336676 375748 336688
rect 375800 336676 375806 336728
rect 380986 336676 380992 336728
rect 381044 336716 381050 336728
rect 381354 336716 381360 336728
rect 381044 336688 381360 336716
rect 381044 336676 381050 336688
rect 381354 336676 381360 336688
rect 381412 336676 381418 336728
rect 524432 336716 524460 336756
rect 524506 336744 524512 336796
rect 524564 336784 524570 336796
rect 525610 336784 525616 336796
rect 524564 336756 525616 336784
rect 524564 336744 524570 336756
rect 525610 336744 525616 336756
rect 525668 336744 525674 336796
rect 525720 336756 527496 336784
rect 525720 336716 525748 336756
rect 524432 336688 525748 336716
rect 527468 336716 527496 336756
rect 527542 336744 527548 336796
rect 527600 336784 527606 336796
rect 528462 336784 528468 336796
rect 527600 336756 528468 336784
rect 527600 336744 527606 336756
rect 528462 336744 528468 336756
rect 528520 336744 528526 336796
rect 528572 336756 529336 336784
rect 528572 336716 528600 336756
rect 527468 336688 528600 336716
rect 529308 336716 529336 336756
rect 529382 336744 529388 336796
rect 529440 336784 529446 336796
rect 529842 336784 529848 336796
rect 529440 336756 529848 336784
rect 529440 336744 529446 336756
rect 529842 336744 529848 336756
rect 529900 336744 529906 336796
rect 531314 336784 531320 336796
rect 529952 336756 531320 336784
rect 529952 336716 529980 336756
rect 531314 336744 531320 336756
rect 531372 336744 531378 336796
rect 529308 336688 529980 336716
rect 252554 336268 252560 336320
rect 252612 336308 252618 336320
rect 253842 336308 253848 336320
rect 252612 336280 253848 336308
rect 252612 336268 252618 336280
rect 253842 336268 253848 336280
rect 253900 336268 253906 336320
rect 229094 335588 229100 335640
rect 229152 335628 229158 335640
rect 229830 335628 229836 335640
rect 229152 335600 229836 335628
rect 229152 335588 229158 335600
rect 229830 335588 229836 335600
rect 229888 335588 229894 335640
rect 230474 335588 230480 335640
rect 230532 335628 230538 335640
rect 230934 335628 230940 335640
rect 230532 335600 230940 335628
rect 230532 335588 230538 335600
rect 230934 335588 230940 335600
rect 230992 335588 230998 335640
rect 241514 335588 241520 335640
rect 241572 335628 241578 335640
rect 241974 335628 241980 335640
rect 241572 335600 241980 335628
rect 241572 335588 241578 335600
rect 241974 335588 241980 335600
rect 242032 335588 242038 335640
rect 259638 335588 259644 335640
rect 259696 335628 259702 335640
rect 260282 335628 260288 335640
rect 259696 335600 260288 335628
rect 259696 335588 259702 335600
rect 260282 335588 260288 335600
rect 260340 335588 260346 335640
rect 296806 335588 296812 335640
rect 296864 335628 296870 335640
rect 297542 335628 297548 335640
rect 296864 335600 297548 335628
rect 296864 335588 296870 335600
rect 297542 335588 297548 335600
rect 297600 335588 297606 335640
rect 299474 335588 299480 335640
rect 299532 335628 299538 335640
rect 300118 335628 300124 335640
rect 299532 335600 300124 335628
rect 299532 335588 299538 335600
rect 300118 335588 300124 335600
rect 300176 335588 300182 335640
rect 302326 335588 302332 335640
rect 302384 335628 302390 335640
rect 303062 335628 303068 335640
rect 302384 335600 303068 335628
rect 302384 335588 302390 335600
rect 303062 335588 303068 335600
rect 303120 335588 303126 335640
rect 303614 335588 303620 335640
rect 303672 335628 303678 335640
rect 304350 335628 304356 335640
rect 303672 335600 304356 335628
rect 303672 335588 303678 335600
rect 304350 335588 304356 335600
rect 304408 335588 304414 335640
rect 306374 335588 306380 335640
rect 306432 335628 306438 335640
rect 306742 335628 306748 335640
rect 306432 335600 306748 335628
rect 306432 335588 306438 335600
rect 306742 335588 306748 335600
rect 306800 335588 306806 335640
rect 307846 335588 307852 335640
rect 307904 335628 307910 335640
rect 308030 335628 308036 335640
rect 307904 335600 308036 335628
rect 307904 335588 307910 335600
rect 308030 335588 308036 335600
rect 308088 335588 308094 335640
rect 310698 335588 310704 335640
rect 310756 335628 310762 335640
rect 311158 335628 311164 335640
rect 310756 335600 311164 335628
rect 310756 335588 310762 335600
rect 311158 335588 311164 335600
rect 311216 335588 311222 335640
rect 323118 335588 323124 335640
rect 323176 335628 323182 335640
rect 323854 335628 323860 335640
rect 323176 335600 323860 335628
rect 323176 335588 323182 335600
rect 323854 335588 323860 335600
rect 323912 335588 323918 335640
rect 328638 335588 328644 335640
rect 328696 335628 328702 335640
rect 329374 335628 329380 335640
rect 328696 335600 329380 335628
rect 328696 335588 328702 335600
rect 329374 335588 329380 335600
rect 329432 335588 329438 335640
rect 335354 335588 335360 335640
rect 335412 335628 335418 335640
rect 336182 335628 336188 335640
rect 335412 335600 336188 335628
rect 335412 335588 335418 335600
rect 336182 335588 336188 335600
rect 336240 335588 336246 335640
rect 339494 335588 339500 335640
rect 339552 335628 339558 335640
rect 340414 335628 340420 335640
rect 339552 335600 340420 335628
rect 339552 335588 339558 335600
rect 340414 335588 340420 335600
rect 340472 335588 340478 335640
rect 345014 335588 345020 335640
rect 345072 335628 345078 335640
rect 345934 335628 345940 335640
rect 345072 335600 345940 335628
rect 345072 335588 345078 335600
rect 345934 335588 345940 335600
rect 345992 335588 345998 335640
rect 350534 335588 350540 335640
rect 350592 335628 350598 335640
rect 351454 335628 351460 335640
rect 350592 335600 351460 335628
rect 350592 335588 350598 335600
rect 351454 335588 351460 335600
rect 351512 335588 351518 335640
rect 354674 335588 354680 335640
rect 354732 335628 354738 335640
rect 355134 335628 355140 335640
rect 354732 335600 355140 335628
rect 354732 335588 354738 335600
rect 355134 335588 355140 335600
rect 355192 335588 355198 335640
rect 357618 335588 357624 335640
rect 357676 335628 357682 335640
rect 358262 335628 358268 335640
rect 357676 335600 358268 335628
rect 357676 335588 357682 335600
rect 358262 335588 358268 335600
rect 358320 335588 358326 335640
rect 360194 335588 360200 335640
rect 360252 335628 360258 335640
rect 360654 335628 360660 335640
rect 360252 335600 360660 335628
rect 360252 335588 360258 335600
rect 360654 335588 360660 335600
rect 360712 335588 360718 335640
rect 361666 335588 361672 335640
rect 361724 335628 361730 335640
rect 362494 335628 362500 335640
rect 361724 335600 362500 335628
rect 361724 335588 361730 335600
rect 362494 335588 362500 335600
rect 362552 335588 362558 335640
rect 367186 335588 367192 335640
rect 367244 335628 367250 335640
rect 368014 335628 368020 335640
rect 367244 335600 368020 335628
rect 367244 335588 367250 335600
rect 368014 335588 368020 335600
rect 368072 335588 368078 335640
rect 378226 335588 378232 335640
rect 378284 335628 378290 335640
rect 379054 335628 379060 335640
rect 378284 335600 379060 335628
rect 378284 335588 378290 335600
rect 379054 335588 379060 335600
rect 379112 335588 379118 335640
rect 405918 335588 405924 335640
rect 405976 335628 405982 335640
rect 406654 335628 406660 335640
rect 405976 335600 406660 335628
rect 405976 335588 405982 335600
rect 406654 335588 406660 335600
rect 406712 335588 406718 335640
rect 422294 335588 422300 335640
rect 422352 335628 422358 335640
rect 423214 335628 423220 335640
rect 422352 335600 423220 335628
rect 422352 335588 422358 335600
rect 423214 335588 423220 335600
rect 423272 335588 423278 335640
rect 430574 335588 430580 335640
rect 430632 335628 430638 335640
rect 431126 335628 431132 335640
rect 430632 335600 431132 335628
rect 430632 335588 430638 335600
rect 431126 335588 431132 335600
rect 431184 335588 431190 335640
rect 470686 335588 470692 335640
rect 470744 335628 470750 335640
rect 471422 335628 471428 335640
rect 470744 335600 471428 335628
rect 470744 335588 470750 335600
rect 471422 335588 471428 335600
rect 471480 335588 471486 335640
rect 245654 335520 245660 335572
rect 245712 335560 245718 335572
rect 246482 335560 246488 335572
rect 245712 335532 246488 335560
rect 245712 335520 245718 335532
rect 246482 335520 246488 335532
rect 246540 335520 246546 335572
rect 334066 335384 334072 335436
rect 334124 335424 334130 335436
rect 334124 335396 334204 335424
rect 334124 335384 334130 335396
rect 334176 335232 334204 335396
rect 357618 335288 357624 335300
rect 357579 335260 357624 335288
rect 357618 335248 357624 335260
rect 357676 335248 357682 335300
rect 334158 335180 334164 335232
rect 334216 335180 334222 335232
rect 254118 335112 254124 335164
rect 254176 335152 254182 335164
rect 255038 335152 255044 335164
rect 254176 335124 255044 335152
rect 254176 335112 254182 335124
rect 255038 335112 255044 335124
rect 255096 335112 255102 335164
rect 340874 334568 340880 334620
rect 340932 334608 340938 334620
rect 341702 334608 341708 334620
rect 340932 334580 341708 334608
rect 340932 334568 340938 334580
rect 341702 334568 341708 334580
rect 341760 334568 341766 334620
rect 251818 334364 251824 334416
rect 251876 334404 251882 334416
rect 253198 334404 253204 334416
rect 251876 334376 253204 334404
rect 251876 334364 251882 334376
rect 253198 334364 253204 334376
rect 253256 334364 253262 334416
rect 362954 334364 362960 334416
rect 363012 334404 363018 334416
rect 363782 334404 363788 334416
rect 363012 334376 363788 334404
rect 363012 334364 363018 334376
rect 363782 334364 363788 334376
rect 363840 334364 363846 334416
rect 253198 334228 253204 334280
rect 253256 334268 253262 334280
rect 255682 334268 255688 334280
rect 253256 334240 255688 334268
rect 253256 334228 253262 334240
rect 255682 334228 255688 334240
rect 255740 334228 255746 334280
rect 294046 333928 294052 333940
rect 294007 333900 294052 333928
rect 294046 333888 294052 333900
rect 294104 333888 294110 333940
rect 237466 333616 237472 333668
rect 237524 333656 237530 333668
rect 238294 333656 238300 333668
rect 237524 333628 238300 333656
rect 237524 333616 237530 333628
rect 238294 333616 238300 333628
rect 238352 333616 238358 333668
rect 324406 333276 324412 333328
rect 324464 333316 324470 333328
rect 325050 333316 325056 333328
rect 324464 333288 325056 333316
rect 324464 333276 324470 333288
rect 325050 333276 325056 333288
rect 325108 333276 325114 333328
rect 433702 333276 433708 333328
rect 433760 333316 433766 333328
rect 434162 333316 434168 333328
rect 433760 333288 434168 333316
rect 433760 333276 433766 333288
rect 434162 333276 434168 333288
rect 434220 333276 434226 333328
rect 466546 333276 466552 333328
rect 466604 333316 466610 333328
rect 467098 333316 467104 333328
rect 466604 333288 467104 333316
rect 466604 333276 466610 333288
rect 467098 333276 467104 333288
rect 467156 333276 467162 333328
rect 325694 332732 325700 332784
rect 325752 332772 325758 332784
rect 326430 332772 326436 332784
rect 325752 332744 326436 332772
rect 325752 332732 325758 332744
rect 326430 332732 326436 332744
rect 326488 332732 326494 332784
rect 359090 331848 359096 331900
rect 359148 331888 359154 331900
rect 359274 331888 359280 331900
rect 359148 331860 359280 331888
rect 359148 331848 359154 331860
rect 359274 331848 359280 331860
rect 359332 331848 359338 331900
rect 349154 331780 349160 331832
rect 349212 331820 349218 331832
rect 349614 331820 349620 331832
rect 349212 331792 349620 331820
rect 349212 331780 349218 331792
rect 349614 331780 349620 331792
rect 349672 331780 349678 331832
rect 333974 331576 333980 331628
rect 334032 331616 334038 331628
rect 334250 331616 334256 331628
rect 334032 331588 334256 331616
rect 334032 331576 334038 331588
rect 334250 331576 334256 331588
rect 334308 331576 334314 331628
rect 343634 331508 343640 331560
rect 343692 331548 343698 331560
rect 344094 331548 344100 331560
rect 343692 331520 344100 331548
rect 343692 331508 343698 331520
rect 344094 331508 344100 331520
rect 344152 331508 344158 331560
rect 364518 331372 364524 331424
rect 364576 331412 364582 331424
rect 364978 331412 364984 331424
rect 364576 331384 364984 331412
rect 364576 331372 364582 331384
rect 364978 331372 364984 331384
rect 365036 331372 365042 331424
rect 231946 331236 231952 331288
rect 232004 331276 232010 331288
rect 232774 331276 232780 331288
rect 232004 331248 232780 331276
rect 232004 331236 232010 331248
rect 232774 331236 232780 331248
rect 232832 331236 232838 331288
rect 309413 331279 309471 331285
rect 309413 331245 309425 331279
rect 309459 331276 309471 331279
rect 309686 331276 309692 331288
rect 309459 331248 309692 331276
rect 309459 331245 309471 331248
rect 309413 331239 309471 331245
rect 309686 331236 309692 331248
rect 309744 331236 309750 331288
rect 342622 331276 342628 331288
rect 342583 331248 342628 331276
rect 342622 331236 342628 331248
rect 342680 331236 342686 331288
rect 393130 331276 393136 331288
rect 393091 331248 393136 331276
rect 393130 331236 393136 331248
rect 393188 331236 393194 331288
rect 305178 331168 305184 331220
rect 305236 331168 305242 331220
rect 416774 331168 416780 331220
rect 416832 331208 416838 331220
rect 416958 331208 416964 331220
rect 416832 331180 416964 331208
rect 416832 331168 416838 331180
rect 416958 331168 416964 331180
rect 417016 331168 417022 331220
rect 422294 331168 422300 331220
rect 422352 331208 422358 331220
rect 422478 331208 422484 331220
rect 422352 331180 422484 331208
rect 422352 331168 422358 331180
rect 422478 331168 422484 331180
rect 422536 331168 422542 331220
rect 305196 331140 305224 331168
rect 305270 331140 305276 331152
rect 305196 331112 305276 331140
rect 305270 331100 305276 331112
rect 305328 331100 305334 331152
rect 451461 330531 451519 330537
rect 451461 330497 451473 330531
rect 451507 330528 451519 330531
rect 451550 330528 451556 330540
rect 451507 330500 451556 330528
rect 451507 330497 451519 330500
rect 451461 330491 451519 330497
rect 451550 330488 451556 330500
rect 451608 330488 451614 330540
rect 292758 328992 292764 329044
rect 292816 329032 292822 329044
rect 293218 329032 293224 329044
rect 292816 329004 293224 329032
rect 292816 328992 292822 329004
rect 293218 328992 293224 329004
rect 293276 328992 293282 329044
rect 241790 328448 241796 328500
rect 241848 328488 241854 328500
rect 242434 328488 242440 328500
rect 241848 328460 242440 328488
rect 241848 328448 241854 328460
rect 242434 328448 242440 328460
rect 242492 328448 242498 328500
rect 265250 328448 265256 328500
rect 265308 328488 265314 328500
rect 265526 328488 265532 328500
rect 265308 328460 265532 328488
rect 265308 328448 265314 328460
rect 265526 328448 265532 328460
rect 265584 328448 265590 328500
rect 267090 328448 267096 328500
rect 267148 328488 267154 328500
rect 267553 328491 267611 328497
rect 267553 328488 267565 328491
rect 267148 328460 267565 328488
rect 267148 328448 267154 328460
rect 267553 328457 267565 328460
rect 267599 328457 267611 328491
rect 267553 328451 267611 328457
rect 270770 328448 270776 328500
rect 270828 328488 270834 328500
rect 271046 328488 271052 328500
rect 270828 328460 271052 328488
rect 270828 328448 270834 328460
rect 271046 328448 271052 328460
rect 271104 328448 271110 328500
rect 295610 328488 295616 328500
rect 295571 328460 295616 328488
rect 295610 328448 295616 328460
rect 295668 328448 295674 328500
rect 309410 328488 309416 328500
rect 309371 328460 309416 328488
rect 309410 328448 309416 328460
rect 309468 328448 309474 328500
rect 330018 328448 330024 328500
rect 330076 328488 330082 328500
rect 330570 328488 330576 328500
rect 330076 328460 330576 328488
rect 330076 328448 330082 328460
rect 330570 328448 330576 328460
rect 330628 328448 330634 328500
rect 331490 328448 331496 328500
rect 331548 328488 331554 328500
rect 331674 328488 331680 328500
rect 331548 328460 331680 328488
rect 331548 328448 331554 328460
rect 331674 328448 331680 328460
rect 331732 328448 331738 328500
rect 332686 328448 332692 328500
rect 332744 328488 332750 328500
rect 332962 328488 332968 328500
rect 332744 328460 332968 328488
rect 332744 328448 332750 328460
rect 332962 328448 332968 328460
rect 333020 328448 333026 328500
rect 334434 328448 334440 328500
rect 334492 328488 334498 328500
rect 334802 328488 334808 328500
rect 334492 328460 334808 328488
rect 334492 328448 334498 328460
rect 334802 328448 334808 328460
rect 334860 328448 334866 328500
rect 336918 328448 336924 328500
rect 336976 328488 336982 328500
rect 337194 328488 337200 328500
rect 336976 328460 337200 328488
rect 336976 328448 336982 328460
rect 337194 328448 337200 328460
rect 337252 328448 337258 328500
rect 342622 328488 342628 328500
rect 342583 328460 342628 328488
rect 342622 328448 342628 328460
rect 342680 328448 342686 328500
rect 397730 328448 397736 328500
rect 397788 328488 397794 328500
rect 397914 328488 397920 328500
rect 397788 328460 397920 328488
rect 397788 328448 397794 328460
rect 397914 328448 397920 328460
rect 397972 328448 397978 328500
rect 252646 328420 252652 328432
rect 252607 328392 252652 328420
rect 252646 328380 252652 328392
rect 252704 328380 252710 328432
rect 416869 328423 416927 328429
rect 416869 328389 416881 328423
rect 416915 328420 416927 328423
rect 416958 328420 416964 328432
rect 416915 328392 416964 328420
rect 416915 328389 416927 328392
rect 416869 328383 416927 328389
rect 416958 328380 416964 328392
rect 417016 328380 417022 328432
rect 422389 328423 422447 328429
rect 422389 328389 422401 328423
rect 422435 328420 422447 328423
rect 422478 328420 422484 328432
rect 422435 328392 422484 328420
rect 422435 328389 422447 328392
rect 422389 328383 422447 328389
rect 422478 328380 422484 328392
rect 422536 328380 422542 328432
rect 427909 328423 427967 328429
rect 427909 328389 427921 328423
rect 427955 328420 427967 328423
rect 427998 328420 428004 328432
rect 427955 328392 428004 328420
rect 427955 328389 427967 328392
rect 427909 328383 427967 328389
rect 427998 328380 428004 328392
rect 428056 328380 428062 328432
rect 433702 328420 433708 328432
rect 433663 328392 433708 328420
rect 433702 328380 433708 328392
rect 433760 328380 433766 328432
rect 472069 328423 472127 328429
rect 472069 328389 472081 328423
rect 472115 328420 472127 328423
rect 472158 328420 472164 328432
rect 472115 328392 472164 328420
rect 472115 328389 472127 328392
rect 472069 328383 472127 328389
rect 472158 328380 472164 328392
rect 472216 328380 472222 328432
rect 236270 327088 236276 327140
rect 236328 327128 236334 327140
rect 236914 327128 236920 327140
rect 236328 327100 236920 327128
rect 236328 327088 236334 327100
rect 236914 327088 236920 327100
rect 236972 327088 236978 327140
rect 370038 327128 370044 327140
rect 369999 327100 370044 327128
rect 370038 327088 370044 327100
rect 370096 327088 370102 327140
rect 375558 327128 375564 327140
rect 375519 327100 375564 327128
rect 375558 327088 375564 327100
rect 375616 327088 375622 327140
rect 393038 327088 393044 327140
rect 393096 327128 393102 327140
rect 393133 327131 393191 327137
rect 393133 327128 393145 327131
rect 393096 327100 393145 327128
rect 393096 327088 393102 327100
rect 393133 327097 393145 327100
rect 393179 327097 393191 327131
rect 393133 327091 393191 327097
rect 292758 327060 292764 327072
rect 292719 327032 292764 327060
rect 292758 327020 292764 327032
rect 292816 327020 292822 327072
rect 318978 326176 318984 326188
rect 318939 326148 318984 326176
rect 318978 326136 318984 326148
rect 319036 326136 319042 326188
rect 357618 325836 357624 325848
rect 357579 325808 357624 325836
rect 357618 325796 357624 325808
rect 357676 325796 357682 325848
rect 356514 325700 356520 325712
rect 356475 325672 356520 325700
rect 356514 325660 356520 325672
rect 356572 325660 356578 325712
rect 230658 325564 230664 325576
rect 230619 325536 230664 325564
rect 230658 325524 230664 325536
rect 230716 325524 230722 325576
rect 393038 324164 393044 324216
rect 393096 324204 393102 324216
rect 393225 324207 393283 324213
rect 393225 324204 393237 324207
rect 393096 324176 393237 324204
rect 393096 324164 393102 324176
rect 393225 324173 393237 324176
rect 393271 324173 393283 324207
rect 393225 324167 393283 324173
rect 2774 323552 2780 323604
rect 2832 323592 2838 323604
rect 5074 323592 5080 323604
rect 2832 323564 5080 323592
rect 2832 323552 2838 323564
rect 5074 323552 5080 323564
rect 5132 323552 5138 323604
rect 530854 322872 530860 322924
rect 530912 322912 530918 322924
rect 580074 322912 580080 322924
rect 530912 322884 580080 322912
rect 530912 322872 530918 322884
rect 580074 322872 580080 322884
rect 580132 322872 580138 322924
rect 249978 321688 249984 321700
rect 249939 321660 249984 321688
rect 249978 321648 249984 321660
rect 250036 321648 250042 321700
rect 261018 321648 261024 321700
rect 261076 321648 261082 321700
rect 231946 321580 231952 321632
rect 232004 321580 232010 321632
rect 259641 321623 259699 321629
rect 259641 321589 259653 321623
rect 259687 321620 259699 321623
rect 259730 321620 259736 321632
rect 259687 321592 259736 321620
rect 259687 321589 259699 321592
rect 259641 321583 259699 321589
rect 259730 321580 259736 321592
rect 259788 321580 259794 321632
rect 231964 321484 231992 321580
rect 261036 321564 261064 321648
rect 324498 321620 324504 321632
rect 324424 321592 324504 321620
rect 324424 321564 324452 321592
rect 324498 321580 324504 321592
rect 324556 321580 324562 321632
rect 359001 321623 359059 321629
rect 359001 321589 359013 321623
rect 359047 321620 359059 321623
rect 359090 321620 359096 321632
rect 359047 321592 359096 321620
rect 359047 321589 359059 321592
rect 359001 321583 359059 321589
rect 359090 321580 359096 321592
rect 359148 321580 359154 321632
rect 392121 321623 392179 321629
rect 392121 321589 392133 321623
rect 392167 321620 392179 321623
rect 392210 321620 392216 321632
rect 392167 321592 392216 321620
rect 392167 321589 392179 321592
rect 392121 321583 392179 321589
rect 392210 321580 392216 321592
rect 392268 321580 392274 321632
rect 408678 321580 408684 321632
rect 408736 321580 408742 321632
rect 466546 321620 466552 321632
rect 466507 321592 466552 321620
rect 466546 321580 466552 321592
rect 466604 321580 466610 321632
rect 261018 321512 261024 321564
rect 261076 321512 261082 321564
rect 324406 321512 324412 321564
rect 324464 321512 324470 321564
rect 400398 321512 400404 321564
rect 400456 321552 400462 321564
rect 400582 321552 400588 321564
rect 400456 321524 400588 321552
rect 400456 321512 400462 321524
rect 400582 321512 400588 321524
rect 400640 321512 400646 321564
rect 232038 321484 232044 321496
rect 231964 321456 232044 321484
rect 232038 321444 232044 321456
rect 232096 321444 232102 321496
rect 408696 321484 408724 321580
rect 408770 321484 408776 321496
rect 408696 321456 408776 321484
rect 408770 321444 408776 321456
rect 408828 321444 408834 321496
rect 252646 320124 252652 320136
rect 252607 320096 252652 320124
rect 252646 320084 252652 320096
rect 252704 320084 252710 320136
rect 230661 318835 230719 318841
rect 230661 318801 230673 318835
rect 230707 318832 230719 318835
rect 230842 318832 230848 318844
rect 230707 318804 230848 318832
rect 230707 318801 230719 318804
rect 230661 318795 230719 318801
rect 230842 318792 230848 318804
rect 230900 318792 230906 318844
rect 259638 318832 259644 318844
rect 259599 318804 259644 318832
rect 259638 318792 259644 318804
rect 259696 318792 259702 318844
rect 358998 318832 359004 318844
rect 358959 318804 359004 318832
rect 358998 318792 359004 318804
rect 359056 318792 359062 318844
rect 392118 318832 392124 318844
rect 392079 318804 392124 318832
rect 392118 318792 392124 318804
rect 392176 318792 392182 318844
rect 416866 318832 416872 318844
rect 416827 318804 416872 318832
rect 416866 318792 416872 318804
rect 416924 318792 416930 318844
rect 422386 318832 422392 318844
rect 422347 318804 422392 318832
rect 422386 318792 422392 318804
rect 422444 318792 422450 318844
rect 427906 318832 427912 318844
rect 427867 318804 427912 318832
rect 427906 318792 427912 318804
rect 427964 318792 427970 318844
rect 433705 318835 433763 318841
rect 433705 318801 433717 318835
rect 433751 318832 433763 318835
rect 433794 318832 433800 318844
rect 433751 318804 433800 318832
rect 433751 318801 433763 318804
rect 433705 318795 433763 318801
rect 433794 318792 433800 318804
rect 433852 318792 433858 318844
rect 466546 318832 466552 318844
rect 466507 318804 466552 318832
rect 466546 318792 466552 318804
rect 466604 318792 466610 318844
rect 472066 318832 472072 318844
rect 472027 318804 472072 318832
rect 472066 318792 472072 318804
rect 472124 318792 472130 318844
rect 283006 318724 283012 318776
rect 283064 318764 283070 318776
rect 283098 318764 283104 318776
rect 283064 318736 283104 318764
rect 283064 318724 283070 318736
rect 283098 318724 283104 318736
rect 283156 318724 283162 318776
rect 288618 318764 288624 318776
rect 288579 318736 288624 318764
rect 288618 318724 288624 318736
rect 288676 318724 288682 318776
rect 327258 318764 327264 318776
rect 327219 318736 327264 318764
rect 327258 318724 327264 318736
rect 327316 318724 327322 318776
rect 332778 318764 332784 318776
rect 332739 318736 332784 318764
rect 332778 318724 332784 318736
rect 332836 318724 332842 318776
rect 347958 318724 347964 318776
rect 348016 318764 348022 318776
rect 348050 318764 348056 318776
rect 348016 318736 348056 318764
rect 348016 318724 348022 318736
rect 348050 318724 348056 318736
rect 348108 318724 348114 318776
rect 352006 318724 352012 318776
rect 352064 318724 352070 318776
rect 353478 318724 353484 318776
rect 353536 318764 353542 318776
rect 353570 318764 353576 318776
rect 353536 318736 353576 318764
rect 353536 318724 353542 318736
rect 353570 318724 353576 318736
rect 353628 318724 353634 318776
rect 371329 318767 371387 318773
rect 371329 318733 371341 318767
rect 371375 318764 371387 318767
rect 371418 318764 371424 318776
rect 371375 318736 371424 318764
rect 371375 318733 371387 318736
rect 371329 318727 371387 318733
rect 371418 318724 371424 318736
rect 371476 318724 371482 318776
rect 375558 318724 375564 318776
rect 375616 318764 375622 318776
rect 375742 318764 375748 318776
rect 375616 318736 375748 318764
rect 375616 318724 375622 318736
rect 375742 318724 375748 318736
rect 375800 318724 375806 318776
rect 376849 318767 376907 318773
rect 376849 318733 376861 318767
rect 376895 318764 376907 318767
rect 376938 318764 376944 318776
rect 376895 318736 376944 318764
rect 376895 318733 376907 318736
rect 376849 318727 376907 318733
rect 376938 318724 376944 318736
rect 376996 318724 377002 318776
rect 381078 318724 381084 318776
rect 381136 318764 381142 318776
rect 381262 318764 381268 318776
rect 381136 318736 381268 318764
rect 381136 318724 381142 318736
rect 381262 318724 381268 318736
rect 381320 318724 381326 318776
rect 382274 318724 382280 318776
rect 382332 318764 382338 318776
rect 382458 318764 382464 318776
rect 382332 318736 382464 318764
rect 382332 318724 382338 318736
rect 382458 318724 382464 318736
rect 382516 318724 382522 318776
rect 387886 318724 387892 318776
rect 387944 318764 387950 318776
rect 387978 318764 387984 318776
rect 387944 318736 387984 318764
rect 387944 318724 387950 318736
rect 387978 318724 387984 318736
rect 388036 318724 388042 318776
rect 397730 318764 397736 318776
rect 397691 318736 397736 318764
rect 397730 318724 397736 318736
rect 397788 318724 397794 318776
rect 352024 318696 352052 318724
rect 352098 318696 352104 318708
rect 352024 318668 352104 318696
rect 352098 318656 352104 318668
rect 352156 318656 352162 318708
rect 249978 317472 249984 317484
rect 249939 317444 249984 317472
rect 249978 317432 249984 317444
rect 250036 317432 250042 317484
rect 292758 317472 292764 317484
rect 292719 317444 292764 317472
rect 292758 317432 292764 317444
rect 292816 317432 292822 317484
rect 318981 317475 319039 317481
rect 318981 317441 318993 317475
rect 319027 317472 319039 317475
rect 319162 317472 319168 317484
rect 319027 317444 319168 317472
rect 319027 317441 319039 317444
rect 318981 317435 319039 317441
rect 319162 317432 319168 317444
rect 319220 317432 319226 317484
rect 255406 317364 255412 317416
rect 255464 317404 255470 317416
rect 255590 317404 255596 317416
rect 255464 317376 255596 317404
rect 255464 317364 255470 317376
rect 255590 317364 255596 317376
rect 255648 317364 255654 317416
rect 283006 317364 283012 317416
rect 283064 317404 283070 317416
rect 283282 317404 283288 317416
rect 283064 317376 283288 317404
rect 283064 317364 283070 317376
rect 283282 317364 283288 317376
rect 283340 317364 283346 317416
rect 375742 317404 375748 317416
rect 375703 317376 375748 317404
rect 375742 317364 375748 317376
rect 375800 317364 375806 317416
rect 381262 317404 381268 317416
rect 381223 317376 381268 317404
rect 381262 317364 381268 317376
rect 381320 317364 381326 317416
rect 382274 317404 382280 317416
rect 382235 317376 382280 317404
rect 382274 317364 382280 317376
rect 382332 317364 382338 317416
rect 387886 317404 387892 317416
rect 387847 317376 387892 317404
rect 387886 317364 387892 317376
rect 387944 317364 387950 317416
rect 451550 316072 451556 316124
rect 451608 316112 451614 316124
rect 451734 316112 451740 316124
rect 451608 316084 451740 316112
rect 451608 316072 451614 316084
rect 451734 316072 451740 316084
rect 451792 316072 451798 316124
rect 277670 316004 277676 316056
rect 277728 316044 277734 316056
rect 277854 316044 277860 316056
rect 277728 316016 277860 316044
rect 277728 316004 277734 316016
rect 277854 316004 277860 316016
rect 277912 316004 277918 316056
rect 294049 316047 294107 316053
rect 294049 316013 294061 316047
rect 294095 316044 294107 316047
rect 294138 316044 294144 316056
rect 294095 316016 294144 316044
rect 294095 316013 294107 316016
rect 294049 316007 294107 316013
rect 294138 316004 294144 316016
rect 294196 316004 294202 316056
rect 357526 316004 357532 316056
rect 357584 316044 357590 316056
rect 357802 316044 357808 316056
rect 357584 316016 357808 316044
rect 357584 316004 357590 316016
rect 357802 316004 357808 316016
rect 357860 316004 357866 316056
rect 231949 315979 232007 315985
rect 231949 315945 231961 315979
rect 231995 315976 232007 315979
rect 232038 315976 232044 315988
rect 231995 315948 232044 315976
rect 231995 315945 232007 315948
rect 231949 315939 232007 315945
rect 232038 315936 232044 315948
rect 232096 315936 232102 315988
rect 356514 315976 356520 315988
rect 356475 315948 356520 315976
rect 356514 315936 356520 315948
rect 356572 315936 356578 315988
rect 451550 315976 451556 315988
rect 451511 315948 451556 315976
rect 451550 315936 451556 315948
rect 451608 315936 451614 315988
rect 397730 312168 397736 312180
rect 397691 312140 397736 312168
rect 397730 312128 397736 312140
rect 397788 312128 397794 312180
rect 294138 311924 294144 311976
rect 294196 311924 294202 311976
rect 230658 311856 230664 311908
rect 230716 311896 230722 311908
rect 230842 311896 230848 311908
rect 230716 311868 230848 311896
rect 230716 311856 230722 311868
rect 230842 311856 230848 311868
rect 230900 311856 230906 311908
rect 249978 311896 249984 311908
rect 249904 311868 249984 311896
rect 249904 311840 249932 311868
rect 249978 311856 249984 311868
rect 250036 311856 250042 311908
rect 277578 311896 277584 311908
rect 277539 311868 277584 311896
rect 277578 311856 277584 311868
rect 277636 311856 277642 311908
rect 294156 311840 294184 311924
rect 433426 311856 433432 311908
rect 433484 311896 433490 311908
rect 433794 311896 433800 311908
rect 433484 311868 433800 311896
rect 433484 311856 433490 311868
rect 433794 311856 433800 311868
rect 433852 311856 433858 311908
rect 249886 311788 249892 311840
rect 249944 311788 249950 311840
rect 294138 311788 294144 311840
rect 294196 311788 294202 311840
rect 346578 311828 346584 311840
rect 346539 311800 346584 311828
rect 346578 311788 346584 311800
rect 346636 311788 346642 311840
rect 416774 311788 416780 311840
rect 416832 311828 416838 311840
rect 416958 311828 416964 311840
rect 416832 311800 416964 311828
rect 416832 311788 416838 311800
rect 416958 311788 416964 311800
rect 417016 311788 417022 311840
rect 422294 311788 422300 311840
rect 422352 311828 422358 311840
rect 422478 311828 422484 311840
rect 422352 311800 422484 311828
rect 422352 311788 422358 311800
rect 422478 311788 422484 311800
rect 422536 311788 422542 311840
rect 427814 311788 427820 311840
rect 427872 311828 427878 311840
rect 427998 311828 428004 311840
rect 427872 311800 428004 311828
rect 427872 311788 427878 311800
rect 427998 311788 428004 311800
rect 428056 311788 428062 311840
rect 466454 311788 466460 311840
rect 466512 311828 466518 311840
rect 466638 311828 466644 311840
rect 466512 311800 466644 311828
rect 466512 311788 466518 311800
rect 466638 311788 466644 311800
rect 466696 311788 466702 311840
rect 471974 311788 471980 311840
rect 472032 311828 472038 311840
rect 472158 311828 472164 311840
rect 472032 311800 472164 311828
rect 472032 311788 472038 311800
rect 472158 311788 472164 311800
rect 472216 311788 472222 311840
rect 371326 309312 371332 309324
rect 371287 309284 371332 309312
rect 371326 309272 371332 309284
rect 371384 309272 371390 309324
rect 376846 309312 376852 309324
rect 376807 309284 376852 309312
rect 376846 309272 376852 309284
rect 376904 309272 376910 309324
rect 319162 309244 319168 309256
rect 318996 309216 319168 309244
rect 252554 309136 252560 309188
rect 252612 309176 252618 309188
rect 252738 309176 252744 309188
rect 252612 309148 252744 309176
rect 252612 309136 252618 309148
rect 252738 309136 252744 309148
rect 252796 309136 252802 309188
rect 267090 309176 267096 309188
rect 267051 309148 267096 309176
rect 267090 309136 267096 309148
rect 267148 309136 267154 309188
rect 287146 309136 287152 309188
rect 287204 309176 287210 309188
rect 287238 309176 287244 309188
rect 287204 309148 287244 309176
rect 287204 309136 287210 309148
rect 287238 309136 287244 309148
rect 287296 309136 287302 309188
rect 288618 309176 288624 309188
rect 288579 309148 288624 309176
rect 288618 309136 288624 309148
rect 288676 309136 288682 309188
rect 305178 309136 305184 309188
rect 305236 309176 305242 309188
rect 305270 309176 305276 309188
rect 305236 309148 305276 309176
rect 305236 309136 305242 309148
rect 305270 309136 305276 309148
rect 305328 309136 305334 309188
rect 318996 309120 319024 309216
rect 319162 309204 319168 309216
rect 319220 309204 319226 309256
rect 342622 309244 342628 309256
rect 342456 309216 342628 309244
rect 342456 309188 342484 309216
rect 342622 309204 342628 309216
rect 342680 309204 342686 309256
rect 324222 309136 324228 309188
rect 324280 309176 324286 309188
rect 324498 309176 324504 309188
rect 324280 309148 324504 309176
rect 324280 309136 324286 309148
rect 324498 309136 324504 309148
rect 324556 309136 324562 309188
rect 327258 309176 327264 309188
rect 327219 309148 327264 309176
rect 327258 309136 327264 309148
rect 327316 309136 327322 309188
rect 332778 309176 332784 309188
rect 332739 309148 332784 309176
rect 332778 309136 332784 309148
rect 332836 309136 332842 309188
rect 334434 309176 334440 309188
rect 334395 309148 334440 309176
rect 334434 309136 334440 309148
rect 334492 309136 334498 309188
rect 336826 309136 336832 309188
rect 336884 309176 336890 309188
rect 336918 309176 336924 309188
rect 336884 309148 336924 309176
rect 336884 309136 336890 309148
rect 336918 309136 336924 309148
rect 336976 309136 336982 309188
rect 342438 309136 342444 309188
rect 342496 309136 342502 309188
rect 346578 309176 346584 309188
rect 346539 309148 346584 309176
rect 346578 309136 346584 309148
rect 346636 309136 346642 309188
rect 393222 309176 393228 309188
rect 393183 309148 393228 309176
rect 393222 309136 393228 309148
rect 393280 309136 393286 309188
rect 400306 309136 400312 309188
rect 400364 309176 400370 309188
rect 400398 309176 400404 309188
rect 400364 309148 400404 309176
rect 400364 309136 400370 309148
rect 400398 309136 400404 309148
rect 400456 309136 400462 309188
rect 236270 309068 236276 309120
rect 236328 309108 236334 309120
rect 236362 309108 236368 309120
rect 236328 309080 236368 309108
rect 236328 309068 236334 309080
rect 236362 309068 236368 309080
rect 236420 309068 236426 309120
rect 270678 309108 270684 309120
rect 270639 309080 270684 309108
rect 270678 309068 270684 309080
rect 270736 309068 270742 309120
rect 309318 309108 309324 309120
rect 309279 309080 309324 309108
rect 309318 309068 309324 309080
rect 309376 309068 309382 309120
rect 318978 309068 318984 309120
rect 319036 309068 319042 309120
rect 375742 309108 375748 309120
rect 375703 309080 375748 309108
rect 375742 309068 375748 309080
rect 375800 309068 375806 309120
rect 376846 309108 376852 309120
rect 376807 309080 376852 309108
rect 376846 309068 376852 309080
rect 376904 309068 376910 309120
rect 416869 309111 416927 309117
rect 416869 309077 416881 309111
rect 416915 309108 416927 309111
rect 416958 309108 416964 309120
rect 416915 309080 416964 309108
rect 416915 309077 416927 309080
rect 416869 309071 416927 309077
rect 416958 309068 416964 309080
rect 417016 309068 417022 309120
rect 422478 309108 422484 309120
rect 422439 309080 422484 309108
rect 422478 309068 422484 309080
rect 422536 309068 422542 309120
rect 427998 309108 428004 309120
rect 427959 309080 428004 309108
rect 427998 309068 428004 309080
rect 428056 309068 428062 309120
rect 433426 309108 433432 309120
rect 433387 309080 433432 309108
rect 433426 309068 433432 309080
rect 433484 309068 433490 309120
rect 466549 309111 466607 309117
rect 466549 309077 466561 309111
rect 466595 309108 466607 309111
rect 466638 309108 466644 309120
rect 466595 309080 466644 309108
rect 466595 309077 466607 309080
rect 466549 309071 466607 309077
rect 466638 309068 466644 309080
rect 466696 309068 466702 309120
rect 472069 309111 472127 309117
rect 472069 309077 472081 309111
rect 472115 309108 472127 309111
rect 472158 309108 472164 309120
rect 472115 309080 472164 309108
rect 472115 309077 472127 309080
rect 472069 309071 472127 309077
rect 472158 309068 472164 309080
rect 472216 309068 472222 309120
rect 342438 309040 342444 309052
rect 342399 309012 342444 309040
rect 342438 309000 342444 309012
rect 342496 309000 342502 309052
rect 261018 307776 261024 307828
rect 261076 307816 261082 307828
rect 261110 307816 261116 307828
rect 261076 307788 261116 307816
rect 261076 307776 261082 307788
rect 261110 307776 261116 307788
rect 261168 307776 261174 307828
rect 267090 307816 267096 307828
rect 267051 307788 267096 307816
rect 267090 307776 267096 307788
rect 267148 307776 267154 307828
rect 334434 307816 334440 307828
rect 334395 307788 334440 307816
rect 334434 307776 334440 307788
rect 334492 307776 334498 307828
rect 381262 307816 381268 307828
rect 381223 307788 381268 307816
rect 381262 307776 381268 307788
rect 381320 307776 381326 307828
rect 387886 307816 387892 307828
rect 387847 307788 387892 307816
rect 387886 307776 387892 307788
rect 387944 307776 387950 307828
rect 242989 307751 243047 307757
rect 242989 307717 243001 307751
rect 243035 307748 243047 307751
rect 243078 307748 243084 307760
rect 243035 307720 243084 307748
rect 243035 307717 243047 307720
rect 242989 307711 243047 307717
rect 243078 307708 243084 307720
rect 243136 307708 243142 307760
rect 292758 307748 292764 307760
rect 292719 307720 292764 307748
rect 292758 307708 292764 307720
rect 292816 307708 292822 307760
rect 277578 306388 277584 306400
rect 277539 306360 277584 306388
rect 277578 306348 277584 306360
rect 277636 306348 277642 306400
rect 357526 306348 357532 306400
rect 357584 306388 357590 306400
rect 357618 306388 357624 306400
rect 357584 306360 357624 306388
rect 357584 306348 357590 306360
rect 357618 306348 357624 306360
rect 357676 306348 357682 306400
rect 365806 306348 365812 306400
rect 365864 306388 365870 306400
rect 365990 306388 365996 306400
rect 365864 306360 365996 306388
rect 365864 306348 365870 306360
rect 365990 306348 365996 306360
rect 366048 306348 366054 306400
rect 387886 304892 387892 304904
rect 387847 304864 387892 304892
rect 387886 304852 387892 304864
rect 387944 304852 387950 304904
rect 230658 304280 230664 304292
rect 230619 304252 230664 304280
rect 230658 304240 230664 304252
rect 230716 304240 230722 304292
rect 298278 302268 298284 302320
rect 298336 302268 298342 302320
rect 347958 302268 347964 302320
rect 348016 302268 348022 302320
rect 400398 302268 400404 302320
rect 400456 302268 400462 302320
rect 298296 302104 298324 302268
rect 347976 302184 348004 302268
rect 347958 302132 347964 302184
rect 348016 302132 348022 302184
rect 298370 302104 298376 302116
rect 298296 302076 298376 302104
rect 298370 302064 298376 302076
rect 298428 302064 298434 302116
rect 382277 302107 382335 302113
rect 382277 302073 382289 302107
rect 382323 302104 382335 302107
rect 382458 302104 382464 302116
rect 382323 302076 382464 302104
rect 382323 302073 382335 302076
rect 382277 302067 382335 302073
rect 382458 302064 382464 302076
rect 382516 302064 382522 302116
rect 400416 302104 400444 302268
rect 408770 302240 408776 302252
rect 408731 302212 408776 302240
rect 408770 302200 408776 302212
rect 408828 302200 408834 302252
rect 400490 302104 400496 302116
rect 400416 302076 400496 302104
rect 400490 302064 400496 302076
rect 400548 302064 400554 302116
rect 451550 302104 451556 302116
rect 451511 302076 451556 302104
rect 451550 302064 451556 302076
rect 451608 302064 451614 302116
rect 422478 299928 422484 299940
rect 422439 299900 422484 299928
rect 422478 299888 422484 299900
rect 422536 299888 422542 299940
rect 277578 299548 277584 299600
rect 277636 299548 277642 299600
rect 342441 299591 342499 299597
rect 342441 299557 342453 299591
rect 342487 299588 342499 299591
rect 342530 299588 342536 299600
rect 342487 299560 342536 299588
rect 342487 299557 342499 299560
rect 342441 299551 342499 299557
rect 342530 299548 342536 299560
rect 342588 299548 342594 299600
rect 230661 299523 230719 299529
rect 230661 299489 230673 299523
rect 230707 299520 230719 299523
rect 230842 299520 230848 299532
rect 230707 299492 230848 299520
rect 230707 299489 230719 299492
rect 230661 299483 230719 299489
rect 230842 299480 230848 299492
rect 230900 299480 230906 299532
rect 265158 299480 265164 299532
rect 265216 299520 265222 299532
rect 265250 299520 265256 299532
rect 265216 299492 265256 299520
rect 265216 299480 265222 299492
rect 265250 299480 265256 299492
rect 265308 299480 265314 299532
rect 270681 299523 270739 299529
rect 270681 299489 270693 299523
rect 270727 299520 270739 299523
rect 270770 299520 270776 299532
rect 270727 299492 270776 299520
rect 270727 299489 270739 299492
rect 270681 299483 270739 299489
rect 270770 299480 270776 299492
rect 270828 299480 270834 299532
rect 277596 299464 277624 299548
rect 309321 299523 309379 299529
rect 309321 299489 309333 299523
rect 309367 299520 309379 299523
rect 309410 299520 309416 299532
rect 309367 299492 309416 299520
rect 309367 299489 309379 299492
rect 309321 299483 309379 299489
rect 309410 299480 309416 299492
rect 309468 299480 309474 299532
rect 370130 299480 370136 299532
rect 370188 299520 370194 299532
rect 370222 299520 370228 299532
rect 370188 299492 370228 299520
rect 370188 299480 370194 299492
rect 370222 299480 370228 299492
rect 370280 299480 370286 299532
rect 375650 299480 375656 299532
rect 375708 299520 375714 299532
rect 375742 299520 375748 299532
rect 375708 299492 375748 299520
rect 375708 299480 375714 299492
rect 375742 299480 375748 299492
rect 375800 299480 375806 299532
rect 376849 299523 376907 299529
rect 376849 299489 376861 299523
rect 376895 299520 376907 299523
rect 376938 299520 376944 299532
rect 376895 299492 376944 299520
rect 376895 299489 376907 299492
rect 376849 299483 376907 299489
rect 376938 299480 376944 299492
rect 376996 299480 377002 299532
rect 416866 299520 416872 299532
rect 416827 299492 416872 299520
rect 416866 299480 416872 299492
rect 416924 299480 416930 299532
rect 427998 299520 428004 299532
rect 427959 299492 428004 299520
rect 427998 299480 428004 299492
rect 428056 299480 428062 299532
rect 433429 299523 433487 299529
rect 433429 299489 433441 299523
rect 433475 299520 433487 299523
rect 433702 299520 433708 299532
rect 433475 299492 433708 299520
rect 433475 299489 433487 299492
rect 433429 299483 433487 299489
rect 433702 299480 433708 299492
rect 433760 299480 433766 299532
rect 466546 299520 466552 299532
rect 466507 299492 466552 299520
rect 466546 299480 466552 299492
rect 466604 299480 466610 299532
rect 472066 299520 472072 299532
rect 472027 299492 472072 299520
rect 472066 299480 472072 299492
rect 472124 299480 472130 299532
rect 241790 299452 241796 299464
rect 241751 299424 241796 299452
rect 241790 299412 241796 299424
rect 241848 299412 241854 299464
rect 277578 299412 277584 299464
rect 277636 299412 277642 299464
rect 281629 299455 281687 299461
rect 281629 299421 281641 299455
rect 281675 299452 281687 299455
rect 281810 299452 281816 299464
rect 281675 299424 281816 299452
rect 281675 299421 281687 299424
rect 281629 299415 281687 299421
rect 281810 299412 281816 299424
rect 281868 299412 281874 299464
rect 305178 299452 305184 299464
rect 305139 299424 305184 299452
rect 305178 299412 305184 299424
rect 305236 299412 305242 299464
rect 310698 299452 310704 299464
rect 310659 299424 310704 299452
rect 310698 299412 310704 299424
rect 310756 299412 310762 299464
rect 331398 299412 331404 299464
rect 331456 299452 331462 299464
rect 331490 299452 331496 299464
rect 331456 299424 331496 299452
rect 331456 299412 331462 299424
rect 331490 299412 331496 299424
rect 331548 299412 331554 299464
rect 334250 299412 334256 299464
rect 334308 299452 334314 299464
rect 334434 299452 334440 299464
rect 334308 299424 334440 299452
rect 334308 299412 334314 299424
rect 334434 299412 334440 299424
rect 334492 299412 334498 299464
rect 346578 299452 346584 299464
rect 346539 299424 346584 299452
rect 346578 299412 346584 299424
rect 346636 299412 346642 299464
rect 382458 299452 382464 299464
rect 382419 299424 382464 299452
rect 382458 299412 382464 299424
rect 382516 299412 382522 299464
rect 324498 299384 324504 299396
rect 324459 299356 324504 299384
rect 324498 299344 324504 299356
rect 324556 299344 324562 299396
rect 292758 298228 292764 298240
rect 292719 298200 292764 298228
rect 292758 298188 292764 298200
rect 292816 298188 292822 298240
rect 231949 298163 232007 298169
rect 231949 298129 231961 298163
rect 231995 298160 232007 298163
rect 232038 298160 232044 298172
rect 231995 298132 232044 298160
rect 231995 298129 232007 298132
rect 231949 298123 232007 298129
rect 232038 298120 232044 298132
rect 232096 298120 232102 298172
rect 242986 298160 242992 298172
rect 242947 298132 242992 298160
rect 242986 298120 242992 298132
rect 243044 298120 243050 298172
rect 261018 298120 261024 298172
rect 261076 298160 261082 298172
rect 261202 298160 261208 298172
rect 261076 298132 261208 298160
rect 261076 298120 261082 298132
rect 261202 298120 261208 298132
rect 261260 298120 261266 298172
rect 356517 298163 356575 298169
rect 356517 298129 356529 298163
rect 356563 298160 356575 298163
rect 356606 298160 356612 298172
rect 356563 298132 356612 298160
rect 356563 298129 356575 298132
rect 356517 298123 356575 298129
rect 356606 298120 356612 298132
rect 356664 298120 356670 298172
rect 371234 298120 371240 298172
rect 371292 298160 371298 298172
rect 371602 298160 371608 298172
rect 371292 298132 371608 298160
rect 371292 298120 371298 298132
rect 371602 298120 371608 298132
rect 371660 298120 371666 298172
rect 387889 298163 387947 298169
rect 387889 298129 387901 298163
rect 387935 298160 387947 298163
rect 387978 298160 387984 298172
rect 387935 298132 387984 298160
rect 387935 298129 387947 298132
rect 387889 298123 387947 298129
rect 387978 298120 387984 298132
rect 388036 298120 388042 298172
rect 408770 298160 408776 298172
rect 408731 298132 408776 298160
rect 408770 298120 408776 298132
rect 408828 298120 408834 298172
rect 236270 298092 236276 298104
rect 236231 298064 236276 298092
rect 236270 298052 236276 298064
rect 236328 298052 236334 298104
rect 249886 298092 249892 298104
rect 249847 298064 249892 298092
rect 249886 298052 249892 298064
rect 249944 298052 249950 298104
rect 254210 298052 254216 298104
rect 254268 298092 254274 298104
rect 254486 298092 254492 298104
rect 254268 298064 254492 298092
rect 254268 298052 254274 298064
rect 254486 298052 254492 298064
rect 254544 298052 254550 298104
rect 255498 298092 255504 298104
rect 255459 298064 255504 298092
rect 255498 298052 255504 298064
rect 255556 298052 255562 298104
rect 265250 298092 265256 298104
rect 265211 298064 265256 298092
rect 265250 298052 265256 298064
rect 265308 298052 265314 298104
rect 267001 298095 267059 298101
rect 267001 298061 267013 298095
rect 267047 298092 267059 298095
rect 267090 298092 267096 298104
rect 267047 298064 267096 298092
rect 267047 298061 267059 298064
rect 267001 298055 267059 298061
rect 267090 298052 267096 298064
rect 267148 298052 267154 298104
rect 270770 298052 270776 298104
rect 270828 298092 270834 298104
rect 270862 298092 270868 298104
rect 270828 298064 270868 298092
rect 270828 298052 270834 298064
rect 270862 298052 270868 298064
rect 270920 298052 270926 298104
rect 277578 298092 277584 298104
rect 277539 298064 277584 298092
rect 277578 298052 277584 298064
rect 277636 298052 277642 298104
rect 292669 298095 292727 298101
rect 292669 298061 292681 298095
rect 292715 298092 292727 298095
rect 292758 298092 292764 298104
rect 292715 298064 292764 298092
rect 292715 298061 292727 298064
rect 292669 298055 292727 298061
rect 292758 298052 292764 298064
rect 292816 298052 292822 298104
rect 295702 298092 295708 298104
rect 295663 298064 295708 298092
rect 295702 298052 295708 298064
rect 295760 298052 295766 298104
rect 331398 298092 331404 298104
rect 331359 298064 331404 298092
rect 331398 298052 331404 298064
rect 331456 298052 331462 298104
rect 334250 298092 334256 298104
rect 334211 298064 334256 298092
rect 334250 298052 334256 298064
rect 334308 298052 334314 298104
rect 352098 298052 352104 298104
rect 352156 298092 352162 298104
rect 353478 298092 353484 298104
rect 352156 298064 352236 298092
rect 353439 298064 353484 298092
rect 352156 298052 352162 298064
rect 352208 298036 352236 298064
rect 353478 298052 353484 298064
rect 353536 298052 353542 298104
rect 365898 298052 365904 298104
rect 365956 298052 365962 298104
rect 370130 298092 370136 298104
rect 370091 298064 370136 298092
rect 370130 298052 370136 298064
rect 370188 298052 370194 298104
rect 400490 298052 400496 298104
rect 400548 298092 400554 298104
rect 400582 298092 400588 298104
rect 400548 298064 400588 298092
rect 400548 298052 400554 298064
rect 400582 298052 400588 298064
rect 400640 298052 400646 298104
rect 261018 297984 261024 298036
rect 261076 298024 261082 298036
rect 261110 298024 261116 298036
rect 261076 297996 261116 298024
rect 261076 297984 261082 297996
rect 261110 297984 261116 297996
rect 261168 297984 261174 298036
rect 352190 297984 352196 298036
rect 352248 297984 352254 298036
rect 365916 297968 365944 298052
rect 365898 297916 365904 297968
rect 365956 297916 365962 297968
rect 298370 296664 298376 296676
rect 298331 296636 298376 296664
rect 298370 296624 298376 296636
rect 298428 296624 298434 296676
rect 3326 294380 3332 294432
rect 3384 294420 3390 294432
rect 7558 294420 7564 294432
rect 3384 294392 7564 294420
rect 3384 294380 3390 294392
rect 7558 294380 7564 294392
rect 7616 294380 7622 294432
rect 295702 293264 295708 293276
rect 295663 293236 295708 293264
rect 295702 293224 295708 293236
rect 295760 293224 295766 293276
rect 408770 293060 408776 293072
rect 408731 293032 408776 293060
rect 408770 293020 408776 293032
rect 408828 293020 408834 293072
rect 327258 292612 327264 292664
rect 327316 292612 327322 292664
rect 330018 292612 330024 292664
rect 330076 292612 330082 292664
rect 332778 292612 332784 292664
rect 332836 292612 332842 292664
rect 387978 292612 387984 292664
rect 388036 292612 388042 292664
rect 451550 292652 451556 292664
rect 451476 292624 451556 292652
rect 230658 292544 230664 292596
rect 230716 292584 230722 292596
rect 230842 292584 230848 292596
rect 230716 292556 230848 292584
rect 230716 292544 230722 292556
rect 230842 292544 230848 292556
rect 230900 292544 230906 292596
rect 327276 292528 327304 292612
rect 330036 292528 330064 292612
rect 332796 292528 332824 292612
rect 387996 292528 388024 292612
rect 451476 292528 451504 292624
rect 451550 292612 451556 292624
rect 451608 292612 451614 292664
rect 288618 292476 288624 292528
rect 288676 292476 288682 292528
rect 327258 292476 327264 292528
rect 327316 292476 327322 292528
rect 330018 292476 330024 292528
rect 330076 292476 330082 292528
rect 332778 292476 332784 292528
rect 332836 292476 332842 292528
rect 387978 292476 387984 292528
rect 388036 292476 388042 292528
rect 451458 292476 451464 292528
rect 451516 292476 451522 292528
rect 466454 292476 466460 292528
rect 466512 292516 466518 292528
rect 466638 292516 466644 292528
rect 466512 292488 466644 292516
rect 466512 292476 466518 292488
rect 466638 292476 466644 292488
rect 466696 292476 466702 292528
rect 471974 292476 471980 292528
rect 472032 292516 472038 292528
rect 472158 292516 472164 292528
rect 472032 292488 472164 292516
rect 472032 292476 472038 292488
rect 472158 292476 472164 292488
rect 472216 292476 472222 292528
rect 288636 292392 288664 292476
rect 288618 292340 288624 292392
rect 288676 292340 288682 292392
rect 357618 291864 357624 291916
rect 357676 291904 357682 291916
rect 357802 291904 357808 291916
rect 357676 291876 357808 291904
rect 357676 291864 357682 291876
rect 357802 291864 357808 291876
rect 357860 291864 357866 291916
rect 376846 289892 376852 289944
rect 376904 289932 376910 289944
rect 376904 289904 376984 289932
rect 376904 289892 376910 289904
rect 376956 289876 376984 289904
rect 241790 289864 241796 289876
rect 241751 289836 241796 289864
rect 241790 289824 241796 289836
rect 241848 289824 241854 289876
rect 281626 289864 281632 289876
rect 281587 289836 281632 289864
rect 281626 289824 281632 289836
rect 281684 289824 281690 289876
rect 305178 289864 305184 289876
rect 305139 289836 305184 289864
rect 305178 289824 305184 289836
rect 305236 289824 305242 289876
rect 309318 289824 309324 289876
rect 309376 289864 309382 289876
rect 309594 289864 309600 289876
rect 309376 289836 309600 289864
rect 309376 289824 309382 289836
rect 309594 289824 309600 289836
rect 309652 289824 309658 289876
rect 310698 289864 310704 289876
rect 310659 289836 310704 289864
rect 310698 289824 310704 289836
rect 310756 289824 310762 289876
rect 324498 289864 324504 289876
rect 324459 289836 324504 289864
rect 324498 289824 324504 289836
rect 324556 289824 324562 289876
rect 346578 289864 346584 289876
rect 346539 289836 346584 289864
rect 346578 289824 346584 289836
rect 346636 289824 346642 289876
rect 376938 289824 376944 289876
rect 376996 289824 377002 289876
rect 381078 289824 381084 289876
rect 381136 289864 381142 289876
rect 381354 289864 381360 289876
rect 381136 289836 381360 289864
rect 381136 289824 381142 289836
rect 381354 289824 381360 289836
rect 381412 289824 381418 289876
rect 382458 289864 382464 289876
rect 382419 289836 382464 289864
rect 382458 289824 382464 289836
rect 382516 289824 382522 289876
rect 259638 289796 259644 289808
rect 259599 289768 259644 289796
rect 259638 289756 259644 289768
rect 259696 289756 259702 289808
rect 287238 289796 287244 289808
rect 287199 289768 287244 289796
rect 287238 289756 287244 289768
rect 287296 289756 287302 289808
rect 347958 289756 347964 289808
rect 348016 289756 348022 289808
rect 356422 289756 356428 289808
rect 356480 289756 356486 289808
rect 375558 289756 375564 289808
rect 375616 289796 375622 289808
rect 375742 289796 375748 289808
rect 375616 289768 375748 289796
rect 375616 289756 375622 289768
rect 375742 289756 375748 289768
rect 375800 289756 375806 289808
rect 392118 289756 392124 289808
rect 392176 289796 392182 289808
rect 392210 289796 392216 289808
rect 392176 289768 392216 289796
rect 392176 289756 392182 289768
rect 392210 289756 392216 289768
rect 392268 289756 392274 289808
rect 236273 289731 236331 289737
rect 236273 289697 236285 289731
rect 236319 289728 236331 289731
rect 236454 289728 236460 289740
rect 236319 289700 236460 289728
rect 236319 289697 236331 289700
rect 236273 289691 236331 289697
rect 236454 289688 236460 289700
rect 236512 289688 236518 289740
rect 309318 289728 309324 289740
rect 309279 289700 309324 289728
rect 309318 289688 309324 289700
rect 309376 289688 309382 289740
rect 347976 289728 348004 289756
rect 348050 289728 348056 289740
rect 347976 289700 348056 289728
rect 348050 289688 348056 289700
rect 348108 289688 348114 289740
rect 356440 289728 356468 289756
rect 356514 289728 356520 289740
rect 356440 289700 356520 289728
rect 356514 289688 356520 289700
rect 356572 289688 356578 289740
rect 370133 289731 370191 289737
rect 370133 289697 370145 289731
rect 370179 289728 370191 289731
rect 370222 289728 370228 289740
rect 370179 289700 370228 289728
rect 370179 289697 370191 289700
rect 370133 289691 370191 289697
rect 370222 289688 370228 289700
rect 370280 289688 370286 289740
rect 249886 288436 249892 288448
rect 249847 288408 249892 288436
rect 249886 288396 249892 288408
rect 249944 288396 249950 288448
rect 255498 288436 255504 288448
rect 255459 288408 255504 288436
rect 255498 288396 255504 288408
rect 255556 288396 255562 288448
rect 265250 288436 265256 288448
rect 265211 288408 265256 288436
rect 265250 288396 265256 288408
rect 265308 288396 265314 288448
rect 292666 288436 292672 288448
rect 292627 288408 292672 288436
rect 292666 288396 292672 288408
rect 292724 288396 292730 288448
rect 331398 288436 331404 288448
rect 331359 288408 331404 288436
rect 331398 288396 331404 288408
rect 331456 288396 331462 288448
rect 353481 288439 353539 288445
rect 353481 288405 353493 288439
rect 353527 288436 353539 288439
rect 353570 288436 353576 288448
rect 353527 288408 353576 288436
rect 353527 288405 353539 288408
rect 353481 288399 353539 288405
rect 353570 288396 353576 288408
rect 353628 288396 353634 288448
rect 298373 287079 298431 287085
rect 298373 287045 298385 287079
rect 298419 287076 298431 287079
rect 298462 287076 298468 287088
rect 298419 287048 298468 287076
rect 298419 287045 298431 287048
rect 298373 287039 298431 287045
rect 298462 287036 298468 287048
rect 298520 287036 298526 287088
rect 352006 287036 352012 287088
rect 352064 287076 352070 287088
rect 352098 287076 352104 287088
rect 352064 287048 352104 287076
rect 352064 287036 352070 287048
rect 352098 287036 352104 287048
rect 352156 287036 352162 287088
rect 231946 285880 231952 285932
rect 232004 285920 232010 285932
rect 232314 285920 232320 285932
rect 232004 285892 232320 285920
rect 232004 285880 232010 285892
rect 232314 285880 232320 285892
rect 232372 285880 232378 285932
rect 249886 285852 249892 285864
rect 249847 285824 249892 285852
rect 249886 285812 249892 285824
rect 249944 285812 249950 285864
rect 230658 282956 230664 283008
rect 230716 282956 230722 283008
rect 230676 282872 230704 282956
rect 331398 282888 331404 282940
rect 331456 282888 331462 282940
rect 342530 282928 342536 282940
rect 342491 282900 342536 282928
rect 342530 282888 342536 282900
rect 342588 282888 342594 282940
rect 364518 282888 364524 282940
rect 364576 282888 364582 282940
rect 381078 282888 381084 282940
rect 381136 282888 381142 282940
rect 422294 282888 422300 282940
rect 422352 282928 422358 282940
rect 422478 282928 422484 282940
rect 422352 282900 422484 282928
rect 422352 282888 422358 282900
rect 422478 282888 422484 282900
rect 422536 282888 422542 282940
rect 427814 282888 427820 282940
rect 427872 282928 427878 282940
rect 427998 282928 428004 282940
rect 427872 282900 428004 282928
rect 427872 282888 427878 282900
rect 427998 282888 428004 282900
rect 428056 282888 428062 282940
rect 230658 282820 230664 282872
rect 230716 282820 230722 282872
rect 242986 282820 242992 282872
rect 243044 282860 243050 282872
rect 243170 282860 243176 282872
rect 243044 282832 243176 282860
rect 243044 282820 243050 282832
rect 243170 282820 243176 282832
rect 243228 282820 243234 282872
rect 259641 282795 259699 282801
rect 259641 282761 259653 282795
rect 259687 282792 259699 282795
rect 259730 282792 259736 282804
rect 259687 282764 259736 282792
rect 259687 282761 259699 282764
rect 259641 282755 259699 282761
rect 259730 282752 259736 282764
rect 259788 282752 259794 282804
rect 331416 282792 331444 282888
rect 331490 282792 331496 282804
rect 331416 282764 331496 282792
rect 331490 282752 331496 282764
rect 331548 282752 331554 282804
rect 334253 282795 334311 282801
rect 334253 282761 334265 282795
rect 334299 282792 334311 282795
rect 334434 282792 334440 282804
rect 334299 282764 334440 282792
rect 334299 282761 334311 282764
rect 334253 282755 334311 282761
rect 334434 282752 334440 282764
rect 334492 282752 334498 282804
rect 364536 282792 364564 282888
rect 364610 282792 364616 282804
rect 364536 282764 364616 282792
rect 364610 282752 364616 282764
rect 364668 282752 364674 282804
rect 381096 282792 381124 282888
rect 381170 282792 381176 282804
rect 381096 282764 381176 282792
rect 381170 282752 381176 282764
rect 381228 282752 381234 282804
rect 408770 282792 408776 282804
rect 408731 282764 408776 282792
rect 408770 282752 408776 282764
rect 408828 282752 408834 282804
rect 342530 280276 342536 280288
rect 342491 280248 342536 280276
rect 342530 280236 342536 280248
rect 342588 280236 342594 280288
rect 266998 280208 267004 280220
rect 266959 280180 267004 280208
rect 266998 280168 267004 280180
rect 267056 280168 267062 280220
rect 277581 280211 277639 280217
rect 277581 280177 277593 280211
rect 277627 280208 277639 280211
rect 277670 280208 277676 280220
rect 277627 280180 277676 280208
rect 277627 280177 277639 280180
rect 277581 280171 277639 280177
rect 277670 280168 277676 280180
rect 277728 280168 277734 280220
rect 281718 280168 281724 280220
rect 281776 280208 281782 280220
rect 281902 280208 281908 280220
rect 281776 280180 281908 280208
rect 281776 280168 281782 280180
rect 281902 280168 281908 280180
rect 281960 280168 281966 280220
rect 287238 280208 287244 280220
rect 287199 280180 287244 280208
rect 287238 280168 287244 280180
rect 287296 280168 287302 280220
rect 292666 280168 292672 280220
rect 292724 280208 292730 280220
rect 292758 280208 292764 280220
rect 292724 280180 292764 280208
rect 292724 280168 292730 280180
rect 292758 280168 292764 280180
rect 292816 280168 292822 280220
rect 309321 280211 309379 280217
rect 309321 280177 309333 280211
rect 309367 280208 309379 280211
rect 309410 280208 309416 280220
rect 309367 280180 309416 280208
rect 309367 280177 309379 280180
rect 309321 280171 309379 280177
rect 309410 280168 309416 280180
rect 309468 280168 309474 280220
rect 324406 280168 324412 280220
rect 324464 280208 324470 280220
rect 324682 280208 324688 280220
rect 324464 280180 324688 280208
rect 324464 280168 324470 280180
rect 324682 280168 324688 280180
rect 324740 280168 324746 280220
rect 352006 280168 352012 280220
rect 352064 280208 352070 280220
rect 352064 280180 352144 280208
rect 352064 280168 352070 280180
rect 352116 280152 352144 280180
rect 3142 280100 3148 280152
rect 3200 280140 3206 280152
rect 6270 280140 6276 280152
rect 3200 280112 6276 280140
rect 3200 280100 3206 280112
rect 6270 280100 6276 280112
rect 6328 280100 6334 280152
rect 230658 280100 230664 280152
rect 230716 280140 230722 280152
rect 230845 280143 230903 280149
rect 230845 280140 230857 280143
rect 230716 280112 230857 280140
rect 230716 280100 230722 280112
rect 230845 280109 230857 280112
rect 230891 280109 230903 280143
rect 230845 280103 230903 280109
rect 233326 280100 233332 280152
rect 233384 280140 233390 280152
rect 233510 280140 233516 280152
rect 233384 280112 233516 280140
rect 233384 280100 233390 280112
rect 233510 280100 233516 280112
rect 233568 280100 233574 280152
rect 241790 280140 241796 280152
rect 241751 280112 241796 280140
rect 241790 280100 241796 280112
rect 241848 280100 241854 280152
rect 242802 280100 242808 280152
rect 242860 280140 242866 280152
rect 243170 280140 243176 280152
rect 242860 280112 243176 280140
rect 242860 280100 242866 280112
rect 243170 280100 243176 280112
rect 243228 280100 243234 280152
rect 244458 280100 244464 280152
rect 244516 280140 244522 280152
rect 244550 280140 244556 280152
rect 244516 280112 244556 280140
rect 244516 280100 244522 280112
rect 244550 280100 244556 280112
rect 244608 280100 244614 280152
rect 265158 280100 265164 280152
rect 265216 280140 265222 280152
rect 265250 280140 265256 280152
rect 265216 280112 265256 280140
rect 265216 280100 265222 280112
rect 265250 280100 265256 280112
rect 265308 280100 265314 280152
rect 270586 280100 270592 280152
rect 270644 280140 270650 280152
rect 270862 280140 270868 280152
rect 270644 280112 270868 280140
rect 270644 280100 270650 280112
rect 270862 280100 270868 280112
rect 270920 280100 270926 280152
rect 283098 280140 283104 280152
rect 283059 280112 283104 280140
rect 283098 280100 283104 280112
rect 283156 280100 283162 280152
rect 295426 280100 295432 280152
rect 295484 280140 295490 280152
rect 295702 280140 295708 280152
rect 295484 280112 295708 280140
rect 295484 280100 295490 280112
rect 295702 280100 295708 280112
rect 295760 280100 295766 280152
rect 298462 280140 298468 280152
rect 298296 280112 298468 280140
rect 298296 280084 298324 280112
rect 298462 280100 298468 280112
rect 298520 280100 298526 280152
rect 305178 280140 305184 280152
rect 305139 280112 305184 280140
rect 305178 280100 305184 280112
rect 305236 280100 305242 280152
rect 310698 280140 310704 280152
rect 310659 280112 310704 280140
rect 310698 280100 310704 280112
rect 310756 280100 310762 280152
rect 318978 280100 318984 280152
rect 319036 280140 319042 280152
rect 319070 280140 319076 280152
rect 319036 280112 319076 280140
rect 319036 280100 319042 280112
rect 319070 280100 319076 280112
rect 319128 280100 319134 280152
rect 327258 280140 327264 280152
rect 327219 280112 327264 280140
rect 327258 280100 327264 280112
rect 327316 280100 327322 280152
rect 331122 280100 331128 280152
rect 331180 280140 331186 280152
rect 331490 280140 331496 280152
rect 331180 280112 331496 280140
rect 331180 280100 331186 280112
rect 331490 280100 331496 280112
rect 331548 280100 331554 280152
rect 334345 280143 334403 280149
rect 334345 280109 334357 280143
rect 334391 280140 334403 280143
rect 334434 280140 334440 280152
rect 334391 280112 334440 280140
rect 334391 280109 334403 280112
rect 334345 280103 334403 280109
rect 334434 280100 334440 280112
rect 334492 280100 334498 280152
rect 346578 280140 346584 280152
rect 346539 280112 346584 280140
rect 346578 280100 346584 280112
rect 346636 280100 346642 280152
rect 352098 280100 352104 280152
rect 352156 280100 352162 280152
rect 353570 280100 353576 280152
rect 353628 280140 353634 280152
rect 353662 280140 353668 280152
rect 353628 280112 353668 280140
rect 353628 280100 353634 280112
rect 353662 280100 353668 280112
rect 353720 280100 353726 280152
rect 356422 280100 356428 280152
rect 356480 280140 356486 280152
rect 356514 280140 356520 280152
rect 356480 280112 356520 280140
rect 356480 280100 356486 280112
rect 356514 280100 356520 280112
rect 356572 280100 356578 280152
rect 358998 280100 359004 280152
rect 359056 280140 359062 280152
rect 359090 280140 359096 280152
rect 359056 280112 359096 280140
rect 359056 280100 359062 280112
rect 359090 280100 359096 280112
rect 359148 280100 359154 280152
rect 364521 280143 364579 280149
rect 364521 280109 364533 280143
rect 364567 280140 364579 280143
rect 364610 280140 364616 280152
rect 364567 280112 364616 280140
rect 364567 280109 364579 280112
rect 364521 280103 364579 280109
rect 364610 280100 364616 280112
rect 364668 280100 364674 280152
rect 369946 280100 369952 280152
rect 370004 280140 370010 280152
rect 370222 280140 370228 280152
rect 370004 280112 370228 280140
rect 370004 280100 370010 280112
rect 370222 280100 370228 280112
rect 370280 280100 370286 280152
rect 371418 280140 371424 280152
rect 371379 280112 371424 280140
rect 371418 280100 371424 280112
rect 371476 280100 371482 280152
rect 375466 280100 375472 280152
rect 375524 280140 375530 280152
rect 375742 280140 375748 280152
rect 375524 280112 375748 280140
rect 375524 280100 375530 280112
rect 375742 280100 375748 280112
rect 375800 280100 375806 280152
rect 376938 280140 376944 280152
rect 376899 280112 376944 280140
rect 376938 280100 376944 280112
rect 376996 280100 377002 280152
rect 386690 280100 386696 280152
rect 386748 280140 386754 280152
rect 386782 280140 386788 280152
rect 386748 280112 386788 280140
rect 386748 280100 386754 280112
rect 386782 280100 386788 280112
rect 386840 280100 386846 280152
rect 387978 280100 387984 280152
rect 388036 280140 388042 280152
rect 388070 280140 388076 280152
rect 388036 280112 388076 280140
rect 388036 280100 388042 280112
rect 388070 280100 388076 280112
rect 388128 280100 388134 280152
rect 393222 280140 393228 280152
rect 393183 280112 393228 280140
rect 393222 280100 393228 280112
rect 393280 280100 393286 280152
rect 400490 280140 400496 280152
rect 400451 280112 400496 280140
rect 400490 280100 400496 280112
rect 400548 280100 400554 280152
rect 416866 280140 416872 280152
rect 416827 280112 416872 280140
rect 416866 280100 416872 280112
rect 416924 280100 416930 280152
rect 433610 280140 433616 280152
rect 433571 280112 433616 280140
rect 433610 280100 433616 280112
rect 433668 280100 433674 280152
rect 466546 280140 466552 280152
rect 466507 280112 466552 280140
rect 466546 280100 466552 280112
rect 466604 280100 466610 280152
rect 472066 280140 472072 280152
rect 472027 280112 472072 280140
rect 472066 280100 472072 280112
rect 472124 280100 472130 280152
rect 298278 280032 298284 280084
rect 298336 280032 298342 280084
rect 348050 278848 348056 278860
rect 347976 278820 348056 278848
rect 347976 278792 348004 278820
rect 348050 278808 348056 278820
rect 348108 278808 348114 278860
rect 236362 278740 236368 278792
rect 236420 278780 236426 278792
rect 236638 278780 236644 278792
rect 236420 278752 236644 278780
rect 236420 278740 236426 278752
rect 236638 278740 236644 278752
rect 236696 278740 236702 278792
rect 249889 278783 249947 278789
rect 249889 278749 249901 278783
rect 249935 278780 249947 278783
rect 250070 278780 250076 278792
rect 249935 278752 250076 278780
rect 249935 278749 249947 278752
rect 249889 278743 249947 278749
rect 250070 278740 250076 278752
rect 250128 278740 250134 278792
rect 254210 278740 254216 278792
rect 254268 278780 254274 278792
rect 254486 278780 254492 278792
rect 254268 278752 254492 278780
rect 254268 278740 254274 278752
rect 254486 278740 254492 278752
rect 254544 278740 254550 278792
rect 347958 278740 347964 278792
rect 348016 278740 348022 278792
rect 392118 278740 392124 278792
rect 392176 278780 392182 278792
rect 392210 278780 392216 278792
rect 392176 278752 392216 278780
rect 392176 278740 392182 278752
rect 392210 278740 392216 278752
rect 392268 278740 392274 278792
rect 451274 278740 451280 278792
rect 451332 278780 451338 278792
rect 451550 278780 451556 278792
rect 451332 278752 451556 278780
rect 451332 278740 451338 278752
rect 451550 278740 451556 278752
rect 451608 278740 451614 278792
rect 270586 278712 270592 278724
rect 270547 278684 270592 278712
rect 270586 278672 270592 278684
rect 270644 278672 270650 278724
rect 295426 278712 295432 278724
rect 295387 278684 295432 278712
rect 295426 278672 295432 278684
rect 295484 278672 295490 278724
rect 375466 278712 375472 278724
rect 375427 278684 375472 278712
rect 375466 278672 375472 278684
rect 375524 278672 375530 278724
rect 408770 278712 408776 278724
rect 408731 278684 408776 278712
rect 408770 278672 408776 278684
rect 408828 278672 408834 278724
rect 277670 275108 277676 275120
rect 277631 275080 277676 275108
rect 277670 275068 277676 275080
rect 277728 275068 277734 275120
rect 451550 273748 451556 273760
rect 451511 273720 451556 273748
rect 451550 273708 451556 273720
rect 451608 273708 451614 273760
rect 254210 273340 254216 273352
rect 254136 273312 254216 273340
rect 230842 273272 230848 273284
rect 230803 273244 230848 273272
rect 230842 273232 230848 273244
rect 230900 273232 230906 273284
rect 254136 273216 254164 273312
rect 254210 273300 254216 273312
rect 254268 273300 254274 273352
rect 330018 273300 330024 273352
rect 330076 273300 330082 273352
rect 332778 273300 332784 273352
rect 332836 273300 332842 273352
rect 356422 273300 356428 273352
rect 356480 273300 356486 273352
rect 357618 273300 357624 273352
rect 357676 273300 357682 273352
rect 330036 273216 330064 273300
rect 332796 273216 332824 273300
rect 356440 273216 356468 273300
rect 357636 273216 357664 273300
rect 254118 273164 254124 273216
rect 254176 273164 254182 273216
rect 272058 273164 272064 273216
rect 272116 273164 272122 273216
rect 288618 273164 288624 273216
rect 288676 273164 288682 273216
rect 294138 273164 294144 273216
rect 294196 273164 294202 273216
rect 330018 273164 330024 273216
rect 330076 273164 330082 273216
rect 332778 273164 332784 273216
rect 332836 273164 332842 273216
rect 356422 273164 356428 273216
rect 356480 273164 356486 273216
rect 357618 273164 357624 273216
rect 357676 273164 357682 273216
rect 364518 273204 364524 273216
rect 364479 273176 364524 273204
rect 364518 273164 364524 273176
rect 364576 273164 364582 273216
rect 382458 273164 382464 273216
rect 382516 273164 382522 273216
rect 272076 273080 272104 273164
rect 288636 273080 288664 273164
rect 294156 273080 294184 273164
rect 382476 273080 382504 273164
rect 272058 273028 272064 273080
rect 272116 273028 272122 273080
rect 288618 273028 288624 273080
rect 288676 273028 288682 273080
rect 294138 273028 294144 273080
rect 294196 273028 294202 273080
rect 382458 273028 382464 273080
rect 382516 273028 382522 273080
rect 327258 272184 327264 272196
rect 327219 272156 327264 272184
rect 327258 272144 327264 272156
rect 327316 272144 327322 272196
rect 334342 270620 334348 270632
rect 334303 270592 334348 270620
rect 334342 270580 334348 270592
rect 334400 270580 334406 270632
rect 232038 270512 232044 270564
rect 232096 270552 232102 270564
rect 232314 270552 232320 270564
rect 232096 270524 232320 270552
rect 232096 270512 232102 270524
rect 232314 270512 232320 270524
rect 232372 270512 232378 270564
rect 236362 270552 236368 270564
rect 236288 270524 236368 270552
rect 236288 270496 236316 270524
rect 236362 270512 236368 270524
rect 236420 270512 236426 270564
rect 241790 270552 241796 270564
rect 241751 270524 241796 270552
rect 241790 270512 241796 270524
rect 241848 270512 241854 270564
rect 266998 270512 267004 270564
rect 267056 270552 267062 270564
rect 267090 270552 267096 270564
rect 267056 270524 267096 270552
rect 267056 270512 267062 270524
rect 267090 270512 267096 270524
rect 267148 270512 267154 270564
rect 283098 270552 283104 270564
rect 283059 270524 283104 270552
rect 283098 270512 283104 270524
rect 283156 270512 283162 270564
rect 305178 270552 305184 270564
rect 305139 270524 305184 270552
rect 305178 270512 305184 270524
rect 305236 270512 305242 270564
rect 309318 270512 309324 270564
rect 309376 270552 309382 270564
rect 309594 270552 309600 270564
rect 309376 270524 309600 270552
rect 309376 270512 309382 270524
rect 309594 270512 309600 270524
rect 309652 270512 309658 270564
rect 310698 270552 310704 270564
rect 310659 270524 310704 270552
rect 310698 270512 310704 270524
rect 310756 270512 310762 270564
rect 346578 270552 346584 270564
rect 346539 270524 346584 270552
rect 346578 270512 346584 270524
rect 346636 270512 346642 270564
rect 371418 270552 371424 270564
rect 371379 270524 371424 270552
rect 371418 270512 371424 270524
rect 371476 270512 371482 270564
rect 376938 270552 376944 270564
rect 376899 270524 376944 270552
rect 376938 270512 376944 270524
rect 376996 270512 377002 270564
rect 380986 270512 380992 270564
rect 381044 270552 381050 270564
rect 381078 270552 381084 270564
rect 381044 270524 381084 270552
rect 381044 270512 381050 270524
rect 381078 270512 381084 270524
rect 381136 270512 381142 270564
rect 393222 270552 393228 270564
rect 393183 270524 393228 270552
rect 393222 270512 393228 270524
rect 393280 270512 393286 270564
rect 400493 270555 400551 270561
rect 400493 270521 400505 270555
rect 400539 270552 400551 270555
rect 400582 270552 400588 270564
rect 400539 270524 400588 270552
rect 400539 270521 400551 270524
rect 400493 270515 400551 270521
rect 400582 270512 400588 270524
rect 400640 270512 400646 270564
rect 416869 270555 416927 270561
rect 416869 270521 416881 270555
rect 416915 270552 416927 270555
rect 416958 270552 416964 270564
rect 416915 270524 416964 270552
rect 416915 270521 416927 270524
rect 416869 270515 416927 270521
rect 416958 270512 416964 270524
rect 417016 270512 417022 270564
rect 433613 270555 433671 270561
rect 433613 270521 433625 270555
rect 433659 270552 433671 270555
rect 433702 270552 433708 270564
rect 433659 270524 433708 270552
rect 433659 270521 433671 270524
rect 433613 270515 433671 270521
rect 433702 270512 433708 270524
rect 433760 270512 433766 270564
rect 466549 270555 466607 270561
rect 466549 270521 466561 270555
rect 466595 270552 466607 270555
rect 466638 270552 466644 270564
rect 466595 270524 466644 270552
rect 466595 270521 466607 270524
rect 466549 270515 466607 270521
rect 466638 270512 466644 270524
rect 466696 270512 466702 270564
rect 472069 270555 472127 270561
rect 472069 270521 472081 270555
rect 472115 270552 472127 270555
rect 472158 270552 472164 270564
rect 472115 270524 472164 270552
rect 472115 270521 472127 270524
rect 472069 270515 472127 270521
rect 472158 270512 472164 270524
rect 472216 270512 472222 270564
rect 236270 270444 236276 270496
rect 236328 270444 236334 270496
rect 252738 270484 252744 270496
rect 252699 270456 252744 270484
rect 252738 270444 252744 270456
rect 252796 270444 252802 270496
rect 287238 270484 287244 270496
rect 287199 270456 287244 270484
rect 287238 270444 287244 270456
rect 287296 270444 287302 270496
rect 392118 270484 392124 270496
rect 392079 270456 392124 270484
rect 392118 270444 392124 270456
rect 392176 270444 392182 270496
rect 309318 270416 309324 270428
rect 309279 270388 309324 270416
rect 309318 270376 309324 270388
rect 309376 270376 309382 270428
rect 381078 270416 381084 270428
rect 381039 270388 381084 270416
rect 381078 270376 381084 270388
rect 381136 270376 381142 270428
rect 270589 269127 270647 269133
rect 270589 269093 270601 269127
rect 270635 269124 270647 269127
rect 270770 269124 270776 269136
rect 270635 269096 270776 269124
rect 270635 269093 270647 269096
rect 270589 269087 270647 269093
rect 270770 269084 270776 269096
rect 270828 269084 270834 269136
rect 277673 269127 277731 269133
rect 277673 269093 277685 269127
rect 277719 269124 277731 269127
rect 277762 269124 277768 269136
rect 277719 269096 277768 269124
rect 277719 269093 277731 269096
rect 277673 269087 277731 269093
rect 277762 269084 277768 269096
rect 277820 269084 277826 269136
rect 295429 269127 295487 269133
rect 295429 269093 295441 269127
rect 295475 269124 295487 269127
rect 295610 269124 295616 269136
rect 295475 269096 295616 269124
rect 295475 269093 295487 269096
rect 295429 269087 295487 269093
rect 295610 269084 295616 269096
rect 295668 269084 295674 269136
rect 259362 267724 259368 267776
rect 259420 267764 259426 267776
rect 259546 267764 259552 267776
rect 259420 267736 259552 267764
rect 259420 267724 259426 267736
rect 259546 267724 259552 267736
rect 259604 267724 259610 267776
rect 3326 266296 3332 266348
rect 3384 266336 3390 266348
rect 229738 266336 229744 266348
rect 3384 266308 229744 266336
rect 3384 266296 3390 266308
rect 229738 266296 229744 266308
rect 229796 266296 229802 266348
rect 530762 264868 530768 264920
rect 530820 264908 530826 264920
rect 580166 264908 580172 264920
rect 530820 264880 580172 264908
rect 530820 264868 530826 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 392121 264299 392179 264305
rect 392121 264265 392133 264299
rect 392167 264296 392179 264299
rect 392210 264296 392216 264308
rect 392167 264268 392216 264296
rect 392167 264265 392179 264268
rect 392121 264259 392179 264265
rect 392210 264256 392216 264268
rect 392268 264256 392274 264308
rect 230842 263576 230848 263628
rect 230900 263576 230906 263628
rect 231857 263619 231915 263625
rect 231857 263585 231869 263619
rect 231903 263616 231915 263619
rect 231946 263616 231952 263628
rect 231903 263588 231952 263616
rect 231903 263585 231915 263588
rect 231857 263579 231915 263585
rect 231946 263576 231952 263588
rect 232004 263576 232010 263628
rect 236270 263576 236276 263628
rect 236328 263616 236334 263628
rect 236328 263588 236408 263616
rect 236328 263576 236334 263588
rect 230860 263480 230888 263576
rect 236380 263560 236408 263588
rect 243170 263576 243176 263628
rect 243228 263576 243234 263628
rect 266998 263616 267004 263628
rect 266959 263588 267004 263616
rect 266998 263576 267004 263588
rect 267056 263576 267062 263628
rect 324406 263616 324412 263628
rect 324367 263588 324412 263616
rect 324406 263576 324412 263588
rect 324464 263576 324470 263628
rect 334342 263576 334348 263628
rect 334400 263576 334406 263628
rect 342530 263616 342536 263628
rect 342491 263588 342536 263616
rect 342530 263576 342536 263588
rect 342588 263576 342594 263628
rect 364518 263576 364524 263628
rect 364576 263576 364582 263628
rect 422294 263576 422300 263628
rect 422352 263616 422358 263628
rect 422478 263616 422484 263628
rect 422352 263588 422484 263616
rect 422352 263576 422358 263588
rect 422478 263576 422484 263588
rect 422536 263576 422542 263628
rect 427814 263576 427820 263628
rect 427872 263616 427878 263628
rect 427998 263616 428004 263628
rect 427872 263588 428004 263616
rect 427872 263576 427878 263588
rect 427998 263576 428004 263588
rect 428056 263576 428062 263628
rect 236362 263508 236368 263560
rect 236420 263508 236426 263560
rect 243188 263492 243216 263576
rect 331306 263508 331312 263560
rect 331364 263548 331370 263560
rect 331364 263520 331536 263548
rect 331364 263508 331370 263520
rect 331508 263492 331536 263520
rect 230934 263480 230940 263492
rect 230860 263452 230940 263480
rect 230934 263440 230940 263452
rect 230992 263440 230998 263492
rect 243170 263440 243176 263492
rect 243228 263440 243234 263492
rect 331490 263440 331496 263492
rect 331548 263440 331554 263492
rect 334360 263480 334388 263576
rect 358906 263508 358912 263560
rect 358964 263548 358970 263560
rect 358964 263520 359136 263548
rect 358964 263508 358970 263520
rect 359108 263492 359136 263520
rect 334434 263480 334440 263492
rect 334360 263452 334440 263480
rect 334434 263440 334440 263452
rect 334492 263440 334498 263492
rect 352006 263440 352012 263492
rect 352064 263480 352070 263492
rect 352282 263480 352288 263492
rect 352064 263452 352288 263480
rect 352064 263440 352070 263452
rect 352282 263440 352288 263452
rect 352340 263440 352346 263492
rect 359090 263440 359096 263492
rect 359148 263440 359154 263492
rect 364536 263480 364564 263576
rect 364610 263480 364616 263492
rect 364536 263452 364616 263480
rect 364610 263440 364616 263452
rect 364668 263440 364674 263492
rect 375469 263483 375527 263489
rect 375469 263449 375481 263483
rect 375515 263480 375527 263483
rect 375650 263480 375656 263492
rect 375515 263452 375656 263480
rect 375515 263449 375527 263452
rect 375469 263443 375527 263449
rect 375650 263440 375656 263452
rect 375708 263440 375714 263492
rect 397362 263440 397368 263492
rect 397420 263480 397426 263492
rect 397730 263480 397736 263492
rect 397420 263452 397736 263480
rect 397420 263440 397426 263452
rect 397730 263440 397736 263452
rect 397788 263440 397794 263492
rect 408770 263480 408776 263492
rect 408731 263452 408776 263480
rect 408770 263440 408776 263452
rect 408828 263440 408834 263492
rect 451550 263480 451556 263492
rect 451511 263452 451556 263480
rect 451550 263440 451556 263452
rect 451608 263440 451614 263492
rect 252738 260896 252744 260908
rect 252699 260868 252744 260896
rect 252738 260856 252744 260868
rect 252796 260856 252802 260908
rect 287238 260896 287244 260908
rect 287199 260868 287244 260896
rect 287238 260856 287244 260868
rect 287296 260856 287302 260908
rect 292758 260856 292764 260908
rect 292816 260856 292822 260908
rect 309321 260899 309379 260905
rect 309321 260865 309333 260899
rect 309367 260896 309379 260899
rect 309410 260896 309416 260908
rect 309367 260868 309416 260896
rect 309367 260865 309379 260868
rect 309321 260859 309379 260865
rect 309410 260856 309416 260868
rect 309468 260856 309474 260908
rect 324406 260896 324412 260908
rect 324367 260868 324412 260896
rect 324406 260856 324412 260868
rect 324464 260856 324470 260908
rect 342530 260896 342536 260908
rect 342491 260868 342536 260896
rect 342530 260856 342536 260868
rect 342588 260856 342594 260908
rect 348050 260856 348056 260908
rect 348108 260856 348114 260908
rect 356514 260896 356520 260908
rect 356440 260868 356520 260896
rect 241790 260828 241796 260840
rect 241751 260800 241796 260828
rect 241790 260788 241796 260800
rect 241848 260788 241854 260840
rect 242802 260788 242808 260840
rect 242860 260828 242866 260840
rect 243170 260828 243176 260840
rect 242860 260800 243176 260828
rect 242860 260788 242866 260800
rect 243170 260788 243176 260800
rect 243228 260788 243234 260840
rect 244458 260788 244464 260840
rect 244516 260788 244522 260840
rect 249978 260788 249984 260840
rect 250036 260788 250042 260840
rect 254026 260788 254032 260840
rect 254084 260828 254090 260840
rect 254210 260828 254216 260840
rect 254084 260800 254216 260828
rect 254084 260788 254090 260800
rect 254210 260788 254216 260800
rect 254268 260788 254274 260840
rect 255498 260788 255504 260840
rect 255556 260788 255562 260840
rect 277578 260788 277584 260840
rect 277636 260828 277642 260840
rect 277670 260828 277676 260840
rect 277636 260800 277676 260828
rect 277636 260788 277642 260800
rect 277670 260788 277676 260800
rect 277728 260788 277734 260840
rect 283098 260828 283104 260840
rect 283059 260800 283104 260828
rect 283098 260788 283104 260800
rect 283156 260788 283162 260840
rect 244476 260760 244504 260788
rect 244550 260760 244556 260772
rect 244476 260732 244556 260760
rect 244550 260720 244556 260732
rect 244608 260720 244614 260772
rect 249996 260760 250024 260788
rect 250070 260760 250076 260772
rect 249996 260732 250076 260760
rect 250070 260720 250076 260732
rect 250128 260720 250134 260772
rect 255516 260760 255544 260788
rect 292776 260772 292804 260856
rect 295426 260788 295432 260840
rect 295484 260828 295490 260840
rect 295610 260828 295616 260840
rect 295484 260800 295616 260828
rect 295484 260788 295490 260800
rect 295610 260788 295616 260800
rect 295668 260788 295674 260840
rect 305178 260828 305184 260840
rect 305139 260800 305184 260828
rect 305178 260788 305184 260800
rect 305236 260788 305242 260840
rect 310698 260828 310704 260840
rect 310659 260800 310704 260828
rect 310698 260788 310704 260800
rect 310756 260788 310762 260840
rect 318978 260788 318984 260840
rect 319036 260828 319042 260840
rect 319070 260828 319076 260840
rect 319036 260800 319076 260828
rect 319036 260788 319042 260800
rect 319070 260788 319076 260800
rect 319128 260788 319134 260840
rect 327258 260828 327264 260840
rect 327219 260800 327264 260828
rect 327258 260788 327264 260800
rect 327316 260788 327322 260840
rect 331122 260788 331128 260840
rect 331180 260828 331186 260840
rect 331490 260828 331496 260840
rect 331180 260800 331496 260828
rect 331180 260788 331186 260800
rect 331490 260788 331496 260800
rect 331548 260788 331554 260840
rect 334345 260831 334403 260837
rect 334345 260797 334357 260831
rect 334391 260828 334403 260831
rect 334434 260828 334440 260840
rect 334391 260800 334440 260828
rect 334391 260797 334403 260800
rect 334345 260791 334403 260797
rect 334434 260788 334440 260800
rect 334492 260788 334498 260840
rect 346578 260828 346584 260840
rect 346539 260800 346584 260828
rect 346578 260788 346584 260800
rect 346636 260788 346642 260840
rect 348068 260828 348096 260856
rect 348142 260828 348148 260840
rect 348068 260800 348148 260828
rect 348142 260788 348148 260800
rect 348200 260788 348206 260840
rect 356440 260772 356468 260868
rect 356514 260856 356520 260868
rect 356572 260856 356578 260908
rect 381081 260899 381139 260905
rect 381081 260865 381093 260899
rect 381127 260896 381139 260899
rect 381170 260896 381176 260908
rect 381127 260868 381176 260896
rect 381127 260865 381139 260868
rect 381081 260859 381139 260865
rect 381170 260856 381176 260868
rect 381228 260856 381234 260908
rect 359001 260831 359059 260837
rect 359001 260797 359013 260831
rect 359047 260828 359059 260831
rect 359090 260828 359096 260840
rect 359047 260800 359096 260828
rect 359047 260797 359059 260800
rect 359001 260791 359059 260797
rect 359090 260788 359096 260800
rect 359148 260788 359154 260840
rect 364242 260788 364248 260840
rect 364300 260828 364306 260840
rect 364610 260828 364616 260840
rect 364300 260800 364616 260828
rect 364300 260788 364306 260800
rect 364610 260788 364616 260800
rect 364668 260788 364674 260840
rect 371418 260828 371424 260840
rect 371379 260800 371424 260828
rect 371418 260788 371424 260800
rect 371476 260788 371482 260840
rect 375561 260831 375619 260837
rect 375561 260797 375573 260831
rect 375607 260828 375619 260831
rect 375650 260828 375656 260840
rect 375607 260800 375656 260828
rect 375607 260797 375619 260800
rect 375561 260791 375619 260797
rect 375650 260788 375656 260800
rect 375708 260788 375714 260840
rect 376938 260828 376944 260840
rect 376899 260800 376944 260828
rect 376938 260788 376944 260800
rect 376996 260788 377002 260840
rect 400490 260828 400496 260840
rect 400451 260800 400496 260828
rect 400490 260788 400496 260800
rect 400548 260788 400554 260840
rect 416866 260828 416872 260840
rect 416827 260800 416872 260828
rect 416866 260788 416872 260800
rect 416924 260788 416930 260840
rect 433610 260828 433616 260840
rect 433571 260800 433616 260828
rect 433610 260788 433616 260800
rect 433668 260788 433674 260840
rect 466546 260828 466552 260840
rect 466507 260800 466552 260828
rect 466546 260788 466552 260800
rect 466604 260788 466610 260840
rect 472066 260828 472072 260840
rect 472027 260800 472072 260828
rect 472066 260788 472072 260800
rect 472124 260788 472130 260840
rect 255590 260760 255596 260772
rect 255516 260732 255596 260760
rect 255590 260720 255596 260732
rect 255648 260720 255654 260772
rect 292758 260720 292764 260772
rect 292816 260720 292822 260772
rect 309321 260763 309379 260769
rect 309321 260729 309333 260763
rect 309367 260760 309379 260763
rect 309410 260760 309416 260772
rect 309367 260732 309416 260760
rect 309367 260729 309379 260732
rect 309321 260723 309379 260729
rect 309410 260720 309416 260732
rect 309468 260720 309474 260772
rect 342441 260763 342499 260769
rect 342441 260729 342453 260763
rect 342487 260760 342499 260763
rect 342530 260760 342536 260772
rect 342487 260732 342536 260760
rect 342487 260729 342499 260732
rect 342441 260723 342499 260729
rect 342530 260720 342536 260732
rect 342588 260720 342594 260772
rect 356422 260720 356428 260772
rect 356480 260720 356486 260772
rect 397362 260720 397368 260772
rect 397420 260760 397426 260772
rect 397730 260760 397736 260772
rect 397420 260732 397736 260760
rect 397420 260720 397426 260732
rect 397730 260720 397736 260732
rect 397788 260720 397794 260772
rect 231854 259468 231860 259480
rect 231815 259440 231860 259468
rect 231854 259428 231860 259440
rect 231912 259428 231918 259480
rect 266998 259468 267004 259480
rect 266959 259440 267004 259468
rect 266998 259428 267004 259440
rect 267056 259428 267062 259480
rect 281905 259403 281963 259409
rect 281905 259369 281917 259403
rect 281951 259400 281963 259403
rect 281994 259400 282000 259412
rect 281951 259372 282000 259400
rect 281951 259369 281963 259372
rect 281905 259363 281963 259369
rect 281994 259360 282000 259372
rect 282052 259360 282058 259412
rect 295426 259400 295432 259412
rect 295387 259372 295432 259400
rect 295426 259360 295432 259372
rect 295484 259360 295490 259412
rect 451550 259400 451556 259412
rect 451511 259372 451556 259400
rect 451550 259360 451556 259372
rect 451608 259360 451614 259412
rect 292850 258000 292856 258052
rect 292908 258040 292914 258052
rect 292945 258043 293003 258049
rect 292945 258040 292957 258043
rect 292908 258012 292957 258040
rect 292908 258000 292914 258012
rect 292945 258009 292957 258012
rect 292991 258009 293003 258043
rect 292945 258003 293003 258009
rect 231854 254600 231860 254652
rect 231912 254640 231918 254652
rect 232038 254640 232044 254652
rect 231912 254612 232044 254640
rect 231912 254600 231918 254612
rect 232038 254600 232044 254612
rect 232096 254600 232102 254652
rect 348053 254643 348111 254649
rect 348053 254609 348065 254643
rect 348099 254640 348111 254643
rect 348142 254640 348148 254652
rect 348099 254612 348148 254640
rect 348099 254609 348111 254612
rect 348053 254603 348111 254609
rect 348142 254600 348148 254612
rect 348200 254600 348206 254652
rect 353573 254643 353631 254649
rect 353573 254609 353585 254643
rect 353619 254640 353631 254643
rect 353662 254640 353668 254652
rect 353619 254612 353668 254640
rect 353619 254609 353631 254612
rect 353573 254603 353631 254609
rect 353662 254600 353668 254612
rect 353720 254600 353726 254652
rect 230934 254436 230940 254448
rect 230895 254408 230940 254436
rect 230934 254396 230940 254408
rect 230992 254396 230998 254448
rect 330018 253988 330024 254040
rect 330076 253988 330082 254040
rect 356422 254028 356428 254040
rect 356383 254000 356428 254028
rect 356422 253988 356428 254000
rect 356480 253988 356486 254040
rect 357618 253988 357624 254040
rect 357676 253988 357682 254040
rect 330036 253904 330064 253988
rect 357636 253904 357664 253988
rect 236362 253892 236368 253904
rect 236288 253864 236368 253892
rect 236288 253768 236316 253864
rect 236362 253852 236368 253864
rect 236420 253852 236426 253904
rect 272058 253852 272064 253904
rect 272116 253852 272122 253904
rect 288618 253852 288624 253904
rect 288676 253852 288682 253904
rect 294138 253852 294144 253904
rect 294196 253852 294202 253904
rect 330018 253852 330024 253904
rect 330076 253852 330082 253904
rect 357618 253852 357624 253904
rect 357676 253852 357682 253904
rect 382458 253852 382464 253904
rect 382516 253852 382522 253904
rect 272076 253768 272104 253852
rect 288636 253768 288664 253852
rect 294156 253768 294184 253852
rect 382476 253768 382504 253852
rect 236270 253716 236276 253768
rect 236328 253716 236334 253768
rect 272058 253716 272064 253768
rect 272116 253716 272122 253768
rect 288618 253716 288624 253768
rect 288676 253716 288682 253768
rect 294138 253716 294144 253768
rect 294196 253716 294202 253768
rect 382458 253716 382464 253768
rect 382516 253716 382522 253768
rect 530670 252492 530676 252544
rect 530728 252532 530734 252544
rect 579614 252532 579620 252544
rect 530728 252504 579620 252532
rect 530728 252492 530734 252504
rect 579614 252492 579620 252504
rect 579672 252492 579678 252544
rect 334342 251308 334348 251320
rect 334303 251280 334348 251308
rect 334342 251268 334348 251280
rect 334400 251268 334406 251320
rect 358998 251308 359004 251320
rect 358959 251280 359004 251308
rect 358998 251268 359004 251280
rect 359056 251268 359062 251320
rect 241790 251240 241796 251252
rect 241751 251212 241796 251240
rect 241790 251200 241796 251212
rect 241848 251200 241854 251252
rect 283098 251240 283104 251252
rect 283059 251212 283104 251240
rect 283098 251200 283104 251212
rect 283156 251200 283162 251252
rect 305178 251240 305184 251252
rect 305139 251212 305184 251240
rect 305178 251200 305184 251212
rect 305236 251200 305242 251252
rect 309318 251240 309324 251252
rect 309279 251212 309324 251240
rect 309318 251200 309324 251212
rect 309376 251200 309382 251252
rect 310698 251240 310704 251252
rect 310659 251212 310704 251240
rect 310698 251200 310704 251212
rect 310756 251200 310762 251252
rect 327258 251240 327264 251252
rect 327219 251212 327264 251240
rect 327258 251200 327264 251212
rect 327316 251200 327322 251252
rect 342438 251240 342444 251252
rect 342399 251212 342444 251240
rect 342438 251200 342444 251212
rect 342496 251200 342502 251252
rect 346578 251240 346584 251252
rect 346539 251212 346584 251240
rect 346578 251200 346584 251212
rect 346636 251200 346642 251252
rect 371418 251240 371424 251252
rect 371379 251212 371424 251240
rect 371418 251200 371424 251212
rect 371476 251200 371482 251252
rect 375558 251240 375564 251252
rect 375519 251212 375564 251240
rect 375558 251200 375564 251212
rect 375616 251200 375622 251252
rect 376938 251240 376944 251252
rect 376899 251212 376944 251240
rect 376938 251200 376944 251212
rect 376996 251200 377002 251252
rect 381078 251200 381084 251252
rect 381136 251240 381142 251252
rect 381354 251240 381360 251252
rect 381136 251212 381360 251240
rect 381136 251200 381142 251212
rect 381354 251200 381360 251212
rect 381412 251200 381418 251252
rect 400493 251243 400551 251249
rect 400493 251209 400505 251243
rect 400539 251240 400551 251243
rect 400582 251240 400588 251252
rect 400539 251212 400588 251240
rect 400539 251209 400551 251212
rect 400493 251203 400551 251209
rect 400582 251200 400588 251212
rect 400640 251200 400646 251252
rect 416869 251243 416927 251249
rect 416869 251209 416881 251243
rect 416915 251240 416927 251243
rect 416958 251240 416964 251252
rect 416915 251212 416964 251240
rect 416915 251209 416927 251212
rect 416869 251203 416927 251209
rect 416958 251200 416964 251212
rect 417016 251200 417022 251252
rect 433613 251243 433671 251249
rect 433613 251209 433625 251243
rect 433659 251240 433671 251243
rect 433702 251240 433708 251252
rect 433659 251212 433708 251240
rect 433659 251209 433671 251212
rect 433613 251203 433671 251209
rect 433702 251200 433708 251212
rect 433760 251200 433766 251252
rect 466549 251243 466607 251249
rect 466549 251209 466561 251243
rect 466595 251240 466607 251243
rect 466638 251240 466644 251252
rect 466595 251212 466644 251240
rect 466595 251209 466607 251212
rect 466549 251203 466607 251209
rect 466638 251200 466644 251212
rect 466696 251200 466702 251252
rect 472069 251243 472127 251249
rect 472069 251209 472081 251243
rect 472115 251240 472127 251243
rect 472158 251240 472164 251252
rect 472115 251212 472164 251240
rect 472115 251209 472127 251212
rect 472069 251203 472127 251209
rect 472158 251200 472164 251212
rect 472216 251200 472222 251252
rect 252738 251172 252744 251184
rect 252699 251144 252744 251172
rect 252738 251132 252744 251144
rect 252796 251132 252802 251184
rect 270586 251132 270592 251184
rect 270644 251172 270650 251184
rect 270954 251172 270960 251184
rect 270644 251144 270960 251172
rect 270644 251132 270650 251144
rect 270954 251132 270960 251144
rect 271012 251132 271018 251184
rect 287238 251172 287244 251184
rect 287199 251144 287244 251172
rect 287238 251132 287244 251144
rect 287296 251132 287302 251184
rect 298189 251175 298247 251181
rect 298189 251141 298201 251175
rect 298235 251172 298247 251175
rect 298278 251172 298284 251184
rect 298235 251144 298284 251172
rect 298235 251141 298247 251144
rect 298189 251135 298247 251141
rect 298278 251132 298284 251144
rect 298336 251132 298342 251184
rect 334342 251172 334348 251184
rect 334303 251144 334348 251172
rect 334342 251132 334348 251144
rect 334400 251132 334406 251184
rect 358998 251172 359004 251184
rect 358959 251144 359004 251172
rect 358998 251132 359004 251144
rect 359056 251132 359062 251184
rect 369949 251175 370007 251181
rect 369949 251141 369961 251175
rect 369995 251172 370007 251175
rect 370038 251172 370044 251184
rect 369995 251144 370044 251172
rect 369995 251141 370007 251144
rect 369949 251135 370007 251141
rect 370038 251132 370044 251144
rect 370096 251132 370102 251184
rect 254026 251064 254032 251116
rect 254084 251104 254090 251116
rect 254210 251104 254216 251116
rect 254084 251076 254216 251104
rect 254084 251064 254090 251076
rect 254210 251064 254216 251076
rect 254268 251064 254274 251116
rect 356422 251104 356428 251116
rect 356383 251076 356428 251104
rect 356422 251064 356428 251076
rect 356480 251064 356486 251116
rect 381078 251104 381084 251116
rect 381039 251076 381084 251104
rect 381078 251064 381084 251076
rect 381136 251064 381142 251116
rect 386598 249840 386604 249892
rect 386656 249880 386662 249892
rect 386690 249880 386696 249892
rect 386656 249852 386696 249880
rect 386656 249840 386662 249852
rect 386690 249840 386696 249852
rect 386748 249840 386754 249892
rect 392118 249840 392124 249892
rect 392176 249880 392182 249892
rect 392210 249880 392216 249892
rect 392176 249852 392216 249880
rect 392176 249840 392182 249852
rect 392210 249840 392216 249852
rect 392268 249840 392274 249892
rect 259546 249772 259552 249824
rect 259604 249812 259610 249824
rect 259730 249812 259736 249824
rect 259604 249784 259736 249812
rect 259604 249772 259610 249784
rect 259730 249772 259736 249784
rect 259788 249772 259794 249824
rect 292850 249704 292856 249756
rect 292908 249744 292914 249756
rect 292945 249747 293003 249753
rect 292945 249744 292957 249747
rect 292908 249716 292957 249744
rect 292908 249704 292914 249716
rect 292945 249713 292957 249716
rect 292991 249713 293003 249747
rect 292945 249707 293003 249713
rect 324222 245420 324228 245472
rect 324280 245460 324286 245472
rect 324406 245460 324412 245472
rect 324280 245432 324412 245460
rect 324280 245420 324286 245432
rect 324406 245420 324412 245432
rect 324464 245420 324470 245472
rect 232038 244372 232044 244384
rect 231964 244344 232044 244372
rect 231964 244248 231992 244344
rect 232038 244332 232044 244344
rect 232096 244332 232102 244384
rect 233326 244264 233332 244316
rect 233384 244304 233390 244316
rect 233510 244304 233516 244316
rect 233384 244276 233516 244304
rect 233384 244264 233390 244276
rect 233510 244264 233516 244276
rect 233568 244264 233574 244316
rect 236270 244304 236276 244316
rect 236231 244276 236276 244304
rect 236270 244264 236276 244276
rect 236328 244264 236334 244316
rect 356422 244264 356428 244316
rect 356480 244264 356486 244316
rect 386690 244304 386696 244316
rect 386616 244276 386696 244304
rect 231946 244196 231952 244248
rect 232004 244196 232010 244248
rect 230934 244168 230940 244180
rect 230895 244140 230940 244168
rect 230934 244128 230940 244140
rect 230992 244128 230998 244180
rect 334342 244168 334348 244180
rect 334303 244140 334348 244168
rect 334342 244128 334348 244140
rect 334400 244128 334406 244180
rect 356440 244168 356468 244264
rect 386616 244248 386644 244276
rect 386690 244264 386696 244276
rect 386748 244264 386754 244316
rect 422294 244264 422300 244316
rect 422352 244304 422358 244316
rect 422478 244304 422484 244316
rect 422352 244276 422484 244304
rect 422352 244264 422358 244276
rect 422478 244264 422484 244276
rect 422536 244264 422542 244316
rect 427814 244264 427820 244316
rect 427872 244304 427878 244316
rect 427998 244304 428004 244316
rect 427872 244276 428004 244304
rect 427872 244264 427878 244276
rect 427998 244264 428004 244276
rect 428056 244264 428062 244316
rect 386598 244196 386604 244248
rect 386656 244196 386662 244248
rect 356514 244168 356520 244180
rect 356440 244140 356520 244168
rect 356514 244128 356520 244140
rect 356572 244128 356578 244180
rect 358998 244168 359004 244180
rect 358959 244140 359004 244168
rect 358998 244128 359004 244140
rect 359056 244128 359062 244180
rect 408770 244128 408776 244180
rect 408828 244168 408834 244180
rect 408954 244168 408960 244180
rect 408828 244140 408960 244168
rect 408828 244128 408834 244140
rect 408954 244128 408960 244140
rect 409012 244128 409018 244180
rect 451550 244168 451556 244180
rect 451511 244140 451556 244168
rect 451550 244128 451556 244140
rect 451608 244128 451614 244180
rect 298186 242672 298192 242684
rect 298147 242644 298192 242672
rect 298186 242632 298192 242644
rect 298244 242632 298250 242684
rect 364242 242156 364248 242208
rect 364300 242196 364306 242208
rect 364610 242196 364616 242208
rect 364300 242168 364616 242196
rect 364300 242156 364306 242168
rect 364610 242156 364616 242168
rect 364668 242156 364674 242208
rect 281902 241584 281908 241596
rect 281863 241556 281908 241584
rect 281902 241544 281908 241556
rect 281960 241544 281966 241596
rect 242986 241476 242992 241528
rect 243044 241516 243050 241528
rect 243170 241516 243176 241528
rect 243044 241488 243176 241516
rect 243044 241476 243050 241488
rect 243170 241476 243176 241488
rect 243228 241476 243234 241528
rect 252738 241516 252744 241528
rect 252699 241488 252744 241516
rect 252738 241476 252744 241488
rect 252796 241476 252802 241528
rect 254026 241476 254032 241528
rect 254084 241516 254090 241528
rect 254210 241516 254216 241528
rect 254084 241488 254216 241516
rect 254084 241476 254090 241488
rect 254210 241476 254216 241488
rect 254268 241476 254274 241528
rect 259546 241476 259552 241528
rect 259604 241516 259610 241528
rect 259730 241516 259736 241528
rect 259604 241488 259736 241516
rect 259604 241476 259610 241488
rect 259730 241476 259736 241488
rect 259788 241476 259794 241528
rect 287238 241516 287244 241528
rect 287199 241488 287244 241516
rect 287238 241476 287244 241488
rect 287296 241476 287302 241528
rect 309502 241476 309508 241528
rect 309560 241516 309566 241528
rect 309594 241516 309600 241528
rect 309560 241488 309600 241516
rect 309560 241476 309566 241488
rect 309594 241476 309600 241488
rect 309652 241476 309658 241528
rect 331122 241476 331128 241528
rect 331180 241516 331186 241528
rect 331490 241516 331496 241528
rect 331180 241488 331496 241516
rect 331180 241476 331186 241488
rect 331490 241476 331496 241488
rect 331548 241476 331554 241528
rect 348050 241516 348056 241528
rect 348011 241488 348056 241516
rect 348050 241476 348056 241488
rect 348108 241476 348114 241528
rect 353570 241516 353576 241528
rect 353531 241488 353576 241516
rect 353570 241476 353576 241488
rect 353628 241476 353634 241528
rect 369946 241516 369952 241528
rect 369907 241488 369952 241516
rect 369946 241476 369952 241488
rect 370004 241476 370010 241528
rect 375742 241476 375748 241528
rect 375800 241516 375806 241528
rect 375834 241516 375840 241528
rect 375800 241488 375840 241516
rect 375800 241476 375806 241488
rect 375834 241476 375840 241488
rect 375892 241476 375898 241528
rect 381081 241519 381139 241525
rect 381081 241485 381093 241519
rect 381127 241516 381139 241519
rect 381170 241516 381176 241528
rect 381127 241488 381176 241516
rect 381127 241485 381139 241488
rect 381081 241479 381139 241485
rect 381170 241476 381176 241488
rect 381228 241476 381234 241528
rect 281902 241448 281908 241460
rect 281863 241420 281908 241448
rect 281902 241408 281908 241420
rect 281960 241408 281966 241460
rect 466546 241408 466552 241460
rect 466604 241448 466610 241460
rect 466638 241448 466644 241460
rect 466604 241420 466644 241448
rect 466604 241408 466610 241420
rect 466638 241408 466644 241420
rect 466696 241408 466702 241460
rect 236270 240224 236276 240236
rect 236231 240196 236276 240224
rect 236270 240184 236276 240196
rect 236328 240184 236334 240236
rect 292758 240116 292764 240168
rect 292816 240156 292822 240168
rect 292850 240156 292856 240168
rect 292816 240128 292856 240156
rect 292816 240116 292822 240128
rect 292850 240116 292856 240128
rect 292908 240116 292914 240168
rect 392210 240116 392216 240168
rect 392268 240156 392274 240168
rect 392394 240156 392400 240168
rect 392268 240128 392400 240156
rect 392268 240116 392274 240128
rect 392394 240116 392400 240128
rect 392452 240116 392458 240168
rect 231946 240048 231952 240100
rect 232004 240088 232010 240100
rect 232222 240088 232228 240100
rect 232004 240060 232228 240088
rect 232004 240048 232010 240060
rect 232222 240048 232228 240060
rect 232280 240048 232286 240100
rect 236270 240088 236276 240100
rect 236231 240060 236276 240088
rect 236270 240048 236276 240060
rect 236328 240048 236334 240100
rect 295429 240091 295487 240097
rect 295429 240057 295441 240091
rect 295475 240088 295487 240091
rect 295518 240088 295524 240100
rect 295475 240060 295524 240088
rect 295475 240057 295487 240060
rect 295429 240051 295487 240057
rect 295518 240048 295524 240060
rect 295576 240048 295582 240100
rect 298186 240048 298192 240100
rect 298244 240088 298250 240100
rect 298278 240088 298284 240100
rect 298244 240060 298284 240088
rect 298244 240048 298250 240060
rect 298278 240048 298284 240060
rect 298336 240048 298342 240100
rect 298278 238688 298284 238740
rect 298336 238728 298342 238740
rect 298554 238728 298560 238740
rect 298336 238700 298560 238728
rect 298336 238688 298342 238700
rect 298554 238688 298560 238700
rect 298612 238688 298618 238740
rect 348050 238728 348056 238740
rect 348011 238700 348056 238728
rect 348050 238688 348056 238700
rect 348108 238688 348114 238740
rect 295518 237368 295524 237380
rect 295479 237340 295524 237368
rect 295518 237328 295524 237340
rect 295576 237328 295582 237380
rect 2774 237260 2780 237312
rect 2832 237300 2838 237312
rect 4982 237300 4988 237312
rect 2832 237272 4988 237300
rect 2832 237260 2838 237272
rect 4982 237260 4988 237272
rect 5040 237260 5046 237312
rect 392121 236759 392179 236765
rect 392121 236725 392133 236759
rect 392167 236756 392179 236759
rect 392210 236756 392216 236768
rect 392167 236728 392216 236756
rect 392167 236725 392179 236728
rect 392121 236719 392179 236725
rect 392210 236716 392216 236728
rect 392268 236716 392274 236768
rect 324222 236648 324228 236700
rect 324280 236688 324286 236700
rect 324406 236688 324412 236700
rect 324280 236660 324412 236688
rect 324280 236648 324286 236660
rect 324406 236648 324412 236660
rect 324464 236648 324470 236700
rect 364429 235943 364487 235949
rect 364429 235909 364441 235943
rect 364475 235940 364487 235943
rect 364610 235940 364616 235952
rect 364475 235912 364616 235940
rect 364475 235909 364487 235912
rect 364429 235903 364487 235909
rect 364610 235900 364616 235912
rect 364668 235900 364674 235952
rect 230934 234716 230940 234728
rect 230860 234688 230940 234716
rect 230860 234592 230888 234688
rect 230934 234676 230940 234688
rect 230992 234676 230998 234728
rect 353570 234676 353576 234728
rect 353628 234676 353634 234728
rect 356425 234719 356483 234725
rect 356425 234685 356437 234719
rect 356471 234716 356483 234719
rect 356514 234716 356520 234728
rect 356471 234688 356520 234716
rect 356471 234685 356483 234688
rect 356425 234679 356483 234685
rect 356514 234676 356520 234688
rect 356572 234676 356578 234728
rect 381078 234716 381084 234728
rect 381039 234688 381084 234716
rect 381078 234676 381084 234688
rect 381136 234676 381142 234728
rect 408770 234716 408776 234728
rect 408696 234688 408776 234716
rect 261110 234648 261116 234660
rect 261036 234620 261116 234648
rect 261036 234592 261064 234620
rect 261110 234608 261116 234620
rect 261168 234608 261174 234660
rect 327350 234648 327356 234660
rect 327276 234620 327356 234648
rect 327276 234592 327304 234620
rect 327350 234608 327356 234620
rect 327408 234608 327414 234660
rect 330110 234648 330116 234660
rect 330036 234620 330116 234648
rect 330036 234592 330064 234620
rect 330110 234608 330116 234620
rect 330168 234608 330174 234660
rect 352006 234648 352012 234660
rect 351967 234620 352012 234648
rect 352006 234608 352012 234620
rect 352064 234608 352070 234660
rect 353588 234592 353616 234676
rect 357710 234648 357716 234660
rect 357636 234620 357716 234648
rect 357636 234592 357664 234620
rect 357710 234608 357716 234620
rect 357768 234608 357774 234660
rect 408696 234592 408724 234688
rect 408770 234676 408776 234688
rect 408828 234676 408834 234728
rect 451550 234716 451556 234728
rect 451476 234688 451556 234716
rect 451476 234592 451504 234688
rect 451550 234676 451556 234688
rect 451608 234676 451614 234728
rect 230842 234540 230848 234592
rect 230900 234540 230906 234592
rect 261018 234540 261024 234592
rect 261076 234540 261082 234592
rect 272058 234540 272064 234592
rect 272116 234540 272122 234592
rect 281902 234580 281908 234592
rect 281863 234552 281908 234580
rect 281902 234540 281908 234552
rect 281960 234540 281966 234592
rect 288618 234540 288624 234592
rect 288676 234540 288682 234592
rect 294138 234540 294144 234592
rect 294196 234540 294202 234592
rect 327258 234540 327264 234592
rect 327316 234540 327322 234592
rect 330018 234540 330024 234592
rect 330076 234540 330082 234592
rect 353570 234540 353576 234592
rect 353628 234540 353634 234592
rect 357618 234540 357624 234592
rect 357676 234540 357682 234592
rect 371418 234540 371424 234592
rect 371476 234540 371482 234592
rect 382458 234540 382464 234592
rect 382516 234540 382522 234592
rect 408678 234540 408684 234592
rect 408736 234540 408742 234592
rect 451458 234540 451464 234592
rect 451516 234540 451522 234592
rect 272076 234456 272104 234540
rect 288636 234456 288664 234540
rect 294156 234456 294184 234540
rect 371436 234456 371464 234540
rect 382476 234456 382504 234540
rect 272058 234404 272064 234456
rect 272116 234404 272122 234456
rect 288618 234404 288624 234456
rect 288676 234404 288682 234456
rect 294138 234404 294144 234456
rect 294196 234404 294202 234456
rect 371418 234404 371424 234456
rect 371476 234404 371482 234456
rect 382458 234404 382464 234456
rect 382516 234404 382522 234456
rect 334342 231956 334348 232008
rect 334400 231996 334406 232008
rect 334400 231968 334480 231996
rect 334400 231956 334406 231968
rect 334452 231872 334480 231968
rect 358998 231956 359004 232008
rect 359056 231996 359062 232008
rect 359056 231968 359136 231996
rect 359056 231956 359062 231968
rect 359108 231872 359136 231968
rect 242986 231820 242992 231872
rect 243044 231860 243050 231872
rect 243078 231860 243084 231872
rect 243044 231832 243084 231860
rect 243044 231820 243050 231832
rect 243078 231820 243084 231832
rect 243136 231820 243142 231872
rect 277578 231820 277584 231872
rect 277636 231860 277642 231872
rect 277670 231860 277676 231872
rect 277636 231832 277676 231860
rect 277636 231820 277642 231832
rect 277670 231820 277676 231832
rect 277728 231820 277734 231872
rect 282914 231820 282920 231872
rect 282972 231860 282978 231872
rect 283098 231860 283104 231872
rect 282972 231832 283104 231860
rect 282972 231820 282978 231832
rect 283098 231820 283104 231832
rect 283156 231820 283162 231872
rect 305178 231820 305184 231872
rect 305236 231860 305242 231872
rect 305362 231860 305368 231872
rect 305236 231832 305368 231860
rect 305236 231820 305242 231832
rect 305362 231820 305368 231832
rect 305420 231820 305426 231872
rect 310698 231820 310704 231872
rect 310756 231860 310762 231872
rect 310882 231860 310888 231872
rect 310756 231832 310888 231860
rect 310756 231820 310762 231832
rect 310882 231820 310888 231832
rect 310940 231820 310946 231872
rect 318978 231820 318984 231872
rect 319036 231860 319042 231872
rect 319070 231860 319076 231872
rect 319036 231832 319076 231860
rect 319036 231820 319042 231832
rect 319070 231820 319076 231832
rect 319128 231820 319134 231872
rect 331490 231820 331496 231872
rect 331548 231820 331554 231872
rect 334434 231820 334440 231872
rect 334492 231820 334498 231872
rect 346578 231820 346584 231872
rect 346636 231860 346642 231872
rect 346762 231860 346768 231872
rect 346636 231832 346768 231860
rect 346636 231820 346642 231832
rect 346762 231820 346768 231832
rect 346820 231820 346826 231872
rect 359090 231820 359096 231872
rect 359148 231820 359154 231872
rect 369946 231820 369952 231872
rect 370004 231860 370010 231872
rect 370038 231860 370044 231872
rect 370004 231832 370044 231860
rect 370004 231820 370010 231832
rect 370038 231820 370044 231832
rect 370096 231820 370102 231872
rect 375558 231820 375564 231872
rect 375616 231860 375622 231872
rect 375834 231860 375840 231872
rect 375616 231832 375840 231860
rect 375616 231820 375622 231832
rect 375834 231820 375840 231832
rect 375892 231820 375898 231872
rect 376754 231820 376760 231872
rect 376812 231860 376818 231872
rect 376938 231860 376944 231872
rect 376812 231832 376944 231860
rect 376812 231820 376818 231832
rect 376938 231820 376944 231832
rect 376996 231820 377002 231872
rect 381081 231863 381139 231869
rect 381081 231829 381093 231863
rect 381127 231860 381139 231863
rect 381170 231860 381176 231872
rect 381127 231832 381176 231860
rect 381127 231829 381139 231832
rect 381081 231823 381139 231829
rect 381170 231820 381176 231832
rect 381228 231820 381234 231872
rect 393130 231820 393136 231872
rect 393188 231860 393194 231872
rect 393222 231860 393228 231872
rect 393188 231832 393228 231860
rect 393188 231820 393194 231832
rect 393222 231820 393228 231832
rect 393280 231820 393286 231872
rect 397730 231820 397736 231872
rect 397788 231860 397794 231872
rect 397914 231860 397920 231872
rect 397788 231832 397920 231860
rect 397788 231820 397794 231832
rect 397914 231820 397920 231832
rect 397972 231820 397978 231872
rect 400306 231820 400312 231872
rect 400364 231860 400370 231872
rect 400582 231860 400588 231872
rect 400364 231832 400588 231860
rect 400364 231820 400370 231832
rect 400582 231820 400588 231832
rect 400640 231820 400646 231872
rect 416958 231820 416964 231872
rect 417016 231860 417022 231872
rect 417142 231860 417148 231872
rect 417016 231832 417148 231860
rect 417016 231820 417022 231832
rect 417142 231820 417148 231832
rect 417200 231820 417206 231872
rect 433426 231820 433432 231872
rect 433484 231860 433490 231872
rect 433702 231860 433708 231872
rect 433484 231832 433708 231860
rect 433484 231820 433490 231832
rect 433702 231820 433708 231832
rect 433760 231820 433766 231872
rect 472158 231820 472164 231872
rect 472216 231860 472222 231872
rect 472342 231860 472348 231872
rect 472216 231832 472348 231860
rect 472216 231820 472222 231832
rect 472342 231820 472348 231832
rect 472400 231820 472406 231872
rect 259638 231792 259644 231804
rect 259599 231764 259644 231792
rect 259638 231752 259644 231764
rect 259696 231752 259702 231804
rect 331508 231736 331536 231820
rect 408678 231792 408684 231804
rect 408639 231764 408684 231792
rect 408678 231752 408684 231764
rect 408736 231752 408742 231804
rect 243170 231724 243176 231736
rect 243131 231696 243176 231724
rect 243170 231684 243176 231696
rect 243228 231684 243234 231736
rect 331490 231684 331496 231736
rect 331548 231684 331554 231736
rect 236270 230568 236276 230580
rect 236231 230540 236276 230568
rect 236270 230528 236276 230540
rect 236328 230528 236334 230580
rect 265158 230528 265164 230580
rect 265216 230568 265222 230580
rect 265250 230568 265256 230580
rect 265216 230540 265256 230568
rect 265216 230528 265222 230540
rect 265250 230528 265256 230540
rect 265308 230528 265314 230580
rect 292758 230528 292764 230580
rect 292816 230568 292822 230580
rect 292850 230568 292856 230580
rect 292816 230540 292856 230568
rect 292816 230528 292822 230540
rect 292850 230528 292856 230540
rect 292908 230528 292914 230580
rect 348050 230364 348056 230376
rect 348011 230336 348056 230364
rect 348050 230324 348056 230336
rect 348108 230324 348114 230376
rect 352009 230367 352067 230373
rect 352009 230333 352021 230367
rect 352055 230364 352067 230367
rect 352190 230364 352196 230376
rect 352055 230336 352196 230364
rect 352055 230333 352067 230336
rect 352009 230327 352067 230333
rect 352190 230324 352196 230336
rect 352248 230324 352254 230376
rect 356422 229208 356428 229220
rect 356383 229180 356428 229208
rect 356422 229168 356428 229180
rect 356480 229168 356486 229220
rect 356422 229072 356428 229084
rect 356383 229044 356428 229072
rect 356422 229032 356428 229044
rect 356480 229032 356486 229084
rect 295518 227780 295524 227792
rect 295479 227752 295524 227780
rect 295518 227740 295524 227752
rect 295576 227740 295582 227792
rect 233326 224952 233332 225004
rect 233384 224992 233390 225004
rect 233510 224992 233516 225004
rect 233384 224964 233516 224992
rect 233384 224952 233390 224964
rect 233510 224952 233516 224964
rect 233568 224952 233574 225004
rect 254118 224952 254124 225004
rect 254176 224952 254182 225004
rect 267090 224992 267096 225004
rect 267051 224964 267096 224992
rect 267090 224952 267096 224964
rect 267148 224952 267154 225004
rect 295518 224952 295524 225004
rect 295576 224952 295582 225004
rect 309318 224952 309324 225004
rect 309376 224952 309382 225004
rect 324406 224992 324412 225004
rect 324367 224964 324412 224992
rect 324406 224952 324412 224964
rect 324464 224952 324470 225004
rect 381170 224992 381176 225004
rect 381131 224964 381176 224992
rect 381170 224952 381176 224964
rect 381228 224952 381234 225004
rect 386598 224952 386604 225004
rect 386656 224952 386662 225004
rect 397730 224952 397736 225004
rect 397788 224952 397794 225004
rect 422294 224952 422300 225004
rect 422352 224992 422358 225004
rect 422478 224992 422484 225004
rect 422352 224964 422484 224992
rect 422352 224952 422358 224964
rect 422478 224952 422484 224964
rect 422536 224952 422542 225004
rect 427814 224952 427820 225004
rect 427872 224992 427878 225004
rect 427998 224992 428004 225004
rect 427872 224964 428004 224992
rect 427872 224952 427878 224964
rect 427998 224952 428004 224964
rect 428056 224952 428062 225004
rect 254136 224856 254164 224952
rect 254210 224856 254216 224868
rect 254136 224828 254216 224856
rect 254210 224816 254216 224828
rect 254268 224816 254274 224868
rect 265158 224816 265164 224868
rect 265216 224856 265222 224868
rect 265342 224856 265348 224868
rect 265216 224828 265348 224856
rect 265216 224816 265222 224828
rect 265342 224816 265348 224828
rect 265400 224816 265406 224868
rect 295536 224856 295564 224952
rect 295610 224856 295616 224868
rect 295536 224828 295616 224856
rect 295610 224816 295616 224828
rect 295668 224816 295674 224868
rect 309336 224856 309364 224952
rect 356422 224924 356428 224936
rect 356383 224896 356428 224924
rect 356422 224884 356428 224896
rect 356480 224884 356486 224936
rect 309410 224856 309416 224868
rect 309336 224828 309416 224856
rect 309410 224816 309416 224828
rect 309468 224816 309474 224868
rect 386616 224856 386644 224952
rect 397748 224868 397776 224952
rect 386690 224856 386696 224868
rect 386616 224828 386696 224856
rect 386690 224816 386696 224828
rect 386748 224816 386754 224868
rect 397730 224816 397736 224868
rect 397788 224816 397794 224868
rect 243173 224247 243231 224253
rect 243173 224213 243185 224247
rect 243219 224244 243231 224247
rect 243354 224244 243360 224256
rect 243219 224216 243360 224244
rect 243219 224213 243231 224216
rect 243173 224207 243231 224213
rect 243354 224204 243360 224216
rect 243412 224204 243418 224256
rect 231946 222232 231952 222284
rect 232004 222272 232010 222284
rect 232222 222272 232228 222284
rect 232004 222244 232228 222272
rect 232004 222232 232010 222244
rect 232222 222232 232228 222244
rect 232280 222232 232286 222284
rect 324406 222272 324412 222284
rect 324367 222244 324412 222272
rect 324406 222232 324412 222244
rect 324464 222232 324470 222284
rect 230658 222164 230664 222216
rect 230716 222204 230722 222216
rect 230934 222204 230940 222216
rect 230716 222176 230940 222204
rect 230716 222164 230722 222176
rect 230934 222164 230940 222176
rect 230992 222164 230998 222216
rect 252738 222164 252744 222216
rect 252796 222204 252802 222216
rect 252922 222204 252928 222216
rect 252796 222176 252928 222204
rect 252796 222164 252802 222176
rect 252922 222164 252928 222176
rect 252980 222164 252986 222216
rect 259641 222207 259699 222213
rect 259641 222173 259653 222207
rect 259687 222204 259699 222207
rect 259730 222204 259736 222216
rect 259687 222176 259736 222204
rect 259687 222173 259699 222176
rect 259641 222167 259699 222173
rect 259730 222164 259736 222176
rect 259788 222164 259794 222216
rect 281902 222204 281908 222216
rect 281863 222176 281908 222204
rect 281902 222164 281908 222176
rect 281960 222164 281966 222216
rect 287238 222164 287244 222216
rect 287296 222204 287302 222216
rect 287422 222204 287428 222216
rect 287296 222176 287428 222204
rect 287296 222164 287302 222176
rect 287422 222164 287428 222176
rect 287480 222164 287486 222216
rect 381170 222204 381176 222216
rect 381131 222176 381176 222204
rect 381170 222164 381176 222176
rect 381228 222164 381234 222216
rect 392121 222207 392179 222213
rect 392121 222173 392133 222207
rect 392167 222204 392179 222207
rect 392210 222204 392216 222216
rect 392167 222176 392216 222204
rect 392167 222173 392179 222176
rect 392121 222167 392179 222173
rect 392210 222164 392216 222176
rect 392268 222164 392274 222216
rect 393222 222164 393228 222216
rect 393280 222204 393286 222216
rect 393406 222204 393412 222216
rect 393280 222176 393412 222204
rect 393280 222164 393286 222176
rect 393406 222164 393412 222176
rect 393464 222164 393470 222216
rect 408681 222207 408739 222213
rect 408681 222173 408693 222207
rect 408727 222204 408739 222207
rect 408770 222204 408776 222216
rect 408727 222176 408776 222204
rect 408727 222173 408739 222176
rect 408681 222167 408739 222173
rect 408770 222164 408776 222176
rect 408828 222164 408834 222216
rect 451274 222164 451280 222216
rect 451332 222204 451338 222216
rect 451550 222204 451556 222216
rect 451332 222176 451556 222204
rect 451332 222164 451338 222176
rect 451550 222164 451556 222176
rect 451608 222164 451614 222216
rect 324406 222136 324412 222148
rect 324367 222108 324412 222136
rect 324406 222096 324412 222108
rect 324464 222096 324470 222148
rect 466546 222096 466552 222148
rect 466604 222136 466610 222148
rect 466638 222136 466644 222148
rect 466604 222108 466644 222136
rect 466604 222096 466610 222108
rect 466638 222096 466644 222108
rect 466696 222096 466702 222148
rect 236270 220804 236276 220856
rect 236328 220844 236334 220856
rect 236454 220844 236460 220856
rect 236328 220816 236460 220844
rect 236328 220804 236334 220816
rect 236454 220804 236460 220816
rect 236512 220804 236518 220856
rect 267090 220844 267096 220856
rect 267051 220816 267096 220844
rect 267090 220804 267096 220816
rect 267148 220804 267154 220856
rect 281902 220844 281908 220856
rect 281863 220816 281908 220844
rect 281902 220804 281908 220816
rect 281960 220804 281966 220856
rect 298370 220804 298376 220856
rect 298428 220844 298434 220856
rect 298554 220844 298560 220856
rect 298428 220816 298560 220844
rect 298428 220804 298434 220816
rect 298554 220804 298560 220816
rect 298612 220804 298618 220856
rect 331306 220804 331312 220856
rect 331364 220844 331370 220856
rect 331582 220844 331588 220856
rect 331364 220816 331588 220844
rect 331364 220804 331370 220816
rect 331582 220804 331588 220816
rect 331640 220804 331646 220856
rect 352006 220804 352012 220856
rect 352064 220844 352070 220856
rect 352190 220844 352196 220856
rect 352064 220816 352196 220844
rect 352064 220804 352070 220816
rect 352190 220804 352196 220816
rect 352248 220804 352254 220856
rect 324406 219552 324412 219564
rect 324367 219524 324412 219552
rect 324406 219512 324412 219524
rect 324464 219512 324470 219564
rect 243078 219376 243084 219428
rect 243136 219416 243142 219428
rect 243354 219416 243360 219428
rect 243136 219388 243360 219416
rect 243136 219376 243142 219388
rect 243354 219376 243360 219388
rect 243412 219376 243418 219428
rect 267001 219419 267059 219425
rect 267001 219385 267013 219419
rect 267047 219416 267059 219419
rect 267090 219416 267096 219428
rect 267047 219388 267096 219416
rect 267047 219385 267059 219388
rect 267001 219379 267059 219385
rect 267090 219376 267096 219388
rect 267148 219376 267154 219428
rect 331122 219376 331128 219428
rect 331180 219416 331186 219428
rect 331306 219416 331312 219428
rect 331180 219388 331312 219416
rect 331180 219376 331186 219388
rect 331306 219376 331312 219388
rect 331364 219376 331370 219428
rect 364426 218056 364432 218068
rect 364387 218028 364432 218056
rect 364426 218016 364432 218028
rect 364484 218016 364490 218068
rect 243078 217988 243084 218000
rect 243039 217960 243084 217988
rect 243078 217948 243084 217960
rect 243136 217948 243142 218000
rect 577498 217948 577504 218000
rect 577556 217988 577562 218000
rect 579614 217988 579620 218000
rect 577556 217960 579620 217988
rect 577556 217948 577562 217960
rect 579614 217948 579620 217960
rect 579672 217948 579678 218000
rect 254210 217444 254216 217456
rect 254136 217416 254216 217444
rect 254136 217388 254164 217416
rect 254210 217404 254216 217416
rect 254268 217404 254274 217456
rect 259730 217444 259736 217456
rect 259656 217416 259736 217444
rect 259656 217388 259684 217416
rect 259730 217404 259736 217416
rect 259788 217404 259794 217456
rect 254118 217336 254124 217388
rect 254176 217336 254182 217388
rect 259638 217336 259644 217388
rect 259696 217336 259702 217388
rect 236362 215976 236368 216028
rect 236420 216016 236426 216028
rect 236546 216016 236552 216028
rect 236420 215988 236552 216016
rect 236420 215976 236426 215988
rect 236546 215976 236552 215988
rect 236604 215976 236610 216028
rect 298281 215475 298339 215481
rect 298281 215441 298293 215475
rect 298327 215472 298339 215475
rect 298370 215472 298376 215484
rect 298327 215444 298376 215472
rect 298327 215441 298339 215444
rect 298281 215435 298339 215441
rect 298370 215432 298376 215444
rect 298428 215432 298434 215484
rect 230934 215404 230940 215416
rect 230860 215376 230940 215404
rect 230860 215280 230888 215376
rect 230934 215364 230940 215376
rect 230992 215364 230998 215416
rect 281902 215364 281908 215416
rect 281960 215364 281966 215416
rect 295429 215407 295487 215413
rect 295429 215373 295441 215407
rect 295475 215404 295487 215407
rect 295610 215404 295616 215416
rect 295475 215376 295616 215404
rect 295475 215373 295487 215376
rect 295429 215367 295487 215373
rect 295610 215364 295616 215376
rect 295668 215364 295674 215416
rect 370038 215364 370044 215416
rect 370096 215364 370102 215416
rect 381078 215404 381084 215416
rect 381039 215376 381084 215404
rect 381078 215364 381084 215376
rect 381136 215364 381142 215416
rect 408770 215404 408776 215416
rect 408696 215376 408776 215404
rect 281920 215280 281948 215364
rect 309318 215336 309324 215348
rect 309279 215308 309324 215336
rect 309318 215296 309324 215308
rect 309376 215296 309382 215348
rect 327350 215336 327356 215348
rect 327276 215308 327356 215336
rect 327276 215280 327304 215308
rect 327350 215296 327356 215308
rect 327408 215296 327414 215348
rect 330110 215336 330116 215348
rect 330036 215308 330116 215336
rect 330036 215280 330064 215308
rect 330110 215296 330116 215308
rect 330168 215296 330174 215348
rect 357710 215336 357716 215348
rect 357636 215308 357716 215336
rect 357636 215280 357664 215308
rect 357710 215296 357716 215308
rect 357768 215296 357774 215348
rect 370056 215280 370084 215364
rect 397638 215336 397644 215348
rect 397599 215308 397644 215336
rect 397638 215296 397644 215308
rect 397696 215296 397702 215348
rect 408696 215280 408724 215376
rect 408770 215364 408776 215376
rect 408828 215364 408834 215416
rect 451550 215404 451556 215416
rect 451476 215376 451556 215404
rect 451476 215280 451504 215376
rect 451550 215364 451556 215376
rect 451608 215364 451614 215416
rect 230842 215228 230848 215280
rect 230900 215228 230906 215280
rect 231762 215228 231768 215280
rect 231820 215268 231826 215280
rect 231946 215268 231952 215280
rect 231820 215240 231952 215268
rect 231820 215228 231826 215240
rect 231946 215228 231952 215240
rect 232004 215228 232010 215280
rect 233326 215228 233332 215280
rect 233384 215268 233390 215280
rect 233510 215268 233516 215280
rect 233384 215240 233516 215268
rect 233384 215228 233390 215240
rect 233510 215228 233516 215240
rect 233568 215228 233574 215280
rect 272058 215228 272064 215280
rect 272116 215228 272122 215280
rect 281902 215228 281908 215280
rect 281960 215228 281966 215280
rect 327258 215228 327264 215280
rect 327316 215228 327322 215280
rect 330018 215228 330024 215280
rect 330076 215228 330082 215280
rect 357618 215228 357624 215280
rect 357676 215228 357682 215280
rect 370038 215228 370044 215280
rect 370096 215228 370102 215280
rect 371418 215228 371424 215280
rect 371476 215228 371482 215280
rect 382458 215228 382464 215280
rect 382516 215228 382522 215280
rect 408678 215228 408684 215280
rect 408736 215228 408742 215280
rect 451458 215228 451464 215280
rect 451516 215228 451522 215280
rect 272076 215144 272104 215228
rect 371436 215144 371464 215228
rect 382476 215144 382504 215228
rect 272058 215092 272064 215144
rect 272116 215092 272122 215144
rect 371418 215092 371424 215144
rect 371476 215092 371482 215144
rect 382458 215092 382464 215144
rect 382516 215092 382522 215144
rect 334342 212644 334348 212696
rect 334400 212684 334406 212696
rect 334400 212656 334480 212684
rect 334400 212644 334406 212656
rect 334452 212560 334480 212656
rect 356514 212616 356520 212628
rect 356440 212588 356520 212616
rect 356440 212560 356468 212588
rect 356514 212576 356520 212588
rect 356572 212576 356578 212628
rect 358909 212619 358967 212625
rect 358909 212585 358921 212619
rect 358955 212616 358967 212619
rect 358998 212616 359004 212628
rect 358955 212588 359004 212616
rect 358955 212585 358967 212588
rect 358909 212579 358967 212585
rect 358998 212576 359004 212588
rect 359056 212576 359062 212628
rect 252738 212508 252744 212560
rect 252796 212548 252802 212560
rect 252830 212548 252836 212560
rect 252796 212520 252836 212548
rect 252796 212508 252802 212520
rect 252830 212508 252836 212520
rect 252888 212508 252894 212560
rect 270770 212508 270776 212560
rect 270828 212548 270834 212560
rect 270954 212548 270960 212560
rect 270828 212520 270960 212548
rect 270828 212508 270834 212520
rect 270954 212508 270960 212520
rect 271012 212508 271018 212560
rect 277578 212508 277584 212560
rect 277636 212548 277642 212560
rect 277670 212548 277676 212560
rect 277636 212520 277676 212548
rect 277636 212508 277642 212520
rect 277670 212508 277676 212520
rect 277728 212508 277734 212560
rect 305178 212508 305184 212560
rect 305236 212548 305242 212560
rect 305362 212548 305368 212560
rect 305236 212520 305368 212548
rect 305236 212508 305242 212520
rect 305362 212508 305368 212520
rect 305420 212508 305426 212560
rect 309321 212551 309379 212557
rect 309321 212517 309333 212551
rect 309367 212548 309379 212551
rect 309410 212548 309416 212560
rect 309367 212520 309416 212548
rect 309367 212517 309379 212520
rect 309321 212511 309379 212517
rect 309410 212508 309416 212520
rect 309468 212508 309474 212560
rect 310698 212508 310704 212560
rect 310756 212548 310762 212560
rect 310882 212548 310888 212560
rect 310756 212520 310888 212548
rect 310756 212508 310762 212520
rect 310882 212508 310888 212520
rect 310940 212508 310946 212560
rect 318978 212508 318984 212560
rect 319036 212548 319042 212560
rect 319070 212548 319076 212560
rect 319036 212520 319076 212548
rect 319036 212508 319042 212520
rect 319070 212508 319076 212520
rect 319128 212508 319134 212560
rect 334434 212508 334440 212560
rect 334492 212508 334498 212560
rect 346578 212508 346584 212560
rect 346636 212548 346642 212560
rect 346762 212548 346768 212560
rect 346636 212520 346768 212548
rect 346636 212508 346642 212520
rect 346762 212508 346768 212520
rect 346820 212508 346826 212560
rect 347958 212508 347964 212560
rect 348016 212548 348022 212560
rect 348142 212548 348148 212560
rect 348016 212520 348148 212548
rect 348016 212508 348022 212520
rect 348142 212508 348148 212520
rect 348200 212508 348206 212560
rect 352006 212508 352012 212560
rect 352064 212548 352070 212560
rect 352098 212548 352104 212560
rect 352064 212520 352104 212548
rect 352064 212508 352070 212520
rect 352098 212508 352104 212520
rect 352156 212508 352162 212560
rect 353478 212508 353484 212560
rect 353536 212548 353542 212560
rect 353662 212548 353668 212560
rect 353536 212520 353668 212548
rect 353536 212508 353542 212520
rect 353662 212508 353668 212520
rect 353720 212508 353726 212560
rect 356422 212508 356428 212560
rect 356480 212508 356486 212560
rect 375558 212508 375564 212560
rect 375616 212548 375622 212560
rect 375834 212548 375840 212560
rect 375616 212520 375840 212548
rect 375616 212508 375622 212520
rect 375834 212508 375840 212520
rect 375892 212508 375898 212560
rect 376754 212508 376760 212560
rect 376812 212548 376818 212560
rect 376938 212548 376944 212560
rect 376812 212520 376944 212548
rect 376812 212508 376818 212520
rect 376938 212508 376944 212520
rect 376996 212508 377002 212560
rect 381081 212551 381139 212557
rect 381081 212517 381093 212551
rect 381127 212548 381139 212551
rect 381170 212548 381176 212560
rect 381127 212520 381176 212548
rect 381127 212517 381139 212520
rect 381081 212511 381139 212517
rect 381170 212508 381176 212520
rect 381228 212508 381234 212560
rect 393130 212508 393136 212560
rect 393188 212548 393194 212560
rect 393222 212548 393228 212560
rect 393188 212520 393228 212548
rect 393188 212508 393194 212520
rect 393222 212508 393228 212520
rect 393280 212508 393286 212560
rect 397546 212508 397552 212560
rect 397604 212548 397610 212560
rect 397641 212551 397699 212557
rect 397641 212548 397653 212551
rect 397604 212520 397653 212548
rect 397604 212508 397610 212520
rect 397641 212517 397653 212520
rect 397687 212517 397699 212551
rect 397641 212511 397699 212517
rect 400306 212508 400312 212560
rect 400364 212548 400370 212560
rect 400582 212548 400588 212560
rect 400364 212520 400588 212548
rect 400364 212508 400370 212520
rect 400582 212508 400588 212520
rect 400640 212508 400646 212560
rect 416958 212508 416964 212560
rect 417016 212548 417022 212560
rect 417142 212548 417148 212560
rect 417016 212520 417148 212548
rect 417016 212508 417022 212520
rect 417142 212508 417148 212520
rect 417200 212508 417206 212560
rect 433426 212508 433432 212560
rect 433484 212548 433490 212560
rect 433702 212548 433708 212560
rect 433484 212520 433708 212548
rect 433484 212508 433490 212520
rect 433702 212508 433708 212520
rect 433760 212508 433766 212560
rect 472158 212508 472164 212560
rect 472216 212548 472222 212560
rect 472342 212548 472348 212560
rect 472216 212520 472348 212548
rect 472216 212508 472222 212520
rect 472342 212508 472348 212520
rect 472400 212508 472406 212560
rect 408678 212480 408684 212492
rect 408639 212452 408684 212480
rect 408678 212440 408684 212452
rect 408736 212440 408742 212492
rect 298278 211256 298284 211268
rect 298239 211228 298284 211256
rect 298278 211216 298284 211228
rect 298336 211216 298342 211268
rect 281718 211120 281724 211132
rect 281679 211092 281724 211120
rect 281718 211080 281724 211092
rect 281776 211080 281782 211132
rect 295426 211120 295432 211132
rect 295387 211092 295432 211120
rect 295426 211080 295432 211092
rect 295484 211080 295490 211132
rect 298278 211120 298284 211132
rect 298239 211092 298284 211120
rect 298278 211080 298284 211092
rect 298336 211080 298342 211132
rect 356422 211120 356428 211132
rect 356383 211092 356428 211120
rect 356422 211080 356428 211092
rect 356480 211080 356486 211132
rect 370038 211080 370044 211132
rect 370096 211120 370102 211132
rect 370222 211120 370228 211132
rect 370096 211092 370228 211120
rect 370096 211080 370102 211092
rect 370222 211080 370228 211092
rect 370280 211080 370286 211132
rect 266998 209828 267004 209840
rect 266959 209800 267004 209828
rect 266998 209788 267004 209800
rect 267056 209788 267062 209840
rect 265158 209760 265164 209772
rect 265119 209732 265164 209760
rect 265158 209720 265164 209732
rect 265216 209720 265222 209772
rect 358906 208400 358912 208412
rect 358867 208372 358912 208400
rect 358906 208360 358912 208372
rect 358964 208360 358970 208412
rect 295426 206252 295432 206304
rect 295484 206292 295490 206304
rect 295702 206292 295708 206304
rect 295484 206264 295708 206292
rect 295484 206252 295490 206264
rect 295702 206252 295708 206264
rect 295760 206252 295766 206304
rect 259638 205640 259644 205692
rect 259696 205640 259702 205692
rect 309410 205680 309416 205692
rect 309371 205652 309416 205680
rect 309410 205640 309416 205652
rect 309468 205640 309474 205692
rect 324406 205680 324412 205692
rect 324367 205652 324412 205680
rect 324406 205640 324412 205652
rect 324464 205640 324470 205692
rect 347958 205640 347964 205692
rect 348016 205640 348022 205692
rect 353478 205640 353484 205692
rect 353536 205640 353542 205692
rect 381170 205640 381176 205692
rect 381228 205640 381234 205692
rect 422294 205640 422300 205692
rect 422352 205680 422358 205692
rect 422478 205680 422484 205692
rect 422352 205652 422484 205680
rect 422352 205640 422358 205652
rect 422478 205640 422484 205652
rect 422536 205640 422542 205692
rect 427814 205640 427820 205692
rect 427872 205680 427878 205692
rect 427998 205680 428004 205692
rect 427872 205652 428004 205680
rect 427872 205640 427878 205652
rect 427998 205640 428004 205652
rect 428056 205640 428062 205692
rect 236270 205612 236276 205624
rect 236231 205584 236276 205612
rect 236270 205572 236276 205584
rect 236328 205572 236334 205624
rect 259656 205544 259684 205640
rect 298278 205612 298284 205624
rect 298239 205584 298284 205612
rect 298278 205572 298284 205584
rect 298336 205572 298342 205624
rect 259730 205544 259736 205556
rect 259656 205516 259736 205544
rect 259730 205504 259736 205516
rect 259788 205504 259794 205556
rect 347976 205544 348004 205640
rect 353496 205612 353524 205640
rect 353570 205612 353576 205624
rect 353496 205584 353576 205612
rect 353570 205572 353576 205584
rect 353628 205572 353634 205624
rect 381188 205556 381216 205640
rect 530578 205572 530584 205624
rect 530636 205612 530642 205624
rect 580166 205612 580172 205624
rect 530636 205584 580172 205612
rect 530636 205572 530642 205584
rect 580166 205572 580172 205584
rect 580224 205572 580230 205624
rect 348050 205544 348056 205556
rect 347976 205516 348056 205544
rect 348050 205504 348056 205516
rect 348108 205504 348114 205556
rect 381170 205504 381176 205556
rect 381228 205504 381234 205556
rect 233510 205164 233516 205216
rect 233568 205164 233574 205216
rect 233528 205080 233556 205164
rect 233510 205028 233516 205080
rect 233568 205028 233574 205080
rect 331401 202963 331459 202969
rect 331401 202929 331413 202963
rect 331447 202960 331459 202963
rect 331490 202960 331496 202972
rect 331447 202932 331496 202960
rect 331447 202929 331459 202932
rect 331401 202923 331459 202929
rect 331490 202920 331496 202932
rect 331548 202920 331554 202972
rect 230658 202852 230664 202904
rect 230716 202892 230722 202904
rect 230934 202892 230940 202904
rect 230716 202864 230940 202892
rect 230716 202852 230722 202864
rect 230934 202852 230940 202864
rect 230992 202852 230998 202904
rect 231946 202852 231952 202904
rect 232004 202892 232010 202904
rect 232038 202892 232044 202904
rect 232004 202864 232044 202892
rect 232004 202852 232010 202864
rect 232038 202852 232044 202864
rect 232096 202852 232102 202904
rect 236270 202892 236276 202904
rect 236231 202864 236276 202892
rect 236270 202852 236276 202864
rect 236328 202852 236334 202904
rect 252462 202852 252468 202904
rect 252520 202892 252526 202904
rect 252554 202892 252560 202904
rect 252520 202864 252560 202892
rect 252520 202852 252526 202864
rect 252554 202852 252560 202864
rect 252612 202852 252618 202904
rect 309410 202892 309416 202904
rect 309371 202864 309416 202892
rect 309410 202852 309416 202864
rect 309468 202852 309474 202904
rect 324406 202892 324412 202904
rect 324367 202864 324412 202892
rect 324406 202852 324412 202864
rect 324464 202852 324470 202904
rect 342622 202852 342628 202904
rect 342680 202892 342686 202904
rect 342714 202892 342720 202904
rect 342680 202864 342720 202892
rect 342680 202852 342686 202864
rect 342714 202852 342720 202864
rect 342772 202852 342778 202904
rect 352006 202852 352012 202904
rect 352064 202892 352070 202904
rect 352098 202892 352104 202904
rect 352064 202864 352104 202892
rect 352064 202852 352070 202864
rect 352098 202852 352104 202864
rect 352156 202852 352162 202904
rect 393222 202852 393228 202904
rect 393280 202892 393286 202904
rect 393406 202892 393412 202904
rect 393280 202864 393412 202892
rect 393280 202852 393286 202864
rect 393406 202852 393412 202864
rect 393464 202852 393470 202904
rect 397362 202852 397368 202904
rect 397420 202892 397426 202904
rect 397730 202892 397736 202904
rect 397420 202864 397736 202892
rect 397420 202852 397426 202864
rect 397730 202852 397736 202864
rect 397788 202852 397794 202904
rect 408681 202895 408739 202901
rect 408681 202861 408693 202895
rect 408727 202892 408739 202895
rect 408770 202892 408776 202904
rect 408727 202864 408776 202892
rect 408727 202861 408739 202864
rect 408681 202855 408739 202861
rect 408770 202852 408776 202864
rect 408828 202852 408834 202904
rect 451274 202852 451280 202904
rect 451332 202892 451338 202904
rect 451550 202892 451556 202904
rect 451332 202864 451556 202892
rect 451332 202852 451338 202864
rect 451550 202852 451556 202864
rect 451608 202852 451614 202904
rect 265161 202827 265219 202833
rect 265161 202793 265173 202827
rect 265207 202824 265219 202827
rect 265250 202824 265256 202836
rect 265207 202796 265256 202824
rect 265207 202793 265219 202796
rect 265161 202787 265219 202793
rect 265250 202784 265256 202796
rect 265308 202784 265314 202836
rect 281721 202827 281779 202833
rect 281721 202793 281733 202827
rect 281767 202824 281779 202827
rect 281810 202824 281816 202836
rect 281767 202796 281816 202824
rect 281767 202793 281779 202796
rect 281721 202787 281779 202793
rect 281810 202784 281816 202796
rect 281868 202784 281874 202836
rect 356422 202824 356428 202836
rect 356383 202796 356428 202824
rect 356422 202784 356428 202796
rect 356480 202784 356486 202836
rect 466546 202784 466552 202836
rect 466604 202824 466610 202836
rect 466638 202824 466644 202836
rect 466604 202796 466644 202824
rect 466604 202784 466610 202796
rect 466638 202784 466644 202796
rect 466696 202784 466702 202836
rect 331398 201532 331404 201544
rect 331359 201504 331404 201532
rect 331398 201492 331404 201504
rect 331456 201492 331462 201544
rect 243078 201464 243084 201476
rect 243039 201436 243084 201464
rect 243078 201424 243084 201436
rect 243136 201424 243142 201476
rect 375558 201424 375564 201476
rect 375616 201464 375622 201476
rect 375834 201464 375840 201476
rect 375616 201436 375840 201464
rect 375616 201424 375622 201436
rect 375834 201424 375840 201436
rect 375892 201424 375898 201476
rect 381078 201424 381084 201476
rect 381136 201464 381142 201476
rect 381354 201464 381360 201476
rect 381136 201436 381360 201464
rect 381136 201424 381142 201436
rect 381354 201424 381360 201436
rect 381412 201424 381418 201476
rect 292758 200064 292764 200116
rect 292816 200104 292822 200116
rect 292850 200104 292856 200116
rect 292816 200076 292856 200104
rect 292816 200064 292822 200076
rect 292850 200064 292856 200076
rect 292908 200064 292914 200116
rect 295426 200064 295432 200116
rect 295484 200104 295490 200116
rect 295702 200104 295708 200116
rect 295484 200076 295708 200104
rect 295484 200064 295490 200076
rect 295702 200064 295708 200076
rect 295760 200064 295766 200116
rect 236270 198676 236276 198688
rect 236231 198648 236276 198676
rect 236270 198636 236276 198648
rect 236328 198636 236334 198688
rect 292761 198679 292819 198685
rect 292761 198645 292773 198679
rect 292807 198676 292819 198679
rect 292850 198676 292856 198688
rect 292807 198648 292856 198676
rect 292807 198645 292819 198648
rect 292761 198639 292819 198645
rect 292850 198636 292856 198648
rect 292908 198636 292914 198688
rect 331030 196596 331036 196648
rect 331088 196636 331094 196648
rect 331398 196636 331404 196648
rect 331088 196608 331404 196636
rect 331088 196596 331094 196608
rect 331398 196596 331404 196608
rect 331456 196596 331462 196648
rect 342714 196596 342720 196648
rect 342772 196636 342778 196648
rect 342898 196636 342904 196648
rect 342772 196608 342904 196636
rect 342772 196596 342778 196608
rect 342898 196596 342904 196608
rect 342956 196596 342962 196648
rect 230934 196092 230940 196104
rect 230860 196064 230940 196092
rect 230860 195968 230888 196064
rect 230934 196052 230940 196064
rect 230992 196052 230998 196104
rect 243170 196052 243176 196104
rect 243228 196052 243234 196104
rect 270770 196092 270776 196104
rect 270731 196064 270776 196092
rect 270770 196052 270776 196064
rect 270828 196052 270834 196104
rect 281902 196092 281908 196104
rect 281828 196064 281908 196092
rect 243188 195968 243216 196052
rect 261110 196024 261116 196036
rect 261036 195996 261116 196024
rect 261036 195968 261064 195996
rect 261110 195984 261116 195996
rect 261168 195984 261174 196036
rect 281828 195968 281856 196064
rect 281902 196052 281908 196064
rect 281960 196052 281966 196104
rect 324406 196092 324412 196104
rect 324367 196064 324412 196092
rect 324406 196052 324412 196064
rect 324464 196052 324470 196104
rect 364610 196052 364616 196104
rect 364668 196052 364674 196104
rect 370038 196052 370044 196104
rect 370096 196052 370102 196104
rect 408770 196092 408776 196104
rect 408696 196064 408776 196092
rect 309318 196024 309324 196036
rect 309279 195996 309324 196024
rect 309318 195984 309324 195996
rect 309376 195984 309382 196036
rect 330110 196024 330116 196036
rect 330036 195996 330116 196024
rect 330036 195968 330064 195996
rect 330110 195984 330116 195996
rect 330168 195984 330174 196036
rect 358906 195984 358912 196036
rect 358964 196024 358970 196036
rect 359090 196024 359096 196036
rect 358964 195996 359096 196024
rect 358964 195984 358970 195996
rect 359090 195984 359096 195996
rect 359148 195984 359154 196036
rect 364628 195968 364656 196052
rect 370056 195968 370084 196052
rect 397638 196024 397644 196036
rect 397599 195996 397644 196024
rect 397638 195984 397644 195996
rect 397696 195984 397702 196036
rect 408696 195968 408724 196064
rect 408770 196052 408776 196064
rect 408828 196052 408834 196104
rect 451550 196092 451556 196104
rect 451476 196064 451556 196092
rect 451476 195968 451504 196064
rect 451550 196052 451556 196064
rect 451608 196052 451614 196104
rect 230842 195916 230848 195968
rect 230900 195916 230906 195968
rect 243170 195916 243176 195968
rect 243228 195916 243234 195968
rect 261018 195916 261024 195968
rect 261076 195916 261082 195968
rect 277486 195916 277492 195968
rect 277544 195956 277550 195968
rect 277670 195956 277676 195968
rect 277544 195928 277676 195956
rect 277544 195916 277550 195928
rect 277670 195916 277676 195928
rect 277728 195916 277734 195968
rect 281810 195916 281816 195968
rect 281868 195916 281874 195968
rect 318886 195916 318892 195968
rect 318944 195956 318950 195968
rect 319070 195956 319076 195968
rect 318944 195928 319076 195956
rect 318944 195916 318950 195928
rect 319070 195916 319076 195928
rect 319128 195916 319134 195968
rect 330018 195916 330024 195968
rect 330076 195916 330082 195968
rect 364610 195916 364616 195968
rect 364668 195916 364674 195968
rect 370038 195916 370044 195968
rect 370096 195916 370102 195968
rect 371418 195916 371424 195968
rect 371476 195916 371482 195968
rect 382458 195916 382464 195968
rect 382516 195916 382522 195968
rect 408678 195916 408684 195968
rect 408736 195916 408742 195968
rect 451458 195916 451464 195968
rect 451516 195916 451522 195968
rect 371436 195832 371464 195916
rect 382476 195832 382504 195916
rect 371418 195780 371424 195832
rect 371476 195780 371482 195832
rect 382458 195780 382464 195832
rect 382516 195780 382522 195832
rect 392026 195236 392032 195288
rect 392084 195276 392090 195288
rect 392302 195276 392308 195288
rect 392084 195248 392308 195276
rect 392084 195236 392090 195248
rect 392302 195236 392308 195248
rect 392360 195236 392366 195288
rect 3142 194284 3148 194336
rect 3200 194324 3206 194336
rect 6178 194324 6184 194336
rect 3200 194296 6184 194324
rect 3200 194284 3206 194296
rect 6178 194284 6184 194296
rect 6236 194284 6242 194336
rect 334342 193332 334348 193384
rect 334400 193372 334406 193384
rect 334400 193344 334480 193372
rect 334400 193332 334406 193344
rect 265158 193264 265164 193316
rect 265216 193304 265222 193316
rect 265342 193304 265348 193316
rect 265216 193276 265348 193304
rect 265216 193264 265222 193276
rect 265342 193264 265348 193276
rect 265400 193264 265406 193316
rect 327350 193264 327356 193316
rect 327408 193264 327414 193316
rect 331214 193264 331220 193316
rect 331272 193264 331278 193316
rect 252554 193196 252560 193248
rect 252612 193236 252618 193248
rect 252738 193236 252744 193248
rect 252612 193208 252744 193236
rect 252612 193196 252618 193208
rect 252738 193196 252744 193208
rect 252796 193196 252802 193248
rect 254118 193196 254124 193248
rect 254176 193236 254182 193248
rect 254302 193236 254308 193248
rect 254176 193208 254308 193236
rect 254176 193196 254182 193208
rect 254302 193196 254308 193208
rect 254360 193196 254366 193248
rect 259730 193236 259736 193248
rect 259656 193208 259736 193236
rect 259656 193180 259684 193208
rect 259730 193196 259736 193208
rect 259788 193196 259794 193248
rect 266354 193196 266360 193248
rect 266412 193236 266418 193248
rect 266538 193236 266544 193248
rect 266412 193208 266544 193236
rect 266412 193196 266418 193208
rect 266538 193196 266544 193208
rect 266596 193196 266602 193248
rect 266998 193196 267004 193248
rect 267056 193236 267062 193248
rect 267090 193236 267096 193248
rect 267056 193208 267096 193236
rect 267056 193196 267062 193208
rect 267090 193196 267096 193208
rect 267148 193196 267154 193248
rect 294138 193196 294144 193248
rect 294196 193196 294202 193248
rect 298281 193239 298339 193245
rect 298281 193205 298293 193239
rect 298327 193236 298339 193239
rect 298370 193236 298376 193248
rect 298327 193208 298376 193236
rect 298327 193205 298339 193208
rect 298281 193199 298339 193205
rect 298370 193196 298376 193208
rect 298428 193196 298434 193248
rect 305178 193196 305184 193248
rect 305236 193236 305242 193248
rect 305362 193236 305368 193248
rect 305236 193208 305368 193236
rect 305236 193196 305242 193208
rect 305362 193196 305368 193208
rect 305420 193196 305426 193248
rect 309321 193239 309379 193245
rect 309321 193205 309333 193239
rect 309367 193236 309379 193239
rect 309410 193236 309416 193248
rect 309367 193208 309416 193236
rect 309367 193205 309379 193208
rect 309321 193199 309379 193205
rect 309410 193196 309416 193208
rect 309468 193196 309474 193248
rect 310698 193196 310704 193248
rect 310756 193236 310762 193248
rect 310882 193236 310888 193248
rect 310756 193208 310888 193236
rect 310756 193196 310762 193208
rect 310882 193196 310888 193208
rect 310940 193196 310946 193248
rect 259638 193128 259644 193180
rect 259696 193128 259702 193180
rect 270770 193168 270776 193180
rect 270731 193140 270776 193168
rect 270770 193128 270776 193140
rect 270828 193128 270834 193180
rect 294156 193168 294184 193196
rect 327368 193180 327396 193264
rect 331232 193180 331260 193264
rect 334452 193248 334480 193344
rect 356514 193304 356520 193316
rect 356440 193276 356520 193304
rect 356440 193248 356468 193276
rect 356514 193264 356520 193276
rect 356572 193264 356578 193316
rect 386598 193264 386604 193316
rect 386656 193304 386662 193316
rect 386782 193304 386788 193316
rect 386656 193276 386788 193304
rect 386656 193264 386662 193276
rect 386782 193264 386788 193276
rect 386840 193264 386846 193316
rect 334434 193196 334440 193248
rect 334492 193196 334498 193248
rect 346578 193196 346584 193248
rect 346636 193236 346642 193248
rect 346762 193236 346768 193248
rect 346636 193208 346768 193236
rect 346636 193196 346642 193208
rect 346762 193196 346768 193208
rect 346820 193196 346826 193248
rect 347958 193196 347964 193248
rect 348016 193236 348022 193248
rect 348142 193236 348148 193248
rect 348016 193208 348148 193236
rect 348016 193196 348022 193208
rect 348142 193196 348148 193208
rect 348200 193196 348206 193248
rect 353478 193196 353484 193248
rect 353536 193236 353542 193248
rect 353662 193236 353668 193248
rect 353536 193208 353668 193236
rect 353536 193196 353542 193208
rect 353662 193196 353668 193208
rect 353720 193196 353726 193248
rect 356422 193196 356428 193248
rect 356480 193196 356486 193248
rect 376754 193196 376760 193248
rect 376812 193236 376818 193248
rect 376938 193236 376944 193248
rect 376812 193208 376944 193236
rect 376812 193196 376818 193208
rect 376938 193196 376944 193208
rect 376996 193196 377002 193248
rect 393130 193196 393136 193248
rect 393188 193236 393194 193248
rect 393222 193236 393228 193248
rect 393188 193208 393228 193236
rect 393188 193196 393194 193208
rect 393222 193196 393228 193208
rect 393280 193196 393286 193248
rect 397546 193196 397552 193248
rect 397604 193236 397610 193248
rect 397641 193239 397699 193245
rect 397641 193236 397653 193239
rect 397604 193208 397653 193236
rect 397604 193196 397610 193208
rect 397641 193205 397653 193208
rect 397687 193205 397699 193239
rect 397641 193199 397699 193205
rect 400306 193196 400312 193248
rect 400364 193236 400370 193248
rect 400582 193236 400588 193248
rect 400364 193208 400588 193236
rect 400364 193196 400370 193208
rect 400582 193196 400588 193208
rect 400640 193196 400646 193248
rect 416958 193196 416964 193248
rect 417016 193236 417022 193248
rect 417142 193236 417148 193248
rect 417016 193208 417148 193236
rect 417016 193196 417022 193208
rect 417142 193196 417148 193208
rect 417200 193196 417206 193248
rect 433426 193196 433432 193248
rect 433484 193236 433490 193248
rect 433702 193236 433708 193248
rect 433484 193208 433708 193236
rect 433484 193196 433490 193208
rect 433702 193196 433708 193208
rect 433760 193196 433766 193248
rect 472158 193196 472164 193248
rect 472216 193236 472222 193248
rect 472342 193236 472348 193248
rect 472216 193208 472348 193236
rect 472216 193196 472222 193208
rect 472342 193196 472348 193208
rect 472400 193196 472406 193248
rect 294230 193168 294236 193180
rect 294156 193140 294236 193168
rect 294230 193128 294236 193140
rect 294288 193128 294294 193180
rect 327350 193128 327356 193180
rect 327408 193128 327414 193180
rect 331214 193128 331220 193180
rect 331272 193128 331278 193180
rect 298278 191876 298284 191888
rect 298239 191848 298284 191876
rect 298278 191836 298284 191848
rect 298336 191836 298342 191888
rect 324406 191876 324412 191888
rect 324367 191848 324412 191876
rect 324406 191836 324412 191848
rect 324464 191836 324470 191888
rect 266449 191811 266507 191817
rect 266449 191777 266461 191811
rect 266495 191808 266507 191811
rect 266538 191808 266544 191820
rect 266495 191780 266544 191808
rect 266495 191777 266507 191780
rect 266449 191771 266507 191777
rect 266538 191768 266544 191780
rect 266596 191768 266602 191820
rect 270402 191768 270408 191820
rect 270460 191808 270466 191820
rect 270770 191808 270776 191820
rect 270460 191780 270776 191808
rect 270460 191768 270466 191780
rect 270770 191768 270776 191780
rect 270828 191768 270834 191820
rect 369762 191768 369768 191820
rect 369820 191808 369826 191820
rect 370038 191808 370044 191820
rect 369820 191780 370044 191808
rect 369820 191768 369826 191780
rect 370038 191768 370044 191780
rect 370096 191768 370102 191820
rect 375466 191768 375472 191820
rect 375524 191808 375530 191820
rect 375558 191808 375564 191820
rect 375524 191780 375564 191808
rect 375524 191768 375530 191780
rect 375558 191768 375564 191780
rect 375616 191768 375622 191820
rect 324222 191700 324228 191752
rect 324280 191740 324286 191752
rect 324406 191740 324412 191752
rect 324280 191712 324412 191740
rect 324280 191700 324286 191712
rect 324406 191700 324412 191712
rect 324464 191700 324470 191752
rect 236273 189091 236331 189097
rect 236273 189057 236285 189091
rect 236319 189088 236331 189091
rect 236362 189088 236368 189100
rect 236319 189060 236368 189088
rect 236319 189057 236331 189060
rect 236273 189051 236331 189057
rect 236362 189048 236368 189060
rect 236420 189048 236426 189100
rect 295610 188476 295616 188488
rect 295571 188448 295616 188476
rect 295610 188436 295616 188448
rect 295668 188436 295674 188488
rect 327166 188096 327172 188148
rect 327224 188136 327230 188148
rect 327350 188136 327356 188148
rect 327224 188108 327356 188136
rect 327224 188096 327230 188108
rect 327350 188096 327356 188108
rect 327408 188096 327414 188148
rect 244458 186940 244464 186992
rect 244516 186980 244522 186992
rect 244642 186980 244648 186992
rect 244516 186952 244648 186980
rect 244516 186940 244522 186952
rect 244642 186940 244648 186952
rect 244700 186940 244706 186992
rect 298278 186464 298284 186516
rect 298336 186504 298342 186516
rect 298373 186507 298431 186513
rect 298373 186504 298385 186507
rect 298336 186476 298385 186504
rect 298336 186464 298342 186476
rect 298373 186473 298385 186476
rect 298419 186473 298431 186507
rect 298373 186467 298431 186473
rect 267090 186436 267096 186448
rect 267016 186408 267096 186436
rect 233326 186328 233332 186380
rect 233384 186368 233390 186380
rect 233510 186368 233516 186380
rect 233384 186340 233516 186368
rect 233384 186328 233390 186340
rect 233510 186328 233516 186340
rect 233568 186328 233574 186380
rect 267016 186312 267044 186408
rect 267090 186396 267096 186408
rect 267148 186396 267154 186448
rect 334434 186436 334440 186448
rect 334395 186408 334440 186436
rect 334434 186396 334440 186408
rect 334492 186396 334498 186448
rect 352098 186436 352104 186448
rect 352024 186408 352104 186436
rect 321738 186368 321744 186380
rect 321664 186340 321744 186368
rect 321664 186312 321692 186340
rect 321738 186328 321744 186340
rect 321796 186328 321802 186380
rect 352024 186312 352052 186408
rect 352098 186396 352104 186408
rect 352156 186396 352162 186448
rect 357529 186439 357587 186445
rect 357529 186405 357541 186439
rect 357575 186436 357587 186439
rect 357618 186436 357624 186448
rect 357575 186408 357624 186436
rect 357575 186405 357587 186408
rect 357529 186399 357587 186405
rect 357618 186396 357624 186408
rect 357676 186396 357682 186448
rect 397730 186328 397736 186380
rect 397788 186328 397794 186380
rect 422294 186328 422300 186380
rect 422352 186368 422358 186380
rect 422478 186368 422484 186380
rect 422352 186340 422484 186368
rect 422352 186328 422358 186340
rect 422478 186328 422484 186340
rect 422536 186328 422542 186380
rect 266998 186260 267004 186312
rect 267056 186260 267062 186312
rect 321646 186260 321652 186312
rect 321704 186260 321710 186312
rect 352006 186260 352012 186312
rect 352064 186260 352070 186312
rect 397748 186244 397776 186328
rect 451458 186260 451464 186312
rect 451516 186300 451522 186312
rect 451642 186300 451648 186312
rect 451516 186272 451648 186300
rect 451516 186260 451522 186272
rect 451642 186260 451648 186272
rect 451700 186260 451706 186312
rect 397730 186192 397736 186244
rect 397788 186192 397794 186244
rect 230658 183540 230664 183592
rect 230716 183580 230722 183592
rect 230934 183580 230940 183592
rect 230716 183552 230940 183580
rect 230716 183540 230722 183552
rect 230934 183540 230940 183552
rect 230992 183540 230998 183592
rect 252738 183540 252744 183592
rect 252796 183540 252802 183592
rect 254302 183580 254308 183592
rect 254228 183552 254308 183580
rect 252756 183444 252784 183540
rect 254228 183524 254256 183552
rect 254302 183540 254308 183552
rect 254360 183540 254366 183592
rect 277578 183540 277584 183592
rect 277636 183580 277642 183592
rect 277670 183580 277676 183592
rect 277636 183552 277676 183580
rect 277636 183540 277642 183552
rect 277670 183540 277676 183552
rect 277728 183540 277734 183592
rect 287238 183540 287244 183592
rect 287296 183580 287302 183592
rect 287422 183580 287428 183592
rect 287296 183552 287428 183580
rect 287296 183540 287302 183552
rect 287422 183540 287428 183552
rect 287480 183540 287486 183592
rect 294046 183540 294052 183592
rect 294104 183580 294110 183592
rect 294230 183580 294236 183592
rect 294104 183552 294236 183580
rect 294104 183540 294110 183552
rect 294230 183540 294236 183552
rect 294288 183540 294294 183592
rect 295610 183580 295616 183592
rect 295571 183552 295616 183580
rect 295610 183540 295616 183552
rect 295668 183540 295674 183592
rect 298370 183580 298376 183592
rect 298331 183552 298376 183580
rect 298370 183540 298376 183552
rect 298428 183540 298434 183592
rect 318978 183540 318984 183592
rect 319036 183580 319042 183592
rect 319070 183580 319076 183592
rect 319036 183552 319076 183580
rect 319036 183540 319042 183552
rect 319070 183540 319076 183552
rect 319128 183540 319134 183592
rect 331122 183540 331128 183592
rect 331180 183580 331186 183592
rect 331490 183580 331496 183592
rect 331180 183552 331496 183580
rect 331180 183540 331186 183552
rect 331490 183540 331496 183552
rect 331548 183540 331554 183592
rect 334434 183580 334440 183592
rect 334395 183552 334440 183580
rect 334434 183540 334440 183552
rect 334492 183540 334498 183592
rect 357526 183580 357532 183592
rect 357487 183552 357532 183580
rect 357526 183540 357532 183552
rect 357584 183540 357590 183592
rect 381170 183540 381176 183592
rect 381228 183580 381234 183592
rect 381354 183580 381360 183592
rect 381228 183552 381360 183580
rect 381228 183540 381234 183552
rect 381354 183540 381360 183552
rect 381412 183540 381418 183592
rect 393222 183540 393228 183592
rect 393280 183580 393286 183592
rect 393406 183580 393412 183592
rect 393280 183552 393412 183580
rect 393280 183540 393286 183552
rect 393406 183540 393412 183552
rect 393464 183540 393470 183592
rect 408770 183540 408776 183592
rect 408828 183580 408834 183592
rect 408954 183580 408960 183592
rect 408828 183552 408960 183580
rect 408828 183540 408834 183552
rect 408954 183540 408960 183552
rect 409012 183540 409018 183592
rect 254210 183472 254216 183524
rect 254268 183472 254274 183524
rect 451642 183512 451648 183524
rect 451603 183484 451648 183512
rect 451642 183472 451648 183484
rect 451700 183472 451706 183524
rect 466546 183472 466552 183524
rect 466604 183512 466610 183524
rect 466638 183512 466644 183524
rect 466604 183484 466644 183512
rect 466604 183472 466610 183484
rect 466638 183472 466644 183484
rect 466696 183472 466702 183524
rect 252830 183444 252836 183456
rect 252756 183416 252836 183444
rect 252830 183404 252836 183416
rect 252888 183404 252894 183456
rect 266446 183376 266452 183388
rect 266407 183348 266452 183376
rect 266446 183336 266452 183348
rect 266504 183336 266510 183388
rect 386690 182180 386696 182232
rect 386748 182220 386754 182232
rect 386782 182220 386788 182232
rect 386748 182192 386788 182220
rect 386748 182180 386754 182192
rect 386782 182180 386788 182192
rect 386840 182180 386846 182232
rect 252830 182152 252836 182164
rect 252791 182124 252836 182152
rect 252830 182112 252836 182124
rect 252888 182112 252894 182164
rect 259730 182112 259736 182164
rect 259788 182152 259794 182164
rect 259914 182152 259920 182164
rect 259788 182124 259920 182152
rect 259788 182112 259794 182124
rect 259914 182112 259920 182124
rect 259972 182112 259978 182164
rect 270586 182112 270592 182164
rect 270644 182152 270650 182164
rect 270862 182152 270868 182164
rect 270644 182124 270868 182152
rect 270644 182112 270650 182124
rect 270862 182112 270868 182124
rect 270920 182112 270926 182164
rect 318978 182112 318984 182164
rect 319036 182152 319042 182164
rect 319070 182152 319076 182164
rect 319036 182124 319076 182152
rect 319036 182112 319042 182124
rect 319070 182112 319076 182124
rect 319128 182112 319134 182164
rect 369946 182112 369952 182164
rect 370004 182152 370010 182164
rect 370406 182152 370412 182164
rect 370004 182124 370412 182152
rect 370004 182112 370010 182124
rect 370406 182112 370412 182124
rect 370464 182112 370470 182164
rect 397362 182112 397368 182164
rect 397420 182152 397426 182164
rect 397730 182152 397736 182164
rect 397420 182124 397736 182152
rect 397420 182112 397426 182124
rect 397730 182112 397736 182124
rect 397788 182112 397794 182164
rect 292758 180860 292764 180872
rect 292719 180832 292764 180860
rect 292758 180820 292764 180832
rect 292816 180820 292822 180872
rect 232130 180792 232136 180804
rect 232091 180764 232136 180792
rect 232130 180752 232136 180764
rect 232188 180752 232194 180804
rect 243170 180752 243176 180804
rect 243228 180792 243234 180804
rect 243354 180792 243360 180804
rect 243228 180764 243360 180792
rect 243228 180752 243234 180764
rect 243354 180752 243360 180764
rect 243412 180752 243418 180804
rect 386601 180795 386659 180801
rect 386601 180761 386613 180795
rect 386647 180792 386659 180795
rect 386690 180792 386696 180804
rect 386647 180764 386696 180792
rect 386647 180761 386659 180764
rect 386601 180755 386659 180761
rect 386690 180752 386696 180764
rect 386748 180752 386754 180804
rect 392121 180795 392179 180801
rect 392121 180761 392133 180795
rect 392167 180792 392179 180795
rect 392210 180792 392216 180804
rect 392167 180764 392216 180792
rect 392167 180761 392179 180764
rect 392121 180755 392179 180761
rect 392210 180752 392216 180764
rect 392268 180752 392274 180804
rect 2774 179460 2780 179512
rect 2832 179500 2838 179512
rect 4890 179500 4896 179512
rect 2832 179472 4896 179500
rect 2832 179460 2838 179472
rect 4890 179460 4896 179472
rect 4948 179460 4954 179512
rect 236362 179364 236368 179376
rect 236323 179336 236368 179364
rect 236362 179324 236368 179336
rect 236420 179324 236426 179376
rect 359090 178820 359096 178832
rect 359016 178792 359096 178820
rect 359016 178764 359044 178792
rect 359090 178780 359096 178792
rect 359148 178780 359154 178832
rect 358998 178712 359004 178764
rect 359056 178712 359062 178764
rect 254121 177327 254179 177333
rect 254121 177293 254133 177327
rect 254167 177324 254179 177327
rect 254210 177324 254216 177336
rect 254167 177296 254216 177324
rect 254167 177293 254179 177296
rect 254121 177287 254179 177293
rect 254210 177284 254216 177296
rect 254268 177284 254274 177336
rect 298370 176780 298376 176792
rect 298296 176752 298376 176780
rect 294046 176672 294052 176724
rect 294104 176672 294110 176724
rect 277578 176604 277584 176656
rect 277636 176604 277642 176656
rect 288618 176604 288624 176656
rect 288676 176604 288682 176656
rect 277596 176520 277624 176604
rect 288636 176520 288664 176604
rect 294064 176576 294092 176672
rect 298296 176656 298324 176752
rect 298370 176740 298376 176752
rect 298428 176740 298434 176792
rect 309410 176780 309416 176792
rect 309336 176752 309416 176780
rect 309336 176656 309364 176752
rect 309410 176740 309416 176752
rect 309468 176740 309474 176792
rect 408770 176740 408776 176792
rect 408828 176740 408834 176792
rect 321646 176672 321652 176724
rect 321704 176672 321710 176724
rect 327166 176672 327172 176724
rect 327224 176672 327230 176724
rect 298278 176604 298284 176656
rect 298336 176604 298342 176656
rect 309318 176604 309324 176656
rect 309376 176604 309382 176656
rect 294138 176576 294144 176588
rect 294064 176548 294144 176576
rect 294138 176536 294144 176548
rect 294196 176536 294202 176588
rect 321664 176576 321692 176672
rect 321738 176576 321744 176588
rect 321664 176548 321744 176576
rect 321738 176536 321744 176548
rect 321796 176536 321802 176588
rect 327184 176576 327212 176672
rect 371418 176604 371424 176656
rect 371476 176604 371482 176656
rect 382458 176604 382464 176656
rect 382516 176604 382522 176656
rect 400398 176604 400404 176656
rect 400456 176644 400462 176656
rect 400582 176644 400588 176656
rect 400456 176616 400588 176644
rect 400456 176604 400462 176616
rect 400582 176604 400588 176616
rect 400640 176604 400646 176656
rect 327258 176576 327264 176588
rect 327184 176548 327264 176576
rect 327258 176536 327264 176548
rect 327316 176536 327322 176588
rect 371436 176520 371464 176604
rect 382476 176520 382504 176604
rect 408788 176588 408816 176740
rect 427906 176712 427912 176724
rect 427867 176684 427912 176712
rect 427906 176672 427912 176684
rect 427964 176672 427970 176724
rect 433610 176644 433616 176656
rect 433571 176616 433616 176644
rect 433610 176604 433616 176616
rect 433668 176604 433674 176656
rect 408770 176536 408776 176588
rect 408828 176536 408834 176588
rect 277578 176468 277584 176520
rect 277636 176468 277642 176520
rect 288618 176468 288624 176520
rect 288676 176468 288682 176520
rect 371418 176468 371424 176520
rect 371476 176468 371482 176520
rect 382458 176468 382464 176520
rect 382516 176468 382522 176520
rect 334342 175896 334348 175908
rect 334303 175868 334348 175896
rect 334342 175856 334348 175868
rect 334400 175856 334406 175908
rect 324222 175380 324228 175432
rect 324280 175420 324286 175432
rect 324498 175420 324504 175432
rect 324280 175392 324504 175420
rect 324280 175380 324286 175392
rect 324498 175380 324504 175392
rect 324556 175380 324562 175432
rect 230750 174360 230756 174412
rect 230808 174400 230814 174412
rect 230934 174400 230940 174412
rect 230808 174372 230940 174400
rect 230808 174360 230814 174372
rect 230934 174360 230940 174372
rect 230992 174360 230998 174412
rect 265250 174020 265256 174072
rect 265308 174020 265314 174072
rect 250070 173992 250076 174004
rect 249996 173964 250076 173992
rect 241790 173884 241796 173936
rect 241848 173924 241854 173936
rect 241974 173924 241980 173936
rect 241848 173896 241980 173924
rect 241848 173884 241854 173896
rect 241974 173884 241980 173896
rect 242032 173884 242038 173936
rect 249996 173868 250024 173964
rect 250070 173952 250076 173964
rect 250128 173952 250134 174004
rect 265268 173936 265296 174020
rect 265250 173884 265256 173936
rect 265308 173884 265314 173936
rect 282914 173884 282920 173936
rect 282972 173924 282978 173936
rect 283098 173924 283104 173936
rect 282972 173896 283104 173924
rect 282972 173884 282978 173896
rect 283098 173884 283104 173896
rect 283156 173884 283162 173936
rect 305178 173884 305184 173936
rect 305236 173924 305242 173936
rect 305362 173924 305368 173936
rect 305236 173896 305368 173924
rect 305236 173884 305242 173896
rect 305362 173884 305368 173896
rect 305420 173884 305426 173936
rect 308122 173884 308128 173936
rect 308180 173924 308186 173936
rect 308306 173924 308312 173936
rect 308180 173896 308312 173924
rect 308180 173884 308186 173896
rect 308306 173884 308312 173896
rect 308364 173884 308370 173936
rect 346578 173884 346584 173936
rect 346636 173924 346642 173936
rect 346762 173924 346768 173936
rect 346636 173896 346768 173924
rect 346636 173884 346642 173896
rect 346762 173884 346768 173896
rect 346820 173884 346826 173936
rect 347958 173884 347964 173936
rect 348016 173924 348022 173936
rect 348142 173924 348148 173936
rect 348016 173896 348148 173924
rect 348016 173884 348022 173896
rect 348142 173884 348148 173896
rect 348200 173884 348206 173936
rect 352006 173884 352012 173936
rect 352064 173924 352070 173936
rect 352098 173924 352104 173936
rect 352064 173896 352104 173924
rect 352064 173884 352070 173896
rect 352098 173884 352104 173896
rect 352156 173884 352162 173936
rect 353478 173884 353484 173936
rect 353536 173924 353542 173936
rect 353662 173924 353668 173936
rect 353536 173896 353668 173924
rect 353536 173884 353542 173896
rect 353662 173884 353668 173896
rect 353720 173884 353726 173936
rect 356422 173884 356428 173936
rect 356480 173924 356486 173936
rect 356606 173924 356612 173936
rect 356480 173896 356612 173924
rect 356480 173884 356486 173896
rect 356606 173884 356612 173896
rect 356664 173884 356670 173936
rect 376754 173884 376760 173936
rect 376812 173924 376818 173936
rect 376938 173924 376944 173936
rect 376812 173896 376944 173924
rect 376812 173884 376818 173896
rect 376938 173884 376944 173896
rect 376996 173884 377002 173936
rect 380802 173884 380808 173936
rect 380860 173924 380866 173936
rect 380986 173924 380992 173936
rect 380860 173896 380992 173924
rect 380860 173884 380866 173896
rect 380986 173884 380992 173896
rect 381044 173884 381050 173936
rect 416958 173884 416964 173936
rect 417016 173924 417022 173936
rect 417142 173924 417148 173936
rect 417016 173896 417148 173924
rect 417016 173884 417022 173896
rect 417142 173884 417148 173896
rect 417200 173884 417206 173936
rect 422478 173884 422484 173936
rect 422536 173924 422542 173936
rect 422662 173924 422668 173936
rect 422536 173896 422668 173924
rect 422536 173884 422542 173896
rect 422662 173884 422668 173896
rect 422720 173884 422726 173936
rect 427906 173924 427912 173936
rect 427867 173896 427912 173924
rect 427906 173884 427912 173896
rect 427964 173884 427970 173936
rect 433610 173924 433616 173936
rect 433571 173896 433616 173924
rect 433610 173884 433616 173896
rect 433668 173884 433674 173936
rect 451645 173927 451703 173933
rect 451645 173893 451657 173927
rect 451691 173924 451703 173927
rect 451734 173924 451740 173936
rect 451691 173896 451740 173924
rect 451691 173893 451703 173896
rect 451645 173887 451703 173893
rect 451734 173884 451740 173896
rect 451792 173884 451798 173936
rect 472158 173884 472164 173936
rect 472216 173924 472222 173936
rect 472342 173924 472348 173936
rect 472216 173896 472348 173924
rect 472216 173884 472222 173896
rect 472342 173884 472348 173896
rect 472400 173884 472406 173936
rect 249978 173816 249984 173868
rect 250036 173816 250042 173868
rect 252830 172564 252836 172576
rect 252791 172536 252836 172564
rect 252830 172524 252836 172536
rect 252888 172524 252894 172576
rect 254118 172564 254124 172576
rect 254079 172536 254124 172564
rect 254118 172524 254124 172536
rect 254176 172524 254182 172576
rect 298278 172496 298284 172508
rect 298239 172468 298284 172496
rect 298278 172456 298284 172468
rect 298336 172456 298342 172508
rect 309318 172496 309324 172508
rect 309279 172468 309324 172496
rect 309318 172456 309324 172468
rect 309376 172456 309382 172508
rect 292758 171232 292764 171284
rect 292816 171232 292822 171284
rect 292776 171148 292804 171232
rect 292758 171096 292764 171148
rect 292816 171096 292822 171148
rect 386598 171136 386604 171148
rect 386559 171108 386604 171136
rect 386598 171096 386604 171108
rect 386656 171096 386662 171148
rect 392118 171136 392124 171148
rect 392079 171108 392124 171136
rect 392118 171096 392124 171108
rect 392176 171096 392182 171148
rect 243078 171068 243084 171080
rect 243039 171040 243084 171068
rect 243078 171028 243084 171040
rect 243136 171028 243142 171080
rect 295518 171068 295524 171080
rect 295479 171040 295524 171068
rect 295518 171028 295524 171040
rect 295576 171028 295582 171080
rect 324498 171068 324504 171080
rect 324459 171040 324504 171068
rect 324498 171028 324504 171040
rect 324556 171028 324562 171080
rect 238754 170280 238760 170332
rect 238812 170320 238818 170332
rect 248322 170320 248328 170332
rect 238812 170292 248328 170320
rect 238812 170280 238818 170292
rect 248322 170280 248328 170292
rect 248380 170280 248386 170332
rect 280062 170144 280068 170196
rect 280120 170144 280126 170196
rect 280080 169992 280108 170144
rect 280062 169940 280068 169992
rect 280120 169940 280126 169992
rect 289630 169940 289636 169992
rect 289688 169980 289694 169992
rect 292942 169980 292948 169992
rect 289688 169952 292948 169980
rect 289688 169940 289694 169952
rect 292942 169940 292948 169952
rect 293000 169940 293006 169992
rect 267734 169872 267740 169924
rect 267792 169912 267798 169924
rect 278682 169912 278688 169924
rect 267792 169884 278688 169912
rect 267792 169872 267798 169884
rect 278682 169872 278688 169884
rect 278740 169872 278746 169924
rect 475930 169872 475936 169924
rect 475988 169912 475994 169924
rect 478138 169912 478144 169924
rect 475988 169884 478144 169912
rect 475988 169872 475994 169884
rect 478138 169872 478144 169884
rect 478196 169872 478202 169924
rect 326062 169804 326068 169856
rect 326120 169844 326126 169856
rect 331306 169844 331312 169856
rect 326120 169816 331312 169844
rect 326120 169804 326126 169816
rect 331306 169804 331312 169816
rect 331364 169804 331370 169856
rect 425054 169804 425060 169856
rect 425112 169844 425118 169856
rect 434530 169844 434536 169856
rect 425112 169816 434536 169844
rect 425112 169804 425118 169816
rect 434530 169804 434536 169816
rect 434588 169804 434594 169856
rect 334345 169779 334403 169785
rect 334345 169745 334357 169779
rect 334391 169776 334403 169779
rect 334526 169776 334532 169788
rect 334391 169748 334532 169776
rect 334391 169745 334403 169748
rect 334345 169739 334403 169745
rect 334526 169736 334532 169748
rect 334584 169736 334590 169788
rect 364518 167668 364524 167680
rect 364479 167640 364524 167668
rect 364518 167628 364524 167640
rect 364576 167628 364582 167680
rect 270678 167016 270684 167068
rect 270736 167016 270742 167068
rect 358998 167016 359004 167068
rect 359056 167016 359062 167068
rect 422294 167016 422300 167068
rect 422352 167056 422358 167068
rect 422478 167056 422484 167068
rect 422352 167028 422484 167056
rect 422352 167016 422358 167028
rect 422478 167016 422484 167028
rect 422536 167016 422542 167068
rect 230750 166948 230756 167000
rect 230808 166988 230814 167000
rect 230934 166988 230940 167000
rect 230808 166960 230940 166988
rect 230808 166948 230814 166960
rect 230934 166948 230940 166960
rect 230992 166948 230998 167000
rect 270696 166920 270724 167016
rect 281718 166948 281724 167000
rect 281776 166988 281782 167000
rect 281902 166988 281908 167000
rect 281776 166960 281908 166988
rect 281776 166948 281782 166960
rect 281902 166948 281908 166960
rect 281960 166948 281966 167000
rect 298278 166988 298284 167000
rect 298239 166960 298284 166988
rect 298278 166948 298284 166960
rect 298336 166948 298342 167000
rect 270770 166920 270776 166932
rect 270696 166892 270776 166920
rect 270770 166880 270776 166892
rect 270828 166880 270834 166932
rect 359016 166920 359044 167016
rect 359090 166920 359096 166932
rect 359016 166892 359096 166920
rect 359090 166880 359096 166892
rect 359148 166880 359154 166932
rect 400306 164228 400312 164280
rect 400364 164268 400370 164280
rect 400398 164268 400404 164280
rect 400364 164240 400404 164268
rect 400364 164228 400370 164240
rect 400398 164228 400404 164240
rect 400456 164228 400462 164280
rect 230658 164160 230664 164212
rect 230716 164200 230722 164212
rect 230934 164200 230940 164212
rect 230716 164172 230940 164200
rect 230716 164160 230722 164172
rect 230934 164160 230940 164172
rect 230992 164160 230998 164212
rect 240134 164160 240140 164212
rect 240192 164200 240198 164212
rect 240318 164200 240324 164212
rect 240192 164172 240324 164200
rect 240192 164160 240198 164172
rect 240318 164160 240324 164172
rect 240376 164160 240382 164212
rect 252554 164160 252560 164212
rect 252612 164200 252618 164212
rect 252830 164200 252836 164212
rect 252612 164172 252836 164200
rect 252612 164160 252618 164172
rect 252830 164160 252836 164172
rect 252888 164160 252894 164212
rect 254118 164160 254124 164212
rect 254176 164200 254182 164212
rect 254302 164200 254308 164212
rect 254176 164172 254308 164200
rect 254176 164160 254182 164172
rect 254302 164160 254308 164172
rect 254360 164160 254366 164212
rect 255498 164160 255504 164212
rect 255556 164200 255562 164212
rect 255590 164200 255596 164212
rect 255556 164172 255596 164200
rect 255556 164160 255562 164172
rect 255590 164160 255596 164172
rect 255648 164160 255654 164212
rect 259638 164200 259644 164212
rect 259599 164172 259644 164200
rect 259638 164160 259644 164172
rect 259696 164160 259702 164212
rect 272058 164160 272064 164212
rect 272116 164200 272122 164212
rect 272242 164200 272248 164212
rect 272116 164172 272248 164200
rect 272116 164160 272122 164172
rect 272242 164160 272248 164172
rect 272300 164160 272306 164212
rect 283098 164200 283104 164212
rect 283059 164172 283104 164200
rect 283098 164160 283104 164172
rect 283156 164160 283162 164212
rect 288618 164200 288624 164212
rect 288579 164172 288624 164200
rect 288618 164160 288624 164172
rect 288676 164160 288682 164212
rect 305178 164160 305184 164212
rect 305236 164200 305242 164212
rect 305270 164200 305276 164212
rect 305236 164172 305276 164200
rect 305236 164160 305242 164172
rect 305270 164160 305276 164172
rect 305328 164160 305334 164212
rect 308122 164160 308128 164212
rect 308180 164200 308186 164212
rect 308306 164200 308312 164212
rect 308180 164172 308312 164200
rect 308180 164160 308186 164172
rect 308306 164160 308312 164172
rect 308364 164160 308370 164212
rect 309318 164200 309324 164212
rect 309279 164172 309324 164200
rect 309318 164160 309324 164172
rect 309376 164160 309382 164212
rect 310698 164160 310704 164212
rect 310756 164200 310762 164212
rect 310882 164200 310888 164212
rect 310756 164172 310888 164200
rect 310756 164160 310762 164172
rect 310882 164160 310888 164172
rect 310940 164160 310946 164212
rect 346578 164160 346584 164212
rect 346636 164200 346642 164212
rect 346762 164200 346768 164212
rect 346636 164172 346768 164200
rect 346636 164160 346642 164172
rect 346762 164160 346768 164172
rect 346820 164160 346826 164212
rect 347958 164200 347964 164212
rect 347919 164172 347964 164200
rect 347958 164160 347964 164172
rect 348016 164160 348022 164212
rect 353478 164160 353484 164212
rect 353536 164200 353542 164212
rect 353570 164200 353576 164212
rect 353536 164172 353576 164200
rect 353536 164160 353542 164172
rect 353570 164160 353576 164172
rect 353628 164160 353634 164212
rect 356422 164160 356428 164212
rect 356480 164200 356486 164212
rect 356514 164200 356520 164212
rect 356480 164172 356520 164200
rect 356480 164160 356486 164172
rect 356514 164160 356520 164172
rect 356572 164160 356578 164212
rect 357618 164200 357624 164212
rect 357579 164172 357624 164200
rect 357618 164160 357624 164172
rect 357676 164160 357682 164212
rect 375190 164160 375196 164212
rect 375248 164200 375254 164212
rect 375558 164200 375564 164212
rect 375248 164172 375564 164200
rect 375248 164160 375254 164172
rect 375558 164160 375564 164172
rect 375616 164160 375622 164212
rect 376754 164160 376760 164212
rect 376812 164200 376818 164212
rect 376938 164200 376944 164212
rect 376812 164172 376944 164200
rect 376812 164160 376818 164172
rect 376938 164160 376944 164172
rect 376996 164160 377002 164212
rect 416866 164160 416872 164212
rect 416924 164200 416930 164212
rect 417142 164200 417148 164212
rect 416924 164172 417148 164200
rect 416924 164160 416930 164172
rect 417142 164160 417148 164172
rect 417200 164160 417206 164212
rect 422386 164200 422392 164212
rect 422347 164172 422392 164200
rect 422386 164160 422392 164172
rect 422444 164160 422450 164212
rect 427906 164200 427912 164212
rect 427867 164172 427912 164200
rect 427906 164160 427912 164172
rect 427964 164160 427970 164212
rect 433242 164160 433248 164212
rect 433300 164200 433306 164212
rect 433426 164200 433432 164212
rect 433300 164172 433432 164200
rect 433300 164160 433306 164172
rect 433426 164160 433432 164172
rect 433484 164160 433490 164212
rect 472066 164160 472072 164212
rect 472124 164200 472130 164212
rect 472342 164200 472348 164212
rect 472124 164172 472348 164200
rect 472124 164160 472130 164172
rect 472342 164160 472348 164172
rect 472400 164160 472406 164212
rect 380986 164092 380992 164144
rect 381044 164132 381050 164144
rect 381078 164132 381084 164144
rect 381044 164104 381084 164132
rect 381044 164092 381050 164104
rect 381078 164092 381084 164104
rect 381136 164092 381142 164144
rect 232130 162908 232136 162920
rect 232091 162880 232136 162908
rect 232130 162868 232136 162880
rect 232188 162868 232194 162920
rect 352006 162840 352012 162852
rect 351967 162812 352012 162840
rect 352006 162800 352012 162812
rect 352064 162800 352070 162852
rect 353478 162840 353484 162852
rect 353439 162812 353484 162840
rect 353478 162800 353484 162812
rect 353536 162800 353542 162852
rect 356422 162840 356428 162852
rect 356383 162812 356428 162840
rect 356422 162800 356428 162812
rect 356480 162800 356486 162852
rect 380986 162840 380992 162852
rect 380947 162812 380992 162840
rect 380986 162800 380992 162812
rect 381044 162800 381050 162852
rect 386598 162800 386604 162852
rect 386656 162840 386662 162852
rect 386782 162840 386788 162852
rect 386656 162812 386788 162840
rect 386656 162800 386662 162812
rect 386782 162800 386788 162812
rect 386840 162800 386846 162852
rect 387978 162840 387984 162852
rect 387939 162812 387984 162840
rect 387978 162800 387984 162812
rect 388036 162800 388042 162852
rect 392118 162800 392124 162852
rect 392176 162840 392182 162852
rect 392302 162840 392308 162852
rect 392176 162812 392308 162840
rect 392176 162800 392182 162812
rect 392302 162800 392308 162812
rect 392360 162800 392366 162852
rect 236362 161480 236368 161492
rect 236323 161452 236368 161480
rect 236362 161440 236368 161452
rect 236420 161440 236426 161492
rect 243081 161483 243139 161489
rect 243081 161449 243093 161483
rect 243127 161480 243139 161483
rect 243170 161480 243176 161492
rect 243127 161452 243176 161480
rect 243127 161449 243139 161452
rect 243081 161443 243139 161449
rect 243170 161440 243176 161452
rect 243228 161440 243234 161492
rect 295518 161480 295524 161492
rect 295479 161452 295524 161480
rect 295518 161440 295524 161452
rect 295576 161440 295582 161492
rect 324498 161480 324504 161492
rect 324459 161452 324504 161480
rect 324498 161440 324504 161452
rect 324556 161440 324562 161492
rect 334342 161440 334348 161492
rect 334400 161480 334406 161492
rect 334526 161480 334532 161492
rect 334400 161452 334532 161480
rect 334400 161440 334406 161452
rect 334526 161440 334532 161452
rect 334584 161440 334590 161492
rect 232130 161412 232136 161424
rect 232091 161384 232136 161412
rect 232130 161372 232136 161384
rect 232188 161372 232194 161424
rect 265250 161412 265256 161424
rect 265211 161384 265256 161412
rect 265250 161372 265256 161384
rect 265308 161372 265314 161424
rect 331398 161412 331404 161424
rect 331359 161384 331404 161412
rect 331398 161372 331404 161384
rect 331456 161372 331462 161424
rect 287238 159332 287244 159384
rect 287296 159372 287302 159384
rect 287422 159372 287428 159384
rect 287296 159344 287428 159372
rect 287296 159332 287302 159344
rect 287422 159332 287428 159344
rect 287480 159332 287486 159384
rect 294138 159332 294144 159384
rect 294196 159372 294202 159384
rect 294322 159372 294328 159384
rect 294196 159344 294328 159372
rect 294196 159332 294202 159344
rect 294322 159332 294328 159344
rect 294380 159332 294386 159384
rect 294049 158695 294107 158701
rect 294049 158661 294061 158695
rect 294095 158692 294107 158695
rect 294322 158692 294328 158704
rect 294095 158664 294328 158692
rect 294095 158661 294107 158664
rect 294049 158655 294107 158661
rect 294322 158652 294328 158664
rect 294380 158652 294386 158704
rect 529658 158652 529664 158704
rect 529716 158692 529722 158704
rect 579706 158692 579712 158704
rect 529716 158664 579712 158692
rect 529716 158652 529722 158664
rect 579706 158652 579712 158664
rect 579764 158652 579770 158704
rect 387978 158012 387984 158024
rect 387939 157984 387984 158012
rect 387978 157972 387984 157984
rect 388036 157972 388042 158024
rect 243170 157428 243176 157480
rect 243228 157428 243234 157480
rect 266998 157468 267004 157480
rect 266959 157440 267004 157468
rect 266998 157428 267004 157440
rect 267056 157428 267062 157480
rect 243188 157344 243216 157428
rect 281902 157400 281908 157412
rect 281828 157372 281908 157400
rect 281828 157344 281856 157372
rect 281902 157360 281908 157372
rect 281960 157360 281966 157412
rect 408586 157360 408592 157412
rect 408644 157360 408650 157412
rect 243170 157292 243176 157344
rect 243228 157292 243234 157344
rect 281810 157292 281816 157344
rect 281868 157292 281874 157344
rect 318886 157292 318892 157344
rect 318944 157332 318950 157344
rect 319070 157332 319076 157344
rect 318944 157304 319076 157332
rect 318944 157292 318950 157304
rect 319070 157292 319076 157304
rect 319128 157292 319134 157344
rect 336826 157292 336832 157344
rect 336884 157292 336890 157344
rect 359001 157335 359059 157341
rect 359001 157301 359013 157335
rect 359047 157332 359059 157335
rect 359090 157332 359096 157344
rect 359047 157304 359096 157332
rect 359047 157301 359059 157304
rect 359001 157295 359059 157301
rect 359090 157292 359096 157304
rect 359148 157292 359154 157344
rect 371418 157292 371424 157344
rect 371476 157292 371482 157344
rect 382458 157292 382464 157344
rect 382516 157292 382522 157344
rect 336844 157264 336872 157292
rect 336918 157264 336924 157276
rect 336844 157236 336924 157264
rect 336918 157224 336924 157236
rect 336976 157224 336982 157276
rect 371436 157208 371464 157292
rect 382476 157208 382504 157292
rect 408604 157264 408632 157360
rect 422386 157332 422392 157344
rect 422347 157304 422392 157332
rect 422386 157292 422392 157304
rect 422444 157292 422450 157344
rect 427906 157332 427912 157344
rect 427867 157304 427912 157332
rect 427906 157292 427912 157304
rect 427964 157292 427970 157344
rect 451642 157292 451648 157344
rect 451700 157292 451706 157344
rect 408678 157264 408684 157276
rect 408604 157236 408684 157264
rect 408678 157224 408684 157236
rect 408736 157224 408742 157276
rect 451660 157208 451688 157292
rect 371418 157156 371424 157208
rect 371476 157156 371482 157208
rect 382458 157156 382464 157208
rect 382516 157156 382522 157208
rect 451642 157156 451648 157208
rect 451700 157156 451706 157208
rect 347958 155768 347964 155780
rect 347919 155740 347964 155768
rect 347958 155728 347964 155740
rect 348016 155728 348022 155780
rect 283098 154952 283104 154964
rect 283059 154924 283104 154952
rect 283098 154912 283104 154924
rect 283156 154912 283162 154964
rect 288618 154952 288624 154964
rect 288579 154924 288624 154952
rect 288618 154912 288624 154924
rect 288676 154912 288682 154964
rect 259638 154612 259644 154624
rect 259599 154584 259644 154612
rect 259638 154572 259644 154584
rect 259696 154572 259702 154624
rect 357618 154612 357624 154624
rect 357579 154584 357624 154612
rect 357618 154572 357624 154584
rect 357676 154572 357682 154624
rect 358998 154612 359004 154624
rect 358959 154584 359004 154612
rect 358998 154572 359004 154584
rect 359056 154572 359062 154624
rect 364521 154615 364579 154621
rect 364521 154581 364533 154615
rect 364567 154612 364579 154615
rect 364610 154612 364616 154624
rect 364567 154584 364616 154612
rect 364567 154581 364579 154584
rect 364521 154575 364579 154581
rect 364610 154572 364616 154584
rect 364668 154572 364674 154624
rect 466546 154572 466552 154624
rect 466604 154612 466610 154624
rect 466638 154612 466644 154624
rect 466604 154584 466644 154612
rect 466604 154572 466610 154584
rect 466638 154572 466644 154584
rect 466696 154572 466702 154624
rect 230842 154504 230848 154556
rect 230900 154544 230906 154556
rect 231026 154544 231032 154556
rect 230900 154516 231032 154544
rect 230900 154504 230906 154516
rect 231026 154504 231032 154516
rect 231084 154504 231090 154556
rect 270678 154544 270684 154556
rect 270639 154516 270684 154544
rect 270678 154504 270684 154516
rect 270736 154504 270742 154556
rect 271782 154504 271788 154556
rect 271840 154544 271846 154556
rect 272058 154544 272064 154556
rect 271840 154516 272064 154544
rect 271840 154504 271846 154516
rect 272058 154504 272064 154516
rect 272116 154504 272122 154556
rect 342346 154504 342352 154556
rect 342404 154544 342410 154556
rect 342530 154544 342536 154556
rect 342404 154516 342536 154544
rect 342404 154504 342410 154516
rect 342530 154504 342536 154516
rect 342588 154504 342594 154556
rect 352006 154544 352012 154556
rect 351967 154516 352012 154544
rect 352006 154504 352012 154516
rect 352064 154504 352070 154556
rect 370038 154544 370044 154556
rect 369999 154516 370044 154544
rect 370038 154504 370044 154516
rect 370096 154504 370102 154556
rect 375558 154504 375564 154556
rect 375616 154544 375622 154556
rect 375742 154544 375748 154556
rect 375616 154516 375748 154544
rect 375616 154504 375622 154516
rect 375742 154504 375748 154516
rect 375800 154504 375806 154556
rect 393222 154504 393228 154556
rect 393280 154544 393286 154556
rect 393406 154544 393412 154556
rect 393280 154516 393412 154544
rect 393280 154504 393286 154516
rect 393406 154504 393412 154516
rect 393464 154504 393470 154556
rect 408678 154544 408684 154556
rect 408639 154516 408684 154544
rect 408678 154504 408684 154516
rect 408736 154504 408742 154556
rect 451642 154544 451648 154556
rect 451603 154516 451648 154544
rect 451642 154504 451648 154516
rect 451700 154504 451706 154556
rect 466546 154476 466552 154488
rect 466507 154448 466552 154476
rect 466546 154436 466552 154448
rect 466604 154436 466610 154488
rect 353478 153252 353484 153264
rect 353439 153224 353484 153252
rect 353478 153212 353484 153224
rect 353536 153212 353542 153264
rect 356422 153252 356428 153264
rect 356383 153224 356428 153252
rect 356422 153212 356428 153224
rect 356480 153212 356486 153264
rect 236270 153144 236276 153196
rect 236328 153184 236334 153196
rect 236362 153184 236368 153196
rect 236328 153156 236368 153184
rect 236328 153144 236334 153156
rect 236362 153144 236368 153156
rect 236420 153144 236426 153196
rect 240134 153144 240140 153196
rect 240192 153184 240198 153196
rect 240226 153184 240232 153196
rect 240192 153156 240232 153184
rect 240192 153144 240198 153156
rect 240226 153144 240232 153156
rect 240284 153144 240290 153196
rect 266998 153184 267004 153196
rect 266959 153156 267004 153184
rect 266998 153144 267004 153156
rect 267056 153144 267062 153196
rect 309318 153144 309324 153196
rect 309376 153184 309382 153196
rect 309502 153184 309508 153196
rect 309376 153156 309508 153184
rect 309376 153144 309382 153156
rect 309502 153144 309508 153156
rect 309560 153144 309566 153196
rect 318978 153144 318984 153196
rect 319036 153184 319042 153196
rect 319070 153184 319076 153196
rect 319036 153156 319076 153184
rect 319036 153144 319042 153156
rect 319070 153144 319076 153156
rect 319128 153144 319134 153196
rect 321738 153184 321744 153196
rect 321699 153156 321744 153184
rect 321738 153144 321744 153156
rect 321796 153144 321802 153196
rect 347958 153184 347964 153196
rect 347919 153156 347964 153184
rect 347958 153144 347964 153156
rect 348016 153144 348022 153196
rect 400490 153184 400496 153196
rect 400451 153156 400496 153184
rect 400490 153144 400496 153156
rect 400548 153144 400554 153196
rect 353478 153116 353484 153128
rect 353439 153088 353484 153116
rect 353478 153076 353484 153088
rect 353536 153076 353542 153128
rect 232133 151827 232191 151833
rect 232133 151793 232145 151827
rect 232179 151824 232191 151827
rect 232222 151824 232228 151836
rect 232179 151796 232228 151824
rect 232179 151793 232191 151796
rect 232133 151787 232191 151793
rect 232222 151784 232228 151796
rect 232280 151784 232286 151836
rect 265250 151824 265256 151836
rect 265211 151796 265256 151824
rect 265250 151784 265256 151796
rect 265308 151784 265314 151836
rect 295610 151784 295616 151836
rect 295668 151824 295674 151836
rect 331398 151824 331404 151836
rect 295668 151796 295748 151824
rect 331359 151796 331404 151824
rect 295668 151784 295674 151796
rect 292758 151756 292764 151768
rect 292719 151728 292764 151756
rect 292758 151716 292764 151728
rect 292816 151716 292822 151768
rect 295720 151700 295748 151796
rect 331398 151784 331404 151796
rect 331456 151784 331462 151836
rect 324590 151756 324596 151768
rect 324551 151728 324596 151756
rect 324590 151716 324596 151728
rect 324648 151716 324654 151768
rect 295702 151648 295708 151700
rect 295760 151648 295766 151700
rect 295613 150399 295671 150405
rect 295613 150365 295625 150399
rect 295659 150396 295671 150399
rect 295702 150396 295708 150408
rect 295659 150368 295708 150396
rect 295659 150365 295671 150368
rect 295613 150359 295671 150365
rect 295702 150356 295708 150368
rect 295760 150356 295766 150408
rect 351822 149676 351828 149728
rect 351880 149716 351886 149728
rect 352006 149716 352012 149728
rect 351880 149688 352012 149716
rect 351880 149676 351886 149688
rect 352006 149676 352012 149688
rect 352064 149676 352070 149728
rect 294046 149104 294052 149116
rect 294007 149076 294052 149104
rect 294046 149064 294052 149076
rect 294104 149064 294110 149116
rect 392121 148359 392179 148365
rect 392121 148325 392133 148359
rect 392167 148356 392179 148359
rect 392302 148356 392308 148368
rect 392167 148328 392308 148356
rect 392167 148325 392179 148328
rect 392121 148319 392179 148325
rect 392302 148316 392308 148328
rect 392360 148316 392366 148368
rect 331398 147704 331404 147756
rect 331456 147704 331462 147756
rect 334342 147704 334348 147756
rect 334400 147704 334406 147756
rect 358998 147704 359004 147756
rect 359056 147704 359062 147756
rect 259638 147636 259644 147688
rect 259696 147636 259702 147688
rect 327258 147676 327264 147688
rect 327184 147648 327264 147676
rect 259656 147608 259684 147636
rect 327184 147620 327212 147648
rect 327258 147636 327264 147648
rect 327316 147636 327322 147688
rect 331416 147620 331444 147704
rect 334360 147620 334388 147704
rect 356422 147636 356428 147688
rect 356480 147676 356486 147688
rect 356480 147648 356560 147676
rect 356480 147636 356486 147648
rect 259730 147608 259736 147620
rect 259656 147580 259736 147608
rect 259730 147568 259736 147580
rect 259788 147568 259794 147620
rect 270678 147608 270684 147620
rect 270639 147580 270684 147608
rect 270678 147568 270684 147580
rect 270736 147568 270742 147620
rect 327166 147568 327172 147620
rect 327224 147568 327230 147620
rect 331398 147568 331404 147620
rect 331456 147568 331462 147620
rect 334342 147568 334348 147620
rect 334400 147568 334406 147620
rect 356532 147484 356560 147648
rect 359016 147620 359044 147704
rect 422294 147636 422300 147688
rect 422352 147676 422358 147688
rect 422478 147676 422484 147688
rect 422352 147648 422484 147676
rect 422352 147636 422358 147648
rect 422478 147636 422484 147648
rect 422536 147636 422542 147688
rect 427814 147636 427820 147688
rect 427872 147676 427878 147688
rect 427998 147676 428004 147688
rect 427872 147648 428004 147676
rect 427872 147636 427878 147648
rect 427998 147636 428004 147648
rect 428056 147636 428062 147688
rect 358998 147568 359004 147620
rect 359056 147568 359062 147620
rect 370038 147608 370044 147620
rect 369999 147580 370044 147608
rect 370038 147568 370044 147580
rect 370096 147568 370102 147620
rect 380989 147611 381047 147617
rect 380989 147577 381001 147611
rect 381035 147608 381047 147611
rect 381078 147608 381084 147620
rect 381035 147580 381084 147608
rect 381035 147577 381047 147580
rect 380989 147571 381047 147577
rect 381078 147568 381084 147580
rect 381136 147568 381142 147620
rect 400490 147608 400496 147620
rect 400451 147580 400496 147608
rect 400490 147568 400496 147580
rect 400548 147568 400554 147620
rect 408678 147608 408684 147620
rect 408639 147580 408684 147608
rect 408678 147568 408684 147580
rect 408736 147568 408742 147620
rect 451642 147608 451648 147620
rect 451603 147580 451648 147608
rect 451642 147568 451648 147580
rect 451700 147568 451706 147620
rect 466546 147608 466552 147620
rect 466507 147580 466552 147608
rect 466546 147568 466552 147580
rect 466604 147568 466610 147620
rect 356514 147432 356520 147484
rect 356572 147432 356578 147484
rect 252554 145528 252560 145580
rect 252612 145568 252618 145580
rect 252738 145568 252744 145580
rect 252612 145540 252744 145568
rect 252612 145528 252618 145540
rect 252738 145528 252744 145540
rect 252796 145528 252802 145580
rect 357618 144916 357624 144968
rect 357676 144956 357682 144968
rect 357710 144956 357716 144968
rect 357676 144928 357716 144956
rect 357676 144916 357682 144928
rect 357710 144916 357716 144928
rect 357768 144916 357774 144968
rect 254210 144848 254216 144900
rect 254268 144888 254274 144900
rect 254302 144888 254308 144900
rect 254268 144860 254308 144888
rect 254268 144848 254274 144860
rect 254302 144848 254308 144860
rect 254360 144848 254366 144900
rect 259730 144848 259736 144900
rect 259788 144888 259794 144900
rect 259822 144888 259828 144900
rect 259788 144860 259828 144888
rect 259788 144848 259794 144860
rect 259822 144848 259828 144860
rect 259880 144848 259886 144900
rect 271966 144848 271972 144900
rect 272024 144888 272030 144900
rect 272058 144888 272064 144900
rect 272024 144860 272064 144888
rect 272024 144848 272030 144860
rect 272058 144848 272064 144860
rect 272116 144848 272122 144900
rect 308122 144848 308128 144900
rect 308180 144888 308186 144900
rect 308306 144888 308312 144900
rect 308180 144860 308312 144888
rect 308180 144848 308186 144860
rect 308306 144848 308312 144860
rect 308364 144848 308370 144900
rect 310698 144848 310704 144900
rect 310756 144888 310762 144900
rect 310882 144888 310888 144900
rect 310756 144860 310888 144888
rect 310756 144848 310762 144860
rect 310882 144848 310888 144860
rect 310940 144848 310946 144900
rect 334345 144891 334403 144897
rect 334345 144857 334357 144891
rect 334391 144888 334403 144891
rect 334434 144888 334440 144900
rect 334391 144860 334440 144888
rect 334391 144857 334403 144860
rect 334345 144851 334403 144857
rect 334434 144848 334440 144860
rect 334492 144848 334498 144900
rect 346578 144848 346584 144900
rect 346636 144888 346642 144900
rect 346762 144888 346768 144900
rect 346636 144860 346768 144888
rect 346636 144848 346642 144860
rect 346762 144848 346768 144860
rect 346820 144848 346826 144900
rect 352006 144848 352012 144900
rect 352064 144888 352070 144900
rect 352190 144888 352196 144900
rect 352064 144860 352196 144888
rect 352064 144848 352070 144860
rect 352190 144848 352196 144860
rect 352248 144848 352254 144900
rect 356514 144848 356520 144900
rect 356572 144888 356578 144900
rect 356606 144888 356612 144900
rect 356572 144860 356612 144888
rect 356572 144848 356578 144860
rect 356606 144848 356612 144860
rect 356664 144848 356670 144900
rect 364610 144848 364616 144900
rect 364668 144888 364674 144900
rect 364702 144888 364708 144900
rect 364668 144860 364708 144888
rect 364668 144848 364674 144860
rect 364702 144848 364708 144860
rect 364760 144848 364766 144900
rect 376754 144848 376760 144900
rect 376812 144888 376818 144900
rect 376938 144888 376944 144900
rect 376812 144860 376944 144888
rect 376812 144848 376818 144860
rect 376938 144848 376944 144860
rect 376996 144848 377002 144900
rect 393222 144888 393228 144900
rect 393183 144860 393228 144888
rect 393222 144848 393228 144860
rect 393280 144848 393286 144900
rect 422386 144888 422392 144900
rect 422347 144860 422392 144888
rect 422386 144848 422392 144860
rect 422444 144848 422450 144900
rect 433610 144848 433616 144900
rect 433668 144888 433674 144900
rect 433794 144888 433800 144900
rect 433668 144860 433800 144888
rect 433668 144848 433674 144860
rect 433794 144848 433800 144860
rect 433852 144848 433858 144900
rect 347958 144820 347964 144832
rect 347919 144792 347964 144820
rect 347958 144780 347964 144792
rect 348016 144780 348022 144832
rect 353478 144820 353484 144832
rect 353439 144792 353484 144820
rect 353478 144780 353484 144792
rect 353536 144780 353542 144832
rect 266998 143556 267004 143608
rect 267056 143596 267062 143608
rect 267090 143596 267096 143608
rect 267056 143568 267096 143596
rect 267056 143556 267062 143568
rect 267090 143556 267096 143568
rect 267148 143556 267154 143608
rect 321738 143596 321744 143608
rect 321699 143568 321744 143596
rect 321738 143556 321744 143568
rect 321796 143556 321802 143608
rect 231946 143488 231952 143540
rect 232004 143528 232010 143540
rect 232038 143528 232044 143540
rect 232004 143500 232044 143528
rect 232004 143488 232010 143500
rect 232038 143488 232044 143500
rect 232096 143488 232102 143540
rect 236270 143488 236276 143540
rect 236328 143528 236334 143540
rect 236454 143528 236460 143540
rect 236328 143500 236460 143528
rect 236328 143488 236334 143500
rect 236454 143488 236460 143500
rect 236512 143488 236518 143540
rect 357526 143488 357532 143540
rect 357584 143528 357590 143540
rect 357618 143528 357624 143540
rect 357584 143500 357624 143528
rect 357584 143488 357590 143500
rect 357618 143488 357624 143500
rect 357676 143488 357682 143540
rect 397730 143528 397736 143540
rect 397691 143500 397736 143528
rect 397730 143488 397736 143500
rect 397788 143488 397794 143540
rect 400398 143488 400404 143540
rect 400456 143528 400462 143540
rect 400490 143528 400496 143540
rect 400456 143500 400496 143528
rect 400456 143488 400462 143500
rect 400490 143488 400496 143500
rect 400548 143488 400554 143540
rect 472066 143528 472072 143540
rect 472027 143500 472072 143528
rect 472066 143488 472072 143500
rect 472124 143488 472130 143540
rect 292758 142168 292764 142180
rect 292719 142140 292764 142168
rect 292758 142128 292764 142140
rect 292816 142128 292822 142180
rect 324590 142168 324596 142180
rect 324551 142140 324596 142168
rect 324590 142128 324596 142140
rect 324648 142128 324654 142180
rect 231949 142103 232007 142109
rect 231949 142069 231961 142103
rect 231995 142100 232007 142103
rect 232038 142100 232044 142112
rect 231995 142072 232044 142100
rect 231995 142069 232007 142072
rect 231949 142063 232007 142069
rect 232038 142060 232044 142072
rect 232096 142060 232102 142112
rect 236454 142100 236460 142112
rect 236415 142072 236460 142100
rect 236454 142060 236460 142072
rect 236512 142060 236518 142112
rect 240134 142100 240140 142112
rect 240095 142072 240140 142100
rect 240134 142060 240140 142072
rect 240192 142060 240198 142112
rect 266446 142100 266452 142112
rect 266407 142072 266452 142100
rect 266446 142060 266452 142072
rect 266504 142060 266510 142112
rect 295610 140808 295616 140820
rect 295571 140780 295616 140808
rect 295610 140768 295616 140780
rect 295668 140768 295674 140820
rect 294046 139380 294052 139392
rect 294007 139352 294052 139380
rect 294046 139340 294052 139352
rect 294104 139340 294110 139392
rect 277578 138048 277584 138100
rect 277636 138048 277642 138100
rect 342530 138048 342536 138100
rect 342588 138048 342594 138100
rect 408770 138088 408776 138100
rect 408696 138060 408776 138088
rect 230750 137980 230756 138032
rect 230808 137980 230814 138032
rect 244458 137980 244464 138032
rect 244516 137980 244522 138032
rect 249978 137980 249984 138032
rect 250036 137980 250042 138032
rect 230768 137952 230796 137980
rect 230842 137952 230848 137964
rect 230768 137924 230848 137952
rect 230842 137912 230848 137924
rect 230900 137912 230906 137964
rect 244476 137896 244504 137980
rect 249996 137896 250024 137980
rect 277596 137964 277624 138048
rect 318978 137980 318984 138032
rect 319036 137980 319042 138032
rect 277578 137912 277584 137964
rect 277636 137912 277642 137964
rect 318996 137952 319024 137980
rect 342548 137964 342576 138048
rect 408696 137964 408724 138060
rect 408770 138048 408776 138060
rect 408828 138048 408834 138100
rect 427909 138091 427967 138097
rect 427909 138057 427921 138091
rect 427955 138088 427967 138091
rect 427998 138088 428004 138100
rect 427955 138060 428004 138088
rect 427955 138057 427967 138060
rect 427909 138051 427967 138057
rect 427998 138048 428004 138060
rect 428056 138048 428062 138100
rect 416866 137980 416872 138032
rect 416924 137980 416930 138032
rect 466454 137980 466460 138032
rect 466512 138020 466518 138032
rect 466638 138020 466644 138032
rect 466512 137992 466644 138020
rect 466512 137980 466518 137992
rect 466638 137980 466644 137992
rect 466696 137980 466702 138032
rect 319070 137952 319076 137964
rect 318996 137924 319076 137952
rect 319070 137912 319076 137924
rect 319128 137912 319134 137964
rect 342530 137912 342536 137964
rect 342588 137912 342594 137964
rect 397730 137952 397736 137964
rect 397691 137924 397736 137952
rect 397730 137912 397736 137924
rect 397788 137912 397794 137964
rect 408678 137912 408684 137964
rect 408736 137912 408742 137964
rect 416774 137912 416780 137964
rect 416832 137952 416838 137964
rect 416884 137952 416912 137980
rect 422386 137952 422392 137964
rect 416832 137924 416912 137952
rect 422347 137924 422392 137952
rect 416832 137912 416838 137924
rect 422386 137912 422392 137924
rect 422444 137912 422450 137964
rect 244458 137844 244464 137896
rect 244516 137844 244522 137896
rect 249978 137844 249984 137896
rect 250036 137844 250042 137896
rect 358998 135328 359004 135380
rect 359056 135328 359062 135380
rect 309318 135260 309324 135312
rect 309376 135300 309382 135312
rect 309594 135300 309600 135312
rect 309376 135272 309600 135300
rect 309376 135260 309382 135272
rect 309594 135260 309600 135272
rect 309652 135260 309658 135312
rect 327166 135300 327172 135312
rect 327127 135272 327172 135300
rect 327166 135260 327172 135272
rect 327224 135260 327230 135312
rect 359016 135244 359044 135328
rect 381078 135260 381084 135312
rect 381136 135300 381142 135312
rect 381262 135300 381268 135312
rect 381136 135272 381268 135300
rect 381136 135260 381142 135272
rect 381262 135260 381268 135272
rect 381320 135260 381326 135312
rect 392118 135300 392124 135312
rect 392079 135272 392124 135300
rect 392118 135260 392124 135272
rect 392176 135260 392182 135312
rect 393222 135300 393228 135312
rect 393183 135272 393228 135300
rect 393222 135260 393228 135272
rect 393280 135260 393286 135312
rect 427906 135300 427912 135312
rect 427867 135272 427912 135300
rect 427906 135260 427912 135272
rect 427964 135260 427970 135312
rect 451642 135260 451648 135312
rect 451700 135300 451706 135312
rect 451734 135300 451740 135312
rect 451700 135272 451740 135300
rect 451700 135260 451706 135272
rect 451734 135260 451740 135272
rect 451792 135260 451798 135312
rect 230842 135192 230848 135244
rect 230900 135232 230906 135244
rect 231026 135232 231032 135244
rect 230900 135204 231032 135232
rect 230900 135192 230906 135204
rect 231026 135192 231032 135204
rect 231084 135192 231090 135244
rect 259638 135192 259644 135244
rect 259696 135232 259702 135244
rect 259822 135232 259828 135244
rect 259696 135204 259828 135232
rect 259696 135192 259702 135204
rect 259822 135192 259828 135204
rect 259880 135192 259886 135244
rect 270678 135232 270684 135244
rect 270639 135204 270684 135232
rect 270678 135192 270684 135204
rect 270736 135192 270742 135244
rect 281626 135232 281632 135244
rect 281587 135204 281632 135232
rect 281626 135192 281632 135204
rect 281684 135192 281690 135244
rect 352098 135192 352104 135244
rect 352156 135232 352162 135244
rect 352190 135232 352196 135244
rect 352156 135204 352196 135232
rect 352156 135192 352162 135204
rect 352190 135192 352196 135204
rect 352248 135192 352254 135244
rect 356422 135192 356428 135244
rect 356480 135192 356486 135244
rect 358998 135192 359004 135244
rect 359056 135192 359062 135244
rect 370038 135232 370044 135244
rect 369999 135204 370044 135232
rect 370038 135192 370044 135204
rect 370096 135192 370102 135244
rect 375558 135192 375564 135244
rect 375616 135192 375622 135244
rect 408678 135232 408684 135244
rect 408639 135204 408684 135232
rect 408678 135192 408684 135204
rect 408736 135192 408742 135244
rect 334345 135167 334403 135173
rect 334345 135133 334357 135167
rect 334391 135164 334403 135167
rect 334434 135164 334440 135176
rect 334391 135136 334440 135164
rect 334391 135133 334403 135136
rect 334345 135127 334403 135133
rect 334434 135124 334440 135136
rect 334492 135124 334498 135176
rect 356440 135164 356468 135192
rect 356514 135164 356520 135176
rect 356440 135136 356520 135164
rect 356514 135124 356520 135136
rect 356572 135124 356578 135176
rect 375576 135164 375604 135192
rect 375742 135164 375748 135176
rect 375576 135136 375748 135164
rect 375742 135124 375748 135136
rect 375800 135124 375806 135176
rect 284294 134036 284300 134088
rect 284352 134076 284358 134088
rect 293770 134076 293776 134088
rect 284352 134048 293776 134076
rect 284352 134036 284358 134048
rect 293770 134036 293776 134048
rect 293828 134036 293834 134088
rect 514570 134036 514576 134088
rect 514628 134076 514634 134088
rect 514846 134076 514852 134088
rect 514628 134048 514852 134076
rect 514628 134036 514634 134048
rect 514846 134036 514852 134048
rect 514904 134036 514910 134088
rect 540974 133900 540980 133952
rect 541032 133940 541038 133952
rect 545850 133940 545856 133952
rect 541032 133912 545856 133940
rect 541032 133900 541038 133912
rect 545850 133900 545856 133912
rect 545908 133900 545914 133952
rect 243078 133872 243084 133884
rect 243039 133844 243084 133872
rect 243078 133832 243084 133844
rect 243136 133832 243142 133884
rect 325602 133832 325608 133884
rect 325660 133872 325666 133884
rect 333882 133872 333888 133884
rect 325660 133844 333888 133872
rect 325660 133832 325666 133844
rect 333882 133832 333888 133844
rect 333940 133832 333946 133884
rect 298370 133804 298376 133816
rect 298331 133776 298376 133804
rect 298370 133764 298376 133776
rect 298428 133764 298434 133816
rect 348418 133696 348424 133748
rect 348476 133736 348482 133748
rect 354582 133736 354588 133748
rect 348476 133708 354588 133736
rect 348476 133696 348482 133708
rect 354582 133696 354588 133708
rect 354640 133696 354646 133748
rect 236454 132512 236460 132524
rect 236415 132484 236460 132512
rect 236454 132472 236460 132484
rect 236512 132472 236518 132524
rect 240137 132515 240195 132521
rect 240137 132481 240149 132515
rect 240183 132512 240195 132515
rect 240318 132512 240324 132524
rect 240183 132484 240324 132512
rect 240183 132481 240195 132484
rect 240137 132475 240195 132481
rect 240318 132472 240324 132484
rect 240376 132472 240382 132524
rect 266449 132515 266507 132521
rect 266449 132481 266461 132515
rect 266495 132512 266507 132515
rect 266538 132512 266544 132524
rect 266495 132484 266544 132512
rect 266495 132481 266507 132484
rect 266449 132475 266507 132481
rect 266538 132472 266544 132484
rect 266596 132472 266602 132524
rect 327166 132512 327172 132524
rect 327127 132484 327172 132512
rect 327166 132472 327172 132484
rect 327224 132472 327230 132524
rect 265342 132444 265348 132456
rect 265303 132416 265348 132444
rect 265342 132404 265348 132416
rect 265400 132404 265406 132456
rect 309318 132444 309324 132456
rect 309279 132416 309324 132444
rect 309318 132404 309324 132416
rect 309376 132404 309382 132456
rect 321738 132444 321744 132456
rect 321699 132416 321744 132444
rect 321738 132404 321744 132416
rect 321796 132404 321802 132456
rect 324409 132447 324467 132453
rect 324409 132413 324421 132447
rect 324455 132444 324467 132447
rect 324498 132444 324504 132456
rect 324455 132416 324504 132444
rect 324455 132413 324467 132416
rect 324409 132407 324467 132413
rect 324498 132404 324504 132416
rect 324556 132404 324562 132456
rect 295518 131084 295524 131096
rect 295479 131056 295524 131084
rect 295518 131044 295524 131056
rect 295576 131044 295582 131096
rect 271966 130364 271972 130416
rect 272024 130404 272030 130416
rect 272150 130404 272156 130416
rect 272024 130376 272156 130404
rect 272024 130364 272030 130376
rect 272150 130364 272156 130376
rect 272208 130364 272214 130416
rect 281629 129047 281687 129053
rect 281629 129013 281641 129047
rect 281675 129044 281687 129047
rect 281810 129044 281816 129056
rect 281675 129016 281816 129044
rect 281675 129013 281687 129016
rect 281629 129007 281687 129013
rect 281810 129004 281816 129016
rect 281868 129004 281874 129056
rect 233326 128324 233332 128376
rect 233384 128364 233390 128376
rect 233510 128364 233516 128376
rect 233384 128336 233516 128364
rect 233384 128324 233390 128336
rect 233510 128324 233516 128336
rect 233568 128324 233574 128376
rect 381078 128324 381084 128376
rect 381136 128324 381142 128376
rect 400398 128324 400404 128376
rect 400456 128324 400462 128376
rect 422294 128324 422300 128376
rect 422352 128364 422358 128376
rect 422478 128364 422484 128376
rect 422352 128336 422484 128364
rect 422352 128324 422358 128336
rect 422478 128324 422484 128336
rect 422536 128324 422542 128376
rect 466454 128324 466460 128376
rect 466512 128324 466518 128376
rect 270678 128296 270684 128308
rect 270639 128268 270684 128296
rect 270678 128256 270684 128268
rect 270736 128256 270742 128308
rect 370038 128296 370044 128308
rect 369999 128268 370044 128296
rect 370038 128256 370044 128268
rect 370096 128256 370102 128308
rect 381096 128296 381124 128324
rect 381170 128296 381176 128308
rect 381096 128268 381176 128296
rect 381170 128256 381176 128268
rect 381228 128256 381234 128308
rect 400416 128296 400444 128324
rect 400490 128296 400496 128308
rect 400416 128268 400496 128296
rect 400490 128256 400496 128268
rect 400548 128256 400554 128308
rect 408678 128296 408684 128308
rect 408639 128268 408684 128296
rect 408678 128256 408684 128268
rect 408736 128256 408742 128308
rect 466472 128296 466500 128324
rect 466546 128296 466552 128308
rect 466472 128268 466552 128296
rect 466546 128256 466552 128268
rect 466604 128256 466610 128308
rect 472066 128296 472072 128308
rect 472027 128268 472072 128296
rect 472066 128256 472072 128268
rect 472124 128256 472130 128308
rect 241790 125536 241796 125588
rect 241848 125576 241854 125588
rect 241974 125576 241980 125588
rect 241848 125548 241980 125576
rect 241848 125536 241854 125548
rect 241974 125536 241980 125548
rect 242032 125536 242038 125588
rect 252738 125536 252744 125588
rect 252796 125576 252802 125588
rect 252922 125576 252928 125588
rect 252796 125548 252928 125576
rect 252796 125536 252802 125548
rect 252922 125536 252928 125548
rect 252980 125536 252986 125588
rect 254210 125536 254216 125588
rect 254268 125576 254274 125588
rect 254302 125576 254308 125588
rect 254268 125548 254308 125576
rect 254268 125536 254274 125548
rect 254302 125536 254308 125548
rect 254360 125536 254366 125588
rect 255498 125536 255504 125588
rect 255556 125576 255562 125588
rect 255590 125576 255596 125588
rect 255556 125548 255596 125576
rect 255556 125536 255562 125548
rect 255590 125536 255596 125548
rect 255648 125536 255654 125588
rect 259730 125536 259736 125588
rect 259788 125576 259794 125588
rect 259822 125576 259828 125588
rect 259788 125548 259828 125576
rect 259788 125536 259794 125548
rect 259822 125536 259828 125548
rect 259880 125536 259886 125588
rect 266538 125536 266544 125588
rect 266596 125576 266602 125588
rect 266722 125576 266728 125588
rect 266596 125548 266728 125576
rect 266596 125536 266602 125548
rect 266722 125536 266728 125548
rect 266780 125536 266786 125588
rect 266998 125536 267004 125588
rect 267056 125576 267062 125588
rect 267274 125576 267280 125588
rect 267056 125548 267280 125576
rect 267056 125536 267062 125548
rect 267274 125536 267280 125548
rect 267332 125536 267338 125588
rect 283098 125576 283104 125588
rect 283059 125548 283104 125576
rect 283098 125536 283104 125548
rect 283156 125536 283162 125588
rect 308122 125536 308128 125588
rect 308180 125576 308186 125588
rect 308306 125576 308312 125588
rect 308180 125548 308312 125576
rect 308180 125536 308186 125548
rect 308306 125536 308312 125548
rect 308364 125536 308370 125588
rect 310698 125576 310704 125588
rect 310659 125548 310704 125576
rect 310698 125536 310704 125548
rect 310756 125536 310762 125588
rect 346578 125576 346584 125588
rect 346539 125548 346584 125576
rect 346578 125536 346584 125548
rect 346636 125536 346642 125588
rect 352006 125536 352012 125588
rect 352064 125576 352070 125588
rect 352190 125576 352196 125588
rect 352064 125548 352196 125576
rect 352064 125536 352070 125548
rect 352190 125536 352196 125548
rect 352248 125536 352254 125588
rect 357618 125536 357624 125588
rect 357676 125576 357682 125588
rect 357710 125576 357716 125588
rect 357676 125548 357716 125576
rect 357676 125536 357682 125548
rect 357710 125536 357716 125548
rect 357768 125536 357774 125588
rect 364521 125579 364579 125585
rect 364521 125545 364533 125579
rect 364567 125576 364579 125579
rect 364610 125576 364616 125588
rect 364567 125548 364616 125576
rect 364567 125545 364579 125548
rect 364521 125539 364579 125545
rect 364610 125536 364616 125548
rect 364668 125536 364674 125588
rect 376938 125576 376944 125588
rect 376899 125548 376944 125576
rect 376938 125536 376944 125548
rect 376996 125536 377002 125588
rect 386690 125536 386696 125588
rect 386748 125576 386754 125588
rect 386782 125576 386788 125588
rect 386748 125548 386788 125576
rect 386748 125536 386754 125548
rect 386782 125536 386788 125548
rect 386840 125536 386846 125588
rect 387978 125536 387984 125588
rect 388036 125576 388042 125588
rect 388070 125576 388076 125588
rect 388036 125548 388076 125576
rect 388036 125536 388042 125548
rect 388070 125536 388076 125548
rect 388128 125536 388134 125588
rect 392210 125536 392216 125588
rect 392268 125576 392274 125588
rect 392302 125576 392308 125588
rect 392268 125548 392308 125576
rect 392268 125536 392274 125548
rect 392302 125536 392308 125548
rect 392360 125536 392366 125588
rect 393222 125576 393228 125588
rect 393183 125548 393228 125576
rect 393222 125536 393228 125548
rect 393280 125536 393286 125588
rect 422386 125576 422392 125588
rect 422347 125548 422392 125576
rect 422386 125536 422392 125548
rect 422444 125536 422450 125588
rect 427906 125576 427912 125588
rect 427867 125548 427912 125576
rect 427906 125536 427912 125548
rect 427964 125536 427970 125588
rect 433610 125576 433616 125588
rect 433571 125548 433616 125576
rect 433610 125536 433616 125548
rect 433668 125536 433674 125588
rect 466638 125536 466644 125588
rect 466696 125576 466702 125588
rect 466730 125576 466736 125588
rect 466696 125548 466736 125576
rect 466696 125536 466702 125548
rect 466730 125536 466736 125548
rect 466788 125536 466794 125588
rect 265342 124624 265348 124636
rect 265303 124596 265348 124624
rect 265342 124584 265348 124596
rect 265400 124584 265406 124636
rect 236362 124244 236368 124296
rect 236420 124284 236426 124296
rect 236454 124284 236460 124296
rect 236420 124256 236460 124284
rect 236420 124244 236426 124256
rect 236454 124244 236460 124256
rect 236512 124244 236518 124296
rect 231946 124216 231952 124228
rect 231907 124188 231952 124216
rect 231946 124176 231952 124188
rect 232004 124176 232010 124228
rect 243081 124219 243139 124225
rect 243081 124185 243093 124219
rect 243127 124216 243139 124219
rect 243262 124216 243268 124228
rect 243127 124188 243268 124216
rect 243127 124185 243139 124188
rect 243081 124179 243139 124185
rect 243262 124176 243268 124188
rect 243320 124176 243326 124228
rect 298370 124216 298376 124228
rect 298331 124188 298376 124216
rect 298370 124176 298376 124188
rect 298428 124176 298434 124228
rect 356422 124176 356428 124228
rect 356480 124216 356486 124228
rect 356514 124216 356520 124228
rect 356480 124188 356520 124216
rect 356480 124176 356486 124188
rect 356514 124176 356520 124188
rect 356572 124176 356578 124228
rect 400309 124151 400367 124157
rect 400309 124117 400321 124151
rect 400355 124148 400367 124151
rect 400490 124148 400496 124160
rect 400355 124120 400496 124148
rect 400355 124117 400367 124120
rect 400309 124111 400367 124117
rect 400490 124108 400496 124120
rect 400548 124108 400554 124160
rect 451458 124148 451464 124160
rect 451419 124120 451464 124148
rect 451458 124108 451464 124120
rect 451516 124108 451522 124160
rect 466641 124151 466699 124157
rect 466641 124117 466653 124151
rect 466687 124148 466699 124151
rect 466730 124148 466736 124160
rect 466687 124120 466736 124148
rect 466687 124117 466699 124120
rect 466641 124111 466699 124117
rect 466730 124108 466736 124120
rect 466788 124108 466794 124160
rect 309321 122859 309379 122865
rect 309321 122825 309333 122859
rect 309367 122856 309379 122859
rect 309502 122856 309508 122868
rect 309367 122828 309508 122856
rect 309367 122825 309379 122828
rect 309321 122819 309379 122825
rect 309502 122816 309508 122828
rect 309560 122816 309566 122868
rect 321738 122856 321744 122868
rect 321699 122828 321744 122856
rect 321738 122816 321744 122828
rect 321796 122816 321802 122868
rect 324406 122856 324412 122868
rect 324367 122828 324412 122856
rect 324406 122816 324412 122828
rect 324464 122816 324470 122868
rect 236362 122788 236368 122800
rect 236323 122760 236368 122788
rect 236362 122748 236368 122760
rect 236420 122748 236426 122800
rect 294049 121499 294107 121505
rect 294049 121465 294061 121499
rect 294095 121496 294107 121499
rect 294138 121496 294144 121508
rect 294095 121468 294144 121496
rect 294095 121465 294107 121468
rect 294049 121459 294107 121465
rect 294138 121456 294144 121468
rect 294196 121456 294202 121508
rect 295521 121499 295579 121505
rect 295521 121465 295533 121499
rect 295567 121496 295579 121499
rect 295610 121496 295616 121508
rect 295567 121468 295616 121496
rect 295567 121465 295579 121468
rect 295521 121459 295579 121465
rect 295610 121456 295616 121468
rect 295668 121456 295674 121508
rect 294138 121360 294144 121372
rect 294099 121332 294144 121360
rect 294138 121320 294144 121332
rect 294196 121320 294202 121372
rect 270770 120708 270776 120760
rect 270828 120708 270834 120760
rect 305181 120751 305239 120757
rect 305181 120717 305193 120751
rect 305227 120748 305239 120751
rect 305270 120748 305276 120760
rect 305227 120720 305276 120748
rect 305227 120717 305239 120720
rect 305181 120711 305239 120717
rect 305270 120708 305276 120720
rect 305328 120708 305334 120760
rect 370130 120708 370136 120760
rect 370188 120708 370194 120760
rect 375466 120708 375472 120760
rect 375524 120748 375530 120760
rect 375742 120748 375748 120760
rect 375524 120720 375748 120748
rect 375524 120708 375530 120720
rect 375742 120708 375748 120720
rect 375800 120708 375806 120760
rect 270788 120624 270816 120708
rect 370148 120624 370176 120708
rect 270770 120572 270776 120624
rect 270828 120572 270834 120624
rect 370130 120572 370136 120624
rect 370188 120572 370194 120624
rect 298370 119388 298376 119400
rect 298331 119360 298376 119388
rect 298370 119348 298376 119360
rect 298428 119348 298434 119400
rect 261018 118736 261024 118788
rect 261076 118736 261082 118788
rect 295610 118736 295616 118788
rect 295668 118736 295674 118788
rect 318978 118776 318984 118788
rect 318939 118748 318984 118776
rect 318978 118736 318984 118748
rect 319036 118736 319042 118788
rect 321738 118736 321744 118788
rect 321796 118736 321802 118788
rect 336918 118776 336924 118788
rect 336844 118748 336924 118776
rect 230750 118668 230756 118720
rect 230808 118668 230814 118720
rect 230768 118640 230796 118668
rect 261036 118652 261064 118736
rect 295628 118652 295656 118736
rect 321756 118652 321784 118736
rect 336844 118720 336872 118748
rect 336918 118736 336924 118748
rect 336976 118736 336982 118788
rect 408770 118776 408776 118788
rect 408696 118748 408776 118776
rect 336826 118668 336832 118720
rect 336884 118668 336890 118720
rect 408696 118652 408724 118748
rect 408770 118736 408776 118748
rect 408828 118736 408834 118788
rect 416866 118668 416872 118720
rect 416924 118668 416930 118720
rect 472066 118668 472072 118720
rect 472124 118668 472130 118720
rect 230842 118640 230848 118652
rect 230768 118612 230848 118640
rect 230842 118600 230848 118612
rect 230900 118600 230906 118652
rect 261018 118600 261024 118652
rect 261076 118600 261082 118652
rect 295610 118600 295616 118652
rect 295668 118600 295674 118652
rect 321738 118600 321744 118652
rect 321796 118600 321802 118652
rect 387978 118600 387984 118652
rect 388036 118640 388042 118652
rect 388070 118640 388076 118652
rect 388036 118612 388076 118640
rect 388036 118600 388042 118612
rect 388070 118600 388076 118612
rect 388128 118600 388134 118652
rect 408678 118600 408684 118652
rect 408736 118600 408742 118652
rect 416774 118600 416780 118652
rect 416832 118640 416838 118652
rect 416884 118640 416912 118668
rect 422386 118640 422392 118652
rect 416832 118612 416912 118640
rect 422347 118612 422392 118640
rect 416832 118600 416838 118612
rect 422386 118600 422392 118612
rect 422444 118600 422450 118652
rect 427906 118640 427912 118652
rect 427867 118612 427912 118640
rect 427906 118600 427912 118612
rect 427964 118600 427970 118652
rect 433610 118640 433616 118652
rect 433571 118612 433616 118640
rect 433610 118600 433616 118612
rect 433668 118600 433674 118652
rect 471974 118600 471980 118652
rect 472032 118640 472038 118652
rect 472084 118640 472112 118668
rect 472032 118612 472112 118640
rect 472032 118600 472038 118612
rect 324222 117988 324228 118040
rect 324280 118028 324286 118040
rect 324406 118028 324412 118040
rect 324280 118000 324412 118028
rect 324280 117988 324286 118000
rect 324406 117988 324412 118000
rect 324464 117988 324470 118040
rect 294138 116600 294144 116612
rect 294099 116572 294144 116600
rect 294138 116560 294144 116572
rect 294196 116560 294202 116612
rect 272058 115948 272064 116000
rect 272116 115988 272122 116000
rect 272150 115988 272156 116000
rect 272116 115960 272156 115988
rect 272116 115948 272122 115960
rect 272150 115948 272156 115960
rect 272208 115948 272214 116000
rect 283098 115988 283104 116000
rect 283059 115960 283104 115988
rect 283098 115948 283104 115960
rect 283156 115948 283162 116000
rect 305178 115988 305184 116000
rect 305139 115960 305184 115988
rect 305178 115948 305184 115960
rect 305236 115948 305242 116000
rect 310698 115988 310704 116000
rect 310659 115960 310704 115988
rect 310698 115948 310704 115960
rect 310756 115948 310762 116000
rect 346578 115988 346584 116000
rect 346539 115960 346584 115988
rect 346578 115948 346584 115960
rect 346636 115948 346642 116000
rect 353570 115988 353576 116000
rect 353531 115960 353576 115988
rect 353570 115948 353576 115960
rect 353628 115948 353634 116000
rect 364518 115988 364524 116000
rect 364479 115960 364524 115988
rect 364518 115948 364524 115960
rect 364576 115948 364582 116000
rect 376938 115988 376944 116000
rect 376899 115960 376944 115988
rect 376938 115948 376944 115960
rect 376996 115948 377002 116000
rect 393222 115988 393228 116000
rect 393183 115960 393228 115988
rect 393222 115948 393228 115960
rect 393280 115948 393286 116000
rect 230842 115880 230848 115932
rect 230900 115920 230906 115932
rect 231026 115920 231032 115932
rect 230900 115892 231032 115920
rect 230900 115880 230906 115892
rect 231026 115880 231032 115892
rect 231084 115880 231090 115932
rect 254118 115920 254124 115932
rect 254079 115892 254124 115920
rect 254118 115880 254124 115892
rect 254176 115880 254182 115932
rect 259638 115880 259644 115932
rect 259696 115920 259702 115932
rect 259822 115920 259828 115932
rect 259696 115892 259828 115920
rect 259696 115880 259702 115892
rect 259822 115880 259828 115892
rect 259880 115880 259886 115932
rect 265158 115880 265164 115932
rect 265216 115920 265222 115932
rect 265250 115920 265256 115932
rect 265216 115892 265256 115920
rect 265216 115880 265222 115892
rect 265250 115880 265256 115892
rect 265308 115880 265314 115932
rect 342438 115920 342444 115932
rect 342399 115892 342444 115920
rect 342438 115880 342444 115892
rect 342496 115880 342502 115932
rect 347958 115880 347964 115932
rect 348016 115920 348022 115932
rect 348050 115920 348056 115932
rect 348016 115892 348056 115920
rect 348016 115880 348022 115892
rect 348050 115880 348056 115892
rect 348108 115880 348114 115932
rect 356422 115880 356428 115932
rect 356480 115920 356486 115932
rect 356606 115920 356612 115932
rect 356480 115892 356612 115920
rect 356480 115880 356486 115892
rect 356606 115880 356612 115892
rect 356664 115880 356670 115932
rect 375466 115880 375472 115932
rect 375524 115920 375530 115932
rect 375742 115920 375748 115932
rect 375524 115892 375748 115920
rect 375524 115880 375530 115892
rect 375742 115880 375748 115892
rect 375800 115880 375806 115932
rect 381078 115880 381084 115932
rect 381136 115920 381142 115932
rect 381262 115920 381268 115932
rect 381136 115892 381268 115920
rect 381136 115880 381142 115892
rect 381262 115880 381268 115892
rect 381320 115880 381326 115932
rect 386598 115880 386604 115932
rect 386656 115920 386662 115932
rect 386782 115920 386788 115932
rect 386656 115892 386788 115920
rect 386656 115880 386662 115892
rect 386782 115880 386788 115892
rect 386840 115880 386846 115932
rect 392118 115880 392124 115932
rect 392176 115920 392182 115932
rect 392302 115920 392308 115932
rect 392176 115892 392308 115920
rect 392176 115880 392182 115892
rect 392302 115880 392308 115892
rect 392360 115880 392366 115932
rect 393222 115812 393228 115864
rect 393280 115852 393286 115864
rect 393314 115852 393320 115864
rect 393280 115824 393320 115852
rect 393280 115812 393286 115824
rect 393314 115812 393320 115824
rect 393372 115812 393378 115864
rect 298186 114520 298192 114572
rect 298244 114560 298250 114572
rect 298373 114563 298431 114569
rect 298373 114560 298385 114563
rect 298244 114532 298385 114560
rect 298244 114520 298250 114532
rect 298373 114529 298385 114532
rect 298419 114529 298431 114563
rect 298373 114523 298431 114529
rect 334345 114563 334403 114569
rect 334345 114529 334357 114563
rect 334391 114560 334403 114563
rect 334434 114560 334440 114572
rect 334391 114532 334440 114560
rect 334391 114529 334403 114532
rect 334345 114523 334403 114529
rect 334434 114520 334440 114532
rect 334492 114520 334498 114572
rect 353570 114560 353576 114572
rect 353531 114532 353576 114560
rect 353570 114520 353576 114532
rect 353628 114520 353634 114572
rect 400306 114560 400312 114572
rect 400267 114532 400312 114560
rect 400306 114520 400312 114532
rect 400364 114520 400370 114572
rect 451461 114563 451519 114569
rect 451461 114529 451473 114563
rect 451507 114560 451519 114563
rect 451550 114560 451556 114572
rect 451507 114532 451556 114560
rect 451507 114529 451519 114532
rect 451461 114523 451519 114529
rect 451550 114520 451556 114532
rect 451608 114520 451614 114572
rect 466638 114560 466644 114572
rect 466599 114532 466644 114560
rect 466638 114520 466644 114532
rect 466696 114520 466702 114572
rect 267001 114495 267059 114501
rect 267001 114461 267013 114495
rect 267047 114492 267059 114495
rect 267090 114492 267096 114504
rect 267047 114464 267096 114492
rect 267047 114461 267059 114464
rect 267001 114455 267059 114461
rect 267090 114452 267096 114464
rect 267148 114452 267154 114504
rect 327166 114492 327172 114504
rect 327127 114464 327172 114492
rect 327166 114452 327172 114464
rect 327224 114452 327230 114504
rect 356425 114495 356483 114501
rect 356425 114461 356437 114495
rect 356471 114492 356483 114495
rect 356606 114492 356612 114504
rect 356471 114464 356612 114492
rect 356471 114461 356483 114464
rect 356425 114455 356483 114461
rect 356606 114452 356612 114464
rect 356664 114452 356670 114504
rect 387978 114492 387984 114504
rect 387939 114464 387984 114492
rect 387978 114452 387984 114464
rect 388036 114452 388042 114504
rect 298186 114424 298192 114436
rect 298147 114396 298192 114424
rect 298186 114384 298192 114396
rect 298244 114384 298250 114436
rect 236365 113203 236423 113209
rect 236365 113169 236377 113203
rect 236411 113200 236423 113203
rect 236454 113200 236460 113212
rect 236411 113172 236460 113200
rect 236411 113169 236423 113172
rect 236365 113163 236423 113169
rect 236454 113160 236460 113172
rect 236512 113160 236518 113212
rect 309318 113160 309324 113212
rect 309376 113200 309382 113212
rect 309502 113200 309508 113212
rect 309376 113172 309508 113200
rect 309376 113160 309382 113172
rect 309502 113160 309508 113172
rect 309560 113160 309566 113212
rect 334342 113200 334348 113212
rect 334303 113172 334348 113200
rect 334342 113160 334348 113172
rect 334400 113160 334406 113212
rect 292758 113132 292764 113144
rect 292719 113104 292764 113132
rect 292758 113092 292764 113104
rect 292816 113092 292822 113144
rect 295610 111772 295616 111784
rect 295571 111744 295616 111772
rect 295610 111732 295616 111744
rect 295668 111732 295674 111784
rect 529566 111732 529572 111784
rect 529624 111772 529630 111784
rect 580166 111772 580172 111784
rect 529624 111744 580172 111772
rect 529624 111732 529630 111744
rect 580166 111732 580172 111744
rect 580224 111732 580230 111784
rect 397638 109080 397644 109132
rect 397696 109080 397702 109132
rect 233326 109012 233332 109064
rect 233384 109052 233390 109064
rect 233510 109052 233516 109064
rect 233384 109024 233516 109052
rect 233384 109012 233390 109024
rect 233510 109012 233516 109024
rect 233568 109012 233574 109064
rect 243078 109012 243084 109064
rect 243136 109012 243142 109064
rect 370130 109052 370136 109064
rect 370091 109024 370136 109052
rect 370130 109012 370136 109024
rect 370188 109012 370194 109064
rect 243096 108984 243124 109012
rect 397656 108996 397684 109080
rect 408678 109012 408684 109064
rect 408736 109012 408742 109064
rect 422294 109012 422300 109064
rect 422352 109052 422358 109064
rect 422478 109052 422484 109064
rect 422352 109024 422484 109052
rect 422352 109012 422358 109024
rect 422478 109012 422484 109024
rect 422536 109012 422542 109064
rect 427814 109012 427820 109064
rect 427872 109052 427878 109064
rect 427998 109052 428004 109064
rect 427872 109024 428004 109052
rect 427872 109012 427878 109024
rect 427998 109012 428004 109024
rect 428056 109012 428062 109064
rect 466638 109052 466644 109064
rect 466564 109024 466644 109052
rect 243170 108984 243176 108996
rect 243096 108956 243176 108984
rect 243170 108944 243176 108956
rect 243228 108944 243234 108996
rect 254118 108984 254124 108996
rect 254079 108956 254124 108984
rect 254118 108944 254124 108956
rect 254176 108944 254182 108996
rect 342438 108984 342444 108996
rect 342399 108956 342444 108984
rect 342438 108944 342444 108956
rect 342496 108944 342502 108996
rect 397638 108944 397644 108996
rect 397696 108944 397702 108996
rect 408696 108984 408724 109012
rect 466564 108996 466592 109024
rect 466638 109012 466644 109024
rect 466696 109012 466702 109064
rect 408770 108984 408776 108996
rect 408696 108956 408776 108984
rect 408770 108944 408776 108956
rect 408828 108944 408834 108996
rect 466546 108944 466552 108996
rect 466604 108944 466610 108996
rect 370130 106332 370136 106344
rect 370091 106304 370136 106332
rect 370130 106292 370136 106304
rect 370188 106292 370194 106344
rect 241790 106224 241796 106276
rect 241848 106264 241854 106276
rect 241974 106264 241980 106276
rect 241848 106236 241980 106264
rect 241848 106224 241854 106236
rect 241974 106224 241980 106236
rect 242032 106224 242038 106276
rect 254118 106224 254124 106276
rect 254176 106264 254182 106276
rect 254210 106264 254216 106276
rect 254176 106236 254216 106264
rect 254176 106224 254182 106236
rect 254210 106224 254216 106236
rect 254268 106224 254274 106276
rect 281810 106224 281816 106276
rect 281868 106264 281874 106276
rect 281902 106264 281908 106276
rect 281868 106236 281908 106264
rect 281868 106224 281874 106236
rect 281902 106224 281908 106236
rect 281960 106224 281966 106276
rect 283098 106264 283104 106276
rect 283059 106236 283104 106264
rect 283098 106224 283104 106236
rect 283156 106224 283162 106276
rect 305178 106264 305184 106276
rect 305139 106236 305184 106264
rect 305178 106224 305184 106236
rect 305236 106224 305242 106276
rect 308030 106224 308036 106276
rect 308088 106264 308094 106276
rect 308214 106264 308220 106276
rect 308088 106236 308220 106264
rect 308088 106224 308094 106236
rect 308214 106224 308220 106236
rect 308272 106224 308278 106276
rect 310698 106264 310704 106276
rect 310659 106236 310704 106264
rect 310698 106224 310704 106236
rect 310756 106224 310762 106276
rect 330018 106224 330024 106276
rect 330076 106264 330082 106276
rect 330202 106264 330208 106276
rect 330076 106236 330208 106264
rect 330076 106224 330082 106236
rect 330202 106224 330208 106236
rect 330260 106224 330266 106276
rect 331398 106224 331404 106276
rect 331456 106264 331462 106276
rect 331490 106264 331496 106276
rect 331456 106236 331496 106264
rect 331456 106224 331462 106236
rect 331490 106224 331496 106236
rect 331548 106224 331554 106276
rect 346578 106264 346584 106276
rect 346539 106236 346584 106264
rect 346578 106224 346584 106236
rect 346636 106224 346642 106276
rect 352006 106224 352012 106276
rect 352064 106264 352070 106276
rect 352190 106264 352196 106276
rect 352064 106236 352196 106264
rect 352064 106224 352070 106236
rect 352190 106224 352196 106236
rect 352248 106224 352254 106276
rect 353478 106224 353484 106276
rect 353536 106264 353542 106276
rect 353570 106264 353576 106276
rect 353536 106236 353576 106264
rect 353536 106224 353542 106236
rect 353570 106224 353576 106236
rect 353628 106224 353634 106276
rect 364518 106224 364524 106276
rect 364576 106264 364582 106276
rect 364610 106264 364616 106276
rect 364576 106236 364616 106264
rect 364576 106224 364582 106236
rect 364610 106224 364616 106236
rect 364668 106224 364674 106276
rect 376938 106264 376944 106276
rect 376899 106236 376944 106264
rect 376938 106224 376944 106236
rect 376996 106224 377002 106276
rect 393222 106224 393228 106276
rect 393280 106264 393286 106276
rect 393406 106264 393412 106276
rect 393280 106236 393412 106264
rect 393280 106224 393286 106236
rect 393406 106224 393412 106236
rect 393464 106224 393470 106276
rect 422386 106264 422392 106276
rect 422347 106236 422392 106264
rect 422386 106224 422392 106236
rect 422444 106224 422450 106276
rect 427906 106264 427912 106276
rect 427867 106236 427912 106264
rect 427906 106224 427912 106236
rect 427964 106224 427970 106276
rect 231946 106156 231952 106208
rect 232004 106196 232010 106208
rect 232130 106196 232136 106208
rect 232004 106168 232136 106196
rect 232004 106156 232010 106168
rect 232130 106156 232136 106168
rect 232188 106156 232194 106208
rect 236270 106156 236276 106208
rect 236328 106196 236334 106208
rect 236546 106196 236552 106208
rect 236328 106168 236552 106196
rect 236328 106156 236334 106168
rect 236546 106156 236552 106168
rect 236604 106156 236610 106208
rect 243170 106196 243176 106208
rect 243131 106168 243176 106196
rect 243170 106156 243176 106168
rect 243228 106156 243234 106208
rect 252738 106196 252744 106208
rect 252699 106168 252744 106196
rect 252738 106156 252744 106168
rect 252796 106156 252802 106208
rect 266998 104972 267004 104984
rect 266959 104944 267004 104972
rect 266998 104932 267004 104944
rect 267056 104932 267062 104984
rect 356422 104972 356428 104984
rect 356383 104944 356428 104972
rect 356422 104932 356428 104944
rect 356480 104932 356486 104984
rect 298189 104907 298247 104913
rect 298189 104873 298201 104907
rect 298235 104904 298247 104907
rect 298370 104904 298376 104916
rect 298235 104876 298376 104904
rect 298235 104873 298247 104876
rect 298189 104867 298247 104873
rect 298370 104864 298376 104876
rect 298428 104864 298434 104916
rect 318978 104904 318984 104916
rect 318939 104876 318984 104904
rect 318978 104864 318984 104876
rect 319036 104864 319042 104916
rect 327169 104907 327227 104913
rect 327169 104873 327181 104907
rect 327215 104904 327227 104907
rect 327258 104904 327264 104916
rect 327215 104876 327264 104904
rect 327215 104873 327227 104876
rect 327169 104867 327227 104873
rect 327258 104864 327264 104876
rect 327316 104864 327322 104916
rect 334342 104864 334348 104916
rect 334400 104904 334406 104916
rect 334434 104904 334440 104916
rect 334400 104876 334440 104904
rect 334400 104864 334406 104876
rect 334434 104864 334440 104876
rect 334492 104864 334498 104916
rect 387978 104904 387984 104916
rect 387939 104876 387984 104904
rect 387978 104864 387984 104876
rect 388036 104864 388042 104916
rect 232130 104836 232136 104848
rect 232091 104808 232136 104836
rect 232130 104796 232136 104808
rect 232188 104796 232194 104848
rect 266998 104836 267004 104848
rect 266959 104808 267004 104836
rect 266998 104796 267004 104808
rect 267056 104796 267062 104848
rect 324406 104796 324412 104848
rect 324464 104836 324470 104848
rect 324682 104836 324688 104848
rect 324464 104808 324688 104836
rect 324464 104796 324470 104808
rect 324682 104796 324688 104808
rect 324740 104796 324746 104848
rect 353478 104836 353484 104848
rect 353439 104808 353484 104836
rect 353478 104796 353484 104808
rect 353536 104796 353542 104848
rect 356422 104836 356428 104848
rect 356383 104808 356428 104836
rect 356422 104796 356428 104808
rect 356480 104796 356486 104848
rect 408681 104839 408739 104845
rect 408681 104805 408693 104839
rect 408727 104836 408739 104839
rect 408770 104836 408776 104848
rect 408727 104808 408776 104836
rect 408727 104805 408739 104808
rect 408681 104799 408739 104805
rect 408770 104796 408776 104808
rect 408828 104796 408834 104848
rect 451550 104836 451556 104848
rect 451511 104808 451556 104836
rect 451550 104796 451556 104808
rect 451608 104796 451614 104848
rect 292758 103612 292764 103624
rect 292719 103584 292764 103612
rect 292758 103572 292764 103584
rect 292816 103572 292822 103624
rect 292669 103479 292727 103485
rect 292669 103445 292681 103479
rect 292715 103476 292727 103479
rect 292758 103476 292764 103488
rect 292715 103448 292764 103476
rect 292715 103445 292727 103448
rect 292669 103439 292727 103445
rect 292758 103436 292764 103448
rect 292816 103436 292822 103488
rect 334345 103479 334403 103485
rect 334345 103445 334357 103479
rect 334391 103476 334403 103479
rect 334434 103476 334440 103488
rect 334391 103448 334440 103476
rect 334391 103445 334403 103448
rect 334345 103439 334403 103445
rect 334434 103436 334440 103448
rect 334492 103436 334498 103488
rect 295613 102187 295671 102193
rect 295613 102153 295625 102187
rect 295659 102184 295671 102187
rect 295702 102184 295708 102196
rect 295659 102156 295708 102184
rect 295659 102153 295671 102156
rect 295613 102147 295671 102153
rect 295702 102144 295708 102156
rect 295760 102144 295766 102196
rect 270862 102116 270868 102128
rect 270823 102088 270868 102116
rect 270862 102076 270868 102088
rect 270920 102076 270926 102128
rect 260834 100036 260840 100088
rect 260892 100076 260898 100088
rect 261018 100076 261024 100088
rect 260892 100048 261024 100076
rect 260892 100036 260898 100048
rect 261018 100036 261024 100048
rect 261076 100036 261082 100088
rect 327258 99492 327264 99544
rect 327316 99492 327322 99544
rect 298370 99464 298376 99476
rect 298331 99436 298376 99464
rect 298370 99424 298376 99436
rect 298428 99424 298434 99476
rect 321738 99424 321744 99476
rect 321796 99424 321802 99476
rect 230750 99356 230756 99408
rect 230808 99356 230814 99408
rect 277578 99356 277584 99408
rect 277636 99356 277642 99408
rect 318978 99356 318984 99408
rect 319036 99356 319042 99408
rect 230768 99328 230796 99356
rect 230842 99328 230848 99340
rect 230768 99300 230848 99328
rect 230842 99288 230848 99300
rect 230900 99288 230906 99340
rect 277596 99328 277624 99356
rect 277670 99328 277676 99340
rect 277596 99300 277676 99328
rect 277670 99288 277676 99300
rect 277728 99288 277734 99340
rect 318996 99328 319024 99356
rect 321756 99340 321784 99424
rect 327276 99340 327304 99492
rect 416866 99356 416872 99408
rect 416924 99356 416930 99408
rect 466546 99356 466552 99408
rect 466604 99356 466610 99408
rect 472066 99356 472072 99408
rect 472124 99356 472130 99408
rect 319070 99328 319076 99340
rect 318996 99300 319076 99328
rect 319070 99288 319076 99300
rect 319128 99288 319134 99340
rect 321738 99288 321744 99340
rect 321796 99288 321802 99340
rect 327258 99288 327264 99340
rect 327316 99288 327322 99340
rect 416774 99288 416780 99340
rect 416832 99328 416838 99340
rect 416884 99328 416912 99356
rect 422386 99328 422392 99340
rect 416832 99300 416912 99328
rect 422347 99300 422392 99328
rect 416832 99288 416838 99300
rect 422386 99288 422392 99300
rect 422444 99288 422450 99340
rect 427906 99328 427912 99340
rect 427867 99300 427912 99328
rect 427906 99288 427912 99300
rect 427964 99288 427970 99340
rect 466454 99288 466460 99340
rect 466512 99328 466518 99340
rect 466564 99328 466592 99356
rect 466512 99300 466592 99328
rect 466512 99288 466518 99300
rect 471974 99288 471980 99340
rect 472032 99328 472038 99340
rect 472084 99328 472112 99356
rect 472032 99300 472112 99328
rect 472032 99288 472038 99300
rect 243170 96744 243176 96756
rect 243131 96716 243176 96744
rect 243170 96704 243176 96716
rect 243228 96704 243234 96756
rect 252738 96676 252744 96688
rect 252699 96648 252744 96676
rect 252738 96636 252744 96648
rect 252796 96636 252802 96688
rect 283098 96676 283104 96688
rect 283059 96648 283104 96676
rect 283098 96636 283104 96648
rect 283156 96636 283162 96688
rect 305178 96676 305184 96688
rect 305139 96648 305184 96676
rect 305178 96636 305184 96648
rect 305236 96636 305242 96688
rect 310698 96676 310704 96688
rect 310659 96648 310704 96676
rect 310698 96636 310704 96648
rect 310756 96636 310762 96688
rect 346578 96676 346584 96688
rect 346539 96648 346584 96676
rect 346578 96636 346584 96648
rect 346636 96636 346642 96688
rect 376938 96676 376944 96688
rect 376899 96648 376944 96676
rect 376938 96636 376944 96648
rect 376996 96636 377002 96688
rect 230842 96608 230848 96620
rect 230803 96580 230848 96608
rect 230842 96568 230848 96580
rect 230900 96568 230906 96620
rect 243078 96568 243084 96620
rect 243136 96608 243142 96620
rect 243170 96608 243176 96620
rect 243136 96580 243176 96608
rect 243136 96568 243142 96580
rect 243170 96568 243176 96580
rect 243228 96568 243234 96620
rect 281810 96568 281816 96620
rect 281868 96608 281874 96620
rect 281994 96608 282000 96620
rect 281868 96580 282000 96608
rect 281868 96568 281874 96580
rect 281994 96568 282000 96580
rect 282052 96568 282058 96620
rect 232133 95251 232191 95257
rect 232133 95217 232145 95251
rect 232179 95248 232191 95251
rect 232222 95248 232228 95260
rect 232179 95220 232228 95248
rect 232179 95217 232191 95220
rect 232133 95211 232191 95217
rect 232222 95208 232228 95220
rect 232280 95208 232286 95260
rect 267001 95251 267059 95257
rect 267001 95217 267013 95251
rect 267047 95248 267059 95251
rect 267090 95248 267096 95260
rect 267047 95220 267096 95248
rect 267047 95217 267059 95220
rect 267001 95211 267059 95217
rect 267090 95208 267096 95220
rect 267148 95208 267154 95260
rect 298370 95248 298376 95260
rect 298331 95220 298376 95248
rect 298370 95208 298376 95220
rect 298428 95208 298434 95260
rect 353478 95248 353484 95260
rect 353439 95220 353484 95248
rect 353478 95208 353484 95220
rect 353536 95208 353542 95260
rect 356425 95251 356483 95257
rect 356425 95217 356437 95251
rect 356471 95248 356483 95251
rect 356606 95248 356612 95260
rect 356471 95220 356612 95248
rect 356471 95217 356483 95220
rect 356425 95211 356483 95217
rect 356606 95208 356612 95220
rect 356664 95208 356670 95260
rect 408678 95248 408684 95260
rect 408639 95220 408684 95248
rect 408678 95208 408684 95220
rect 408736 95208 408742 95260
rect 451550 95248 451556 95260
rect 451511 95220 451556 95248
rect 451550 95208 451556 95220
rect 451608 95208 451614 95260
rect 265158 95180 265164 95192
rect 265119 95152 265164 95180
rect 265158 95140 265164 95152
rect 265216 95140 265222 95192
rect 324498 95180 324504 95192
rect 324459 95152 324504 95180
rect 324498 95140 324504 95152
rect 324556 95140 324562 95192
rect 327258 95180 327264 95192
rect 327219 95152 327264 95180
rect 327258 95140 327264 95152
rect 327316 95140 327322 95192
rect 387978 95180 387984 95192
rect 387939 95152 387984 95180
rect 387978 95140 387984 95152
rect 388036 95140 388042 95192
rect 393222 95180 393228 95192
rect 393183 95152 393228 95180
rect 393222 95140 393228 95152
rect 393280 95140 393286 95192
rect 292666 93888 292672 93900
rect 292627 93860 292672 93888
rect 292666 93848 292672 93860
rect 292724 93848 292730 93900
rect 334342 93888 334348 93900
rect 334303 93860 334348 93888
rect 334342 93848 334348 93860
rect 334400 93848 334406 93900
rect 270865 92531 270923 92537
rect 270865 92497 270877 92531
rect 270911 92528 270923 92531
rect 270954 92528 270960 92540
rect 270911 92500 270960 92528
rect 270911 92497 270923 92500
rect 270865 92491 270923 92497
rect 270954 92488 270960 92500
rect 271012 92488 271018 92540
rect 233326 89700 233332 89752
rect 233384 89740 233390 89752
rect 233510 89740 233516 89752
rect 233384 89712 233516 89740
rect 233384 89700 233390 89712
rect 233510 89700 233516 89712
rect 233568 89700 233574 89752
rect 298370 89740 298376 89752
rect 298331 89712 298376 89740
rect 298370 89700 298376 89712
rect 298428 89700 298434 89752
rect 408678 89700 408684 89752
rect 408736 89700 408742 89752
rect 422294 89700 422300 89752
rect 422352 89740 422358 89752
rect 422478 89740 422484 89752
rect 422352 89712 422484 89740
rect 422352 89700 422358 89712
rect 422478 89700 422484 89712
rect 422536 89700 422542 89752
rect 427814 89700 427820 89752
rect 427872 89740 427878 89752
rect 427998 89740 428004 89752
rect 427872 89712 428004 89740
rect 427872 89700 427878 89712
rect 427998 89700 428004 89712
rect 428056 89700 428062 89752
rect 230842 89672 230848 89684
rect 230803 89644 230848 89672
rect 230842 89632 230848 89644
rect 230900 89632 230906 89684
rect 408696 89604 408724 89700
rect 408770 89604 408776 89616
rect 408696 89576 408776 89604
rect 408770 89564 408776 89576
rect 408828 89564 408834 89616
rect 241790 86952 241796 86964
rect 241751 86924 241796 86952
rect 241790 86912 241796 86924
rect 241848 86912 241854 86964
rect 271966 86912 271972 86964
rect 272024 86952 272030 86964
rect 272058 86952 272064 86964
rect 272024 86924 272064 86952
rect 272024 86912 272030 86924
rect 272058 86912 272064 86924
rect 272116 86912 272122 86964
rect 305178 86952 305184 86964
rect 305139 86924 305184 86952
rect 305178 86912 305184 86924
rect 305236 86912 305242 86964
rect 308030 86952 308036 86964
rect 307991 86924 308036 86952
rect 308030 86912 308036 86924
rect 308088 86912 308094 86964
rect 309318 86952 309324 86964
rect 309279 86924 309324 86952
rect 309318 86912 309324 86924
rect 309376 86912 309382 86964
rect 310698 86952 310704 86964
rect 310659 86924 310704 86952
rect 310698 86912 310704 86924
rect 310756 86912 310762 86964
rect 318978 86912 318984 86964
rect 319036 86912 319042 86964
rect 342438 86952 342444 86964
rect 342399 86924 342444 86952
rect 342438 86912 342444 86924
rect 342496 86912 342502 86964
rect 346578 86952 346584 86964
rect 346539 86924 346584 86952
rect 346578 86912 346584 86924
rect 346636 86912 346642 86964
rect 352006 86912 352012 86964
rect 352064 86912 352070 86964
rect 353478 86912 353484 86964
rect 353536 86952 353542 86964
rect 353570 86952 353576 86964
rect 353536 86924 353576 86952
rect 353536 86912 353542 86924
rect 353570 86912 353576 86924
rect 353628 86912 353634 86964
rect 357618 86912 357624 86964
rect 357676 86952 357682 86964
rect 357802 86952 357808 86964
rect 357676 86924 357808 86952
rect 357676 86912 357682 86924
rect 357802 86912 357808 86924
rect 357860 86912 357866 86964
rect 397638 86952 397644 86964
rect 397599 86924 397644 86952
rect 397638 86912 397644 86924
rect 397696 86912 397702 86964
rect 400309 86955 400367 86961
rect 400309 86921 400321 86955
rect 400355 86952 400367 86955
rect 400398 86952 400404 86964
rect 400355 86924 400404 86952
rect 400355 86921 400367 86924
rect 400309 86915 400367 86921
rect 400398 86912 400404 86924
rect 400456 86912 400462 86964
rect 422386 86952 422392 86964
rect 422347 86924 422392 86952
rect 422386 86912 422392 86924
rect 422444 86912 422450 86964
rect 427906 86952 427912 86964
rect 427867 86924 427912 86952
rect 427906 86912 427912 86924
rect 427964 86912 427970 86964
rect 433429 86955 433487 86961
rect 433429 86921 433441 86955
rect 433475 86952 433487 86955
rect 433518 86952 433524 86964
rect 433475 86924 433524 86952
rect 433475 86921 433487 86924
rect 433429 86915 433487 86921
rect 433518 86912 433524 86924
rect 433576 86912 433582 86964
rect 243078 86844 243084 86896
rect 243136 86884 243142 86896
rect 243262 86884 243268 86896
rect 243136 86856 243268 86884
rect 243136 86844 243142 86856
rect 243262 86844 243268 86856
rect 243320 86844 243326 86896
rect 252738 86884 252744 86896
rect 252699 86856 252744 86884
rect 252738 86844 252744 86856
rect 252796 86844 252802 86896
rect 254118 86884 254124 86896
rect 254079 86856 254124 86884
rect 254118 86844 254124 86856
rect 254176 86844 254182 86896
rect 259638 86884 259644 86896
rect 259599 86856 259644 86884
rect 259638 86844 259644 86856
rect 259696 86844 259702 86896
rect 318996 86884 319024 86912
rect 319070 86884 319076 86896
rect 318996 86856 319076 86884
rect 319070 86844 319076 86856
rect 319128 86844 319134 86896
rect 331398 86884 331404 86896
rect 331359 86856 331404 86884
rect 331398 86844 331404 86856
rect 331456 86844 331462 86896
rect 334342 86884 334348 86896
rect 334303 86856 334348 86884
rect 334342 86844 334348 86856
rect 334400 86844 334406 86896
rect 352024 86884 352052 86912
rect 352098 86884 352104 86896
rect 352024 86856 352104 86884
rect 352098 86844 352104 86856
rect 352156 86844 352162 86896
rect 364518 86884 364524 86896
rect 364479 86856 364524 86884
rect 364518 86844 364524 86856
rect 364576 86844 364582 86896
rect 370038 86884 370044 86896
rect 369999 86856 370044 86884
rect 370038 86844 370044 86856
rect 370096 86844 370102 86896
rect 386598 86884 386604 86896
rect 386559 86856 386604 86884
rect 386598 86844 386604 86856
rect 386656 86844 386662 86896
rect 392118 86884 392124 86896
rect 392079 86856 392124 86884
rect 392118 86844 392124 86856
rect 392176 86844 392182 86896
rect 260742 85620 260748 85672
rect 260800 85660 260806 85672
rect 260800 85632 261064 85660
rect 260800 85620 260806 85632
rect 261036 85604 261064 85632
rect 261018 85552 261024 85604
rect 261076 85552 261082 85604
rect 265158 85592 265164 85604
rect 265119 85564 265164 85592
rect 265158 85552 265164 85564
rect 265216 85552 265222 85604
rect 298370 85592 298376 85604
rect 298331 85564 298376 85592
rect 298370 85552 298376 85564
rect 298428 85552 298434 85604
rect 324498 85592 324504 85604
rect 324459 85564 324504 85592
rect 324498 85552 324504 85564
rect 324556 85552 324562 85604
rect 327258 85592 327264 85604
rect 327219 85564 327264 85592
rect 327258 85552 327264 85564
rect 327316 85552 327322 85604
rect 330018 85552 330024 85604
rect 330076 85592 330082 85604
rect 330110 85592 330116 85604
rect 330076 85564 330116 85592
rect 330076 85552 330082 85564
rect 330110 85552 330116 85564
rect 330168 85552 330174 85604
rect 356422 85552 356428 85604
rect 356480 85592 356486 85604
rect 356606 85592 356612 85604
rect 356480 85564 356612 85592
rect 356480 85552 356486 85564
rect 356606 85552 356612 85564
rect 356664 85552 356670 85604
rect 387978 85592 387984 85604
rect 387939 85564 387984 85592
rect 387978 85552 387984 85564
rect 388036 85552 388042 85604
rect 393225 85595 393283 85601
rect 393225 85561 393237 85595
rect 393271 85592 393283 85595
rect 393406 85592 393412 85604
rect 393271 85564 393412 85592
rect 393271 85561 393283 85564
rect 393225 85555 393283 85561
rect 393406 85552 393412 85564
rect 393464 85552 393470 85604
rect 231946 85524 231952 85536
rect 231907 85496 231952 85524
rect 231946 85484 231952 85496
rect 232004 85484 232010 85536
rect 236270 85524 236276 85536
rect 236231 85496 236276 85524
rect 236270 85484 236276 85496
rect 236328 85484 236334 85536
rect 353478 85484 353484 85536
rect 353536 85484 353542 85536
rect 451461 85527 451519 85533
rect 451461 85493 451473 85527
rect 451507 85524 451519 85527
rect 451550 85524 451556 85536
rect 451507 85496 451556 85524
rect 451507 85493 451519 85496
rect 451461 85487 451519 85493
rect 451550 85484 451556 85496
rect 451608 85484 451614 85536
rect 466546 85524 466552 85536
rect 466507 85496 466552 85524
rect 466546 85484 466552 85496
rect 466604 85484 466610 85536
rect 353496 85456 353524 85484
rect 353570 85456 353576 85468
rect 353496 85428 353576 85456
rect 353570 85416 353576 85428
rect 353628 85416 353634 85468
rect 270681 82807 270739 82813
rect 270681 82773 270693 82807
rect 270727 82804 270739 82807
rect 270954 82804 270960 82816
rect 270727 82776 270960 82804
rect 270727 82773 270739 82776
rect 270681 82767 270739 82773
rect 270954 82764 270960 82776
rect 271012 82764 271018 82816
rect 358998 82804 359004 82816
rect 358959 82776 359004 82804
rect 358998 82764 359004 82776
rect 359056 82764 359062 82816
rect 408770 82124 408776 82136
rect 408731 82096 408776 82124
rect 408770 82084 408776 82096
rect 408828 82084 408834 82136
rect 298281 80767 298339 80773
rect 298281 80733 298293 80767
rect 298327 80764 298339 80767
rect 298370 80764 298376 80776
rect 298327 80736 298376 80764
rect 298327 80733 298339 80736
rect 298281 80727 298339 80733
rect 298370 80724 298376 80736
rect 298428 80724 298434 80776
rect 346486 80724 346492 80776
rect 346544 80764 346550 80776
rect 346581 80767 346639 80773
rect 346581 80764 346593 80767
rect 346544 80736 346593 80764
rect 346544 80724 346550 80736
rect 346581 80733 346593 80736
rect 346627 80733 346639 80767
rect 472066 80764 472072 80776
rect 472027 80736 472072 80764
rect 346581 80727 346639 80733
rect 472066 80724 472072 80736
rect 472124 80724 472130 80776
rect 230934 80152 230940 80164
rect 230895 80124 230940 80152
rect 230934 80112 230940 80124
rect 230992 80112 230998 80164
rect 277486 80152 277492 80164
rect 277412 80124 277492 80152
rect 244458 80044 244464 80096
rect 244516 80044 244522 80096
rect 244476 79960 244504 80044
rect 277412 80028 277440 80124
rect 277486 80112 277492 80124
rect 277544 80112 277550 80164
rect 294138 80112 294144 80164
rect 294196 80112 294202 80164
rect 295518 80112 295524 80164
rect 295576 80152 295582 80164
rect 295702 80152 295708 80164
rect 295576 80124 295708 80152
rect 295576 80112 295582 80124
rect 295702 80112 295708 80124
rect 295760 80112 295766 80164
rect 294156 80028 294184 80112
rect 371418 80044 371424 80096
rect 371476 80044 371482 80096
rect 376938 80044 376944 80096
rect 376996 80044 377002 80096
rect 382458 80044 382464 80096
rect 382516 80044 382522 80096
rect 277394 79976 277400 80028
rect 277452 79976 277458 80028
rect 294138 79976 294144 80028
rect 294196 79976 294202 80028
rect 371436 79960 371464 80044
rect 376956 79960 376984 80044
rect 382476 79960 382504 80044
rect 244458 79908 244464 79960
rect 244516 79908 244522 79960
rect 371418 79908 371424 79960
rect 371476 79908 371482 79960
rect 376938 79908 376944 79960
rect 376996 79908 377002 79960
rect 382458 79908 382464 79960
rect 382516 79908 382522 79960
rect 2774 79840 2780 79892
rect 2832 79880 2838 79892
rect 4798 79880 4804 79892
rect 2832 79852 4804 79880
rect 2832 79840 2838 79852
rect 4798 79840 4804 79852
rect 4856 79840 4862 79892
rect 281810 77324 281816 77376
rect 281868 77364 281874 77376
rect 281994 77364 282000 77376
rect 281868 77336 282000 77364
rect 281868 77324 281874 77336
rect 281994 77324 282000 77336
rect 282052 77324 282058 77376
rect 327258 77364 327264 77376
rect 327184 77336 327264 77364
rect 230934 77296 230940 77308
rect 230895 77268 230940 77296
rect 230934 77256 230940 77268
rect 230992 77256 230998 77308
rect 241790 77296 241796 77308
rect 241751 77268 241796 77296
rect 241790 77256 241796 77268
rect 241848 77256 241854 77308
rect 252738 77296 252744 77308
rect 252699 77268 252744 77296
rect 252738 77256 252744 77268
rect 252796 77256 252802 77308
rect 254118 77296 254124 77308
rect 254079 77268 254124 77296
rect 254118 77256 254124 77268
rect 254176 77256 254182 77308
rect 259638 77296 259644 77308
rect 259599 77268 259644 77296
rect 259638 77256 259644 77268
rect 259696 77256 259702 77308
rect 287146 77256 287152 77308
rect 287204 77296 287210 77308
rect 287238 77296 287244 77308
rect 287204 77268 287244 77296
rect 287204 77256 287210 77268
rect 287238 77256 287244 77268
rect 287296 77256 287302 77308
rect 305178 77296 305184 77308
rect 305139 77268 305184 77296
rect 305178 77256 305184 77268
rect 305236 77256 305242 77308
rect 308030 77296 308036 77308
rect 307991 77268 308036 77296
rect 308030 77256 308036 77268
rect 308088 77256 308094 77308
rect 309318 77296 309324 77308
rect 309279 77268 309324 77296
rect 309318 77256 309324 77268
rect 309376 77256 309382 77308
rect 310698 77296 310704 77308
rect 310659 77268 310704 77296
rect 310698 77256 310704 77268
rect 310756 77256 310762 77308
rect 327184 77240 327212 77336
rect 327258 77324 327264 77336
rect 327316 77324 327322 77376
rect 347866 77324 347872 77376
rect 347924 77324 347930 77376
rect 416774 77324 416780 77376
rect 416832 77364 416838 77376
rect 416958 77364 416964 77376
rect 416832 77336 416964 77364
rect 416832 77324 416838 77336
rect 416958 77324 416964 77336
rect 417016 77324 417022 77376
rect 331398 77296 331404 77308
rect 331359 77268 331404 77296
rect 331398 77256 331404 77268
rect 331456 77256 331462 77308
rect 334342 77296 334348 77308
rect 334303 77268 334348 77296
rect 334342 77256 334348 77268
rect 334400 77256 334406 77308
rect 342438 77296 342444 77308
rect 342399 77268 342444 77296
rect 342438 77256 342444 77268
rect 342496 77256 342502 77308
rect 347884 77240 347912 77324
rect 364518 77296 364524 77308
rect 364479 77268 364524 77296
rect 364518 77256 364524 77268
rect 364576 77256 364582 77308
rect 370038 77296 370044 77308
rect 369999 77268 370044 77296
rect 370038 77256 370044 77268
rect 370096 77256 370102 77308
rect 381078 77256 381084 77308
rect 381136 77296 381142 77308
rect 381170 77296 381176 77308
rect 381136 77268 381176 77296
rect 381136 77256 381142 77268
rect 381170 77256 381176 77268
rect 381228 77256 381234 77308
rect 386598 77296 386604 77308
rect 386559 77268 386604 77296
rect 386598 77256 386604 77268
rect 386656 77256 386662 77308
rect 392118 77296 392124 77308
rect 392079 77268 392124 77296
rect 392118 77256 392124 77268
rect 392176 77256 392182 77308
rect 397638 77296 397644 77308
rect 397599 77268 397644 77296
rect 397638 77256 397644 77268
rect 397696 77256 397702 77308
rect 400306 77296 400312 77308
rect 400267 77268 400312 77296
rect 400306 77256 400312 77268
rect 400364 77256 400370 77308
rect 408770 77296 408776 77308
rect 408731 77268 408776 77296
rect 408770 77256 408776 77268
rect 408828 77256 408834 77308
rect 422389 77299 422447 77305
rect 422389 77265 422401 77299
rect 422435 77296 422447 77299
rect 422478 77296 422484 77308
rect 422435 77268 422484 77296
rect 422435 77265 422447 77268
rect 422389 77259 422447 77265
rect 422478 77256 422484 77268
rect 422536 77256 422542 77308
rect 427909 77299 427967 77305
rect 427909 77265 427921 77299
rect 427955 77296 427967 77299
rect 427998 77296 428004 77308
rect 427955 77268 428004 77296
rect 427955 77265 427967 77268
rect 427909 77259 427967 77265
rect 427998 77256 428004 77268
rect 428056 77256 428062 77308
rect 433426 77296 433432 77308
rect 433387 77268 433432 77296
rect 433426 77256 433432 77268
rect 433484 77256 433490 77308
rect 277394 77228 277400 77240
rect 277355 77200 277400 77228
rect 277394 77188 277400 77200
rect 277452 77188 277458 77240
rect 327166 77188 327172 77240
rect 327224 77188 327230 77240
rect 347866 77188 347872 77240
rect 347924 77188 347930 77240
rect 416869 77231 416927 77237
rect 416869 77197 416881 77231
rect 416915 77228 416927 77231
rect 416958 77228 416964 77240
rect 416915 77200 416964 77228
rect 416915 77197 416927 77200
rect 416869 77191 416927 77197
rect 416958 77188 416964 77200
rect 417016 77188 417022 77240
rect 330018 76032 330024 76084
rect 330076 76072 330082 76084
rect 330076 76044 330156 76072
rect 330076 76032 330082 76044
rect 261018 76004 261024 76016
rect 260852 75976 261024 76004
rect 231946 75936 231952 75948
rect 231907 75908 231952 75936
rect 231946 75896 231952 75908
rect 232004 75896 232010 75948
rect 236270 75936 236276 75948
rect 236231 75908 236276 75936
rect 236270 75896 236276 75908
rect 236328 75896 236334 75948
rect 260852 75880 260880 75976
rect 261018 75964 261024 75976
rect 261076 75964 261082 76016
rect 330128 75948 330156 76044
rect 330110 75896 330116 75948
rect 330168 75896 330174 75948
rect 466549 75939 466607 75945
rect 466549 75905 466561 75939
rect 466595 75936 466607 75939
rect 466638 75936 466644 75948
rect 466595 75908 466644 75936
rect 466595 75905 466607 75908
rect 466549 75899 466607 75905
rect 466638 75896 466644 75908
rect 466696 75896 466702 75948
rect 230934 75868 230940 75880
rect 230895 75840 230940 75868
rect 230934 75828 230940 75840
rect 230992 75828 230998 75880
rect 260834 75828 260840 75880
rect 260892 75828 260898 75880
rect 327166 75868 327172 75880
rect 327127 75840 327172 75868
rect 327166 75828 327172 75840
rect 327224 75828 327230 75880
rect 346486 75828 346492 75880
rect 346544 75868 346550 75880
rect 346578 75868 346584 75880
rect 346544 75840 346584 75868
rect 346544 75828 346550 75840
rect 346578 75828 346584 75840
rect 346636 75828 346642 75880
rect 353570 75868 353576 75880
rect 353531 75840 353576 75868
rect 353570 75828 353576 75840
rect 353628 75828 353634 75880
rect 387978 75828 387984 75880
rect 388036 75868 388042 75880
rect 388162 75868 388168 75880
rect 388036 75840 388168 75868
rect 388036 75828 388042 75840
rect 388162 75828 388168 75840
rect 388220 75828 388226 75880
rect 267090 74536 267096 74588
rect 267148 74576 267154 74588
rect 267274 74576 267280 74588
rect 267148 74548 267280 74576
rect 267148 74536 267154 74548
rect 267274 74536 267280 74548
rect 267332 74536 267338 74588
rect 357529 74511 357587 74517
rect 357529 74477 357541 74511
rect 357575 74508 357587 74511
rect 357618 74508 357624 74520
rect 357575 74480 357624 74508
rect 357575 74477 357587 74480
rect 357529 74471 357587 74477
rect 357618 74468 357624 74480
rect 357676 74468 357682 74520
rect 358998 73216 359004 73228
rect 358959 73188 359004 73216
rect 358998 73176 359004 73188
rect 359056 73176 359062 73228
rect 271969 73151 272027 73157
rect 271969 73117 271981 73151
rect 272015 73148 272027 73151
rect 272058 73148 272064 73160
rect 272015 73120 272064 73148
rect 272015 73117 272027 73120
rect 271969 73111 272027 73117
rect 272058 73108 272064 73120
rect 272116 73108 272122 73160
rect 281810 72428 281816 72480
rect 281868 72468 281874 72480
rect 281994 72468 282000 72480
rect 281868 72440 282000 72468
rect 281868 72428 281874 72440
rect 281994 72428 282000 72440
rect 282052 72428 282058 72480
rect 240226 70456 240232 70508
rect 240284 70456 240290 70508
rect 266538 70496 266544 70508
rect 266464 70468 266544 70496
rect 240244 70372 240272 70456
rect 243078 70388 243084 70440
rect 243136 70388 243142 70440
rect 236270 70360 236276 70372
rect 236231 70332 236276 70360
rect 236270 70320 236276 70332
rect 236328 70320 236334 70372
rect 240226 70320 240232 70372
rect 240284 70320 240290 70372
rect 243096 70292 243124 70388
rect 266464 70372 266492 70468
rect 266538 70456 266544 70468
rect 266596 70456 266602 70508
rect 408770 70428 408776 70440
rect 408731 70400 408776 70428
rect 408770 70388 408776 70400
rect 408828 70388 408834 70440
rect 266446 70320 266452 70372
rect 266504 70320 266510 70372
rect 277397 70363 277455 70369
rect 277397 70329 277409 70363
rect 277443 70360 277455 70363
rect 277486 70360 277492 70372
rect 277443 70332 277492 70360
rect 277443 70329 277455 70332
rect 277397 70323 277455 70329
rect 277486 70320 277492 70332
rect 277544 70320 277550 70372
rect 243170 70292 243176 70304
rect 243096 70264 243176 70292
rect 243170 70252 243176 70264
rect 243228 70252 243234 70304
rect 292758 69028 292764 69080
rect 292816 69028 292822 69080
rect 292776 68944 292804 69028
rect 292758 68892 292764 68944
rect 292816 68892 292822 68944
rect 267274 67708 267280 67720
rect 267200 67680 267280 67708
rect 231854 67600 231860 67652
rect 231912 67640 231918 67652
rect 231946 67640 231952 67652
rect 231912 67612 231952 67640
rect 231912 67600 231918 67612
rect 231946 67600 231952 67612
rect 232004 67600 232010 67652
rect 236270 67640 236276 67652
rect 236231 67612 236276 67640
rect 236270 67600 236276 67612
rect 236328 67600 236334 67652
rect 267200 67584 267228 67680
rect 267274 67668 267280 67680
rect 267332 67668 267338 67720
rect 386598 67668 386604 67720
rect 386656 67668 386662 67720
rect 392118 67668 392124 67720
rect 392176 67668 392182 67720
rect 298281 67643 298339 67649
rect 298281 67609 298293 67643
rect 298327 67640 298339 67643
rect 298370 67640 298376 67652
rect 298327 67612 298376 67640
rect 298327 67609 298339 67612
rect 298281 67603 298339 67609
rect 298370 67600 298376 67612
rect 298428 67600 298434 67652
rect 319070 67640 319076 67652
rect 319031 67612 319076 67640
rect 319070 67600 319076 67612
rect 319128 67600 319134 67652
rect 324406 67600 324412 67652
rect 324464 67640 324470 67652
rect 324498 67640 324504 67652
rect 324464 67612 324504 67640
rect 324464 67600 324470 67612
rect 324498 67600 324504 67612
rect 324556 67600 324562 67652
rect 347866 67600 347872 67652
rect 347924 67640 347930 67652
rect 348050 67640 348056 67652
rect 347924 67612 348056 67640
rect 347924 67600 347930 67612
rect 348050 67600 348056 67612
rect 348108 67600 348114 67652
rect 386616 67640 386644 67668
rect 386690 67640 386696 67652
rect 386616 67612 386696 67640
rect 386690 67600 386696 67612
rect 386748 67600 386754 67652
rect 392136 67640 392164 67668
rect 392210 67640 392216 67652
rect 392136 67612 392216 67640
rect 392210 67600 392216 67612
rect 392268 67600 392274 67652
rect 408770 67640 408776 67652
rect 408731 67612 408776 67640
rect 408770 67600 408776 67612
rect 408828 67600 408834 67652
rect 416866 67640 416872 67652
rect 416827 67612 416872 67640
rect 416866 67600 416872 67612
rect 416924 67600 416930 67652
rect 433426 67600 433432 67652
rect 433484 67640 433490 67652
rect 433518 67640 433524 67652
rect 433484 67612 433524 67640
rect 433484 67600 433490 67612
rect 433518 67600 433524 67612
rect 433576 67600 433582 67652
rect 451458 67640 451464 67652
rect 451419 67612 451464 67640
rect 451458 67600 451464 67612
rect 451516 67600 451522 67652
rect 472066 67640 472072 67652
rect 472027 67612 472072 67640
rect 472066 67600 472072 67612
rect 472124 67600 472130 67652
rect 267182 67532 267188 67584
rect 267240 67532 267246 67584
rect 305178 67532 305184 67584
rect 305236 67572 305242 67584
rect 305270 67572 305276 67584
rect 305236 67544 305276 67572
rect 305236 67532 305242 67544
rect 305270 67532 305276 67544
rect 305328 67532 305334 67584
rect 308030 67572 308036 67584
rect 307991 67544 308036 67572
rect 308030 67532 308036 67544
rect 308088 67532 308094 67584
rect 356425 67575 356483 67581
rect 356425 67541 356437 67575
rect 356471 67572 356483 67575
rect 356514 67572 356520 67584
rect 356471 67544 356520 67572
rect 356471 67541 356483 67544
rect 356425 67535 356483 67541
rect 356514 67532 356520 67544
rect 356572 67532 356578 67584
rect 393222 67572 393228 67584
rect 393183 67544 393228 67572
rect 393222 67532 393228 67544
rect 393280 67532 393286 67584
rect 397638 67572 397644 67584
rect 397599 67544 397644 67572
rect 397638 67532 397644 67544
rect 397696 67532 397702 67584
rect 260834 66308 260840 66360
rect 260892 66348 260898 66360
rect 261018 66348 261024 66360
rect 260892 66320 261024 66348
rect 260892 66308 260898 66320
rect 261018 66308 261024 66320
rect 261076 66308 261082 66360
rect 230937 66283 230995 66289
rect 230937 66249 230949 66283
rect 230983 66280 230995 66283
rect 231026 66280 231032 66292
rect 230983 66252 231032 66280
rect 230983 66249 230995 66252
rect 230937 66243 230995 66249
rect 231026 66240 231032 66252
rect 231084 66240 231090 66292
rect 319070 66280 319076 66292
rect 319031 66252 319076 66280
rect 319070 66240 319076 66252
rect 319128 66240 319134 66292
rect 327169 66283 327227 66289
rect 327169 66249 327181 66283
rect 327215 66280 327227 66283
rect 327258 66280 327264 66292
rect 327215 66252 327264 66280
rect 327215 66249 327227 66252
rect 327169 66243 327227 66249
rect 327258 66240 327264 66252
rect 327316 66240 327322 66292
rect 330018 66280 330024 66292
rect 329979 66252 330024 66280
rect 330018 66240 330024 66252
rect 330076 66240 330082 66292
rect 353573 66283 353631 66289
rect 353573 66249 353585 66283
rect 353619 66280 353631 66283
rect 353662 66280 353668 66292
rect 353619 66252 353668 66280
rect 353619 66249 353631 66252
rect 353573 66243 353631 66249
rect 353662 66240 353668 66252
rect 353720 66240 353726 66292
rect 236270 66172 236276 66224
rect 236328 66212 236334 66224
rect 236365 66215 236423 66221
rect 236365 66212 236377 66215
rect 236328 66184 236377 66212
rect 236328 66172 236334 66184
rect 236365 66181 236377 66184
rect 236411 66181 236423 66215
rect 281718 66212 281724 66224
rect 281679 66184 281724 66212
rect 236365 66175 236423 66181
rect 281718 66172 281724 66184
rect 281776 66172 281782 66224
rect 309410 66172 309416 66224
rect 309468 66172 309474 66224
rect 336826 66172 336832 66224
rect 336884 66212 336890 66224
rect 336918 66212 336924 66224
rect 336884 66184 336924 66212
rect 336884 66172 336890 66184
rect 336918 66172 336924 66184
rect 336976 66172 336982 66224
rect 387978 66212 387984 66224
rect 387939 66184 387984 66212
rect 387978 66172 387984 66184
rect 388036 66172 388042 66224
rect 451458 66212 451464 66224
rect 451419 66184 451464 66212
rect 451458 66172 451464 66184
rect 451516 66172 451522 66224
rect 466454 66212 466460 66224
rect 466415 66184 466460 66212
rect 466454 66172 466460 66184
rect 466512 66172 466518 66224
rect 309428 66085 309456 66172
rect 309413 66079 309471 66085
rect 309413 66045 309425 66079
rect 309459 66045 309471 66079
rect 309413 66039 309471 66045
rect 330018 64988 330024 65000
rect 329979 64960 330024 64988
rect 330018 64948 330024 64960
rect 330076 64948 330082 65000
rect 270678 64920 270684 64932
rect 270639 64892 270684 64920
rect 270678 64880 270684 64892
rect 270736 64880 270742 64932
rect 357526 64920 357532 64932
rect 357487 64892 357532 64920
rect 357526 64880 357532 64892
rect 357584 64880 357590 64932
rect 242989 64855 243047 64861
rect 242989 64821 243001 64855
rect 243035 64852 243047 64855
rect 243170 64852 243176 64864
rect 243035 64824 243176 64852
rect 243035 64821 243047 64824
rect 242989 64815 243047 64821
rect 243170 64812 243176 64824
rect 243228 64812 243234 64864
rect 260837 64855 260895 64861
rect 260837 64821 260849 64855
rect 260883 64852 260895 64855
rect 261018 64852 261024 64864
rect 260883 64824 261024 64852
rect 260883 64821 260895 64824
rect 260837 64815 260895 64821
rect 261018 64812 261024 64824
rect 261076 64812 261082 64864
rect 292482 64812 292488 64864
rect 292540 64852 292546 64864
rect 292758 64852 292764 64864
rect 292540 64824 292764 64852
rect 292540 64812 292546 64824
rect 292758 64812 292764 64824
rect 292816 64812 292822 64864
rect 332778 64812 332784 64864
rect 332836 64852 332842 64864
rect 332870 64852 332876 64864
rect 332836 64824 332876 64852
rect 332836 64812 332842 64824
rect 332870 64812 332876 64824
rect 332928 64812 332934 64864
rect 529474 64812 529480 64864
rect 529532 64852 529538 64864
rect 580166 64852 580172 64864
rect 529532 64824 580172 64852
rect 529532 64812 529538 64824
rect 580166 64812 580172 64824
rect 580224 64812 580230 64864
rect 271966 63560 271972 63572
rect 271927 63532 271972 63560
rect 271966 63520 271972 63532
rect 272024 63520 272030 63572
rect 329929 63495 329987 63501
rect 329929 63461 329941 63495
rect 329975 63492 329987 63495
rect 330018 63492 330024 63504
rect 329975 63464 330024 63492
rect 329975 63461 329987 63464
rect 329929 63455 329987 63461
rect 330018 63452 330024 63464
rect 330076 63452 330082 63504
rect 332870 63492 332876 63504
rect 332831 63464 332876 63492
rect 332870 63452 332876 63464
rect 332928 63452 332934 63504
rect 359090 63492 359096 63504
rect 359051 63464 359096 63492
rect 359090 63452 359096 63464
rect 359148 63452 359154 63504
rect 408770 62812 408776 62824
rect 408731 62784 408776 62812
rect 408770 62772 408776 62784
rect 408828 62772 408834 62824
rect 392210 61684 392216 61736
rect 392268 61724 392274 61736
rect 392394 61724 392400 61736
rect 392268 61696 392400 61724
rect 392268 61684 392274 61696
rect 392394 61684 392400 61696
rect 392452 61684 392458 61736
rect 370038 61112 370044 61124
rect 369999 61084 370044 61112
rect 370038 61072 370044 61084
rect 370096 61072 370102 61124
rect 375558 61112 375564 61124
rect 375519 61084 375564 61112
rect 375558 61072 375564 61084
rect 375616 61072 375622 61124
rect 416774 60664 416780 60716
rect 416832 60704 416838 60716
rect 416958 60704 416964 60716
rect 416832 60676 416964 60704
rect 416832 60664 416838 60676
rect 416958 60664 416964 60676
rect 417016 60664 417022 60716
rect 433518 60664 433524 60716
rect 433576 60704 433582 60716
rect 433702 60704 433708 60716
rect 433576 60676 433708 60704
rect 433576 60664 433582 60676
rect 433702 60664 433708 60676
rect 433760 60664 433766 60716
rect 451461 60707 451519 60713
rect 451461 60673 451473 60707
rect 451507 60704 451519 60707
rect 451642 60704 451648 60716
rect 451507 60676 451648 60704
rect 451507 60673 451519 60676
rect 451461 60667 451519 60673
rect 451642 60664 451648 60676
rect 451700 60664 451706 60716
rect 471974 60664 471980 60716
rect 472032 60704 472038 60716
rect 472158 60704 472164 60716
rect 472032 60676 472164 60704
rect 472032 60664 472038 60676
rect 472158 60664 472164 60676
rect 472216 60664 472222 60716
rect 371418 60636 371424 60648
rect 371379 60608 371424 60636
rect 371418 60596 371424 60608
rect 371476 60596 371482 60648
rect 318978 60024 318984 60036
rect 318939 59996 318984 60024
rect 318978 59984 318984 59996
rect 319036 59984 319042 60036
rect 259638 59752 259644 59764
rect 259599 59724 259644 59752
rect 259638 59712 259644 59724
rect 259696 59712 259702 59764
rect 271966 58596 271972 58608
rect 271927 58568 271972 58596
rect 271966 58556 271972 58568
rect 272024 58556 272030 58608
rect 352006 58120 352012 58132
rect 351967 58092 352012 58120
rect 352006 58080 352012 58092
rect 352064 58080 352070 58132
rect 266446 57944 266452 57996
rect 266504 57984 266510 57996
rect 266538 57984 266544 57996
rect 266504 57956 266544 57984
rect 266504 57944 266510 57956
rect 266538 57944 266544 57956
rect 266596 57944 266602 57996
rect 267090 57944 267096 57996
rect 267148 57984 267154 57996
rect 267182 57984 267188 57996
rect 267148 57956 267188 57984
rect 267148 57944 267154 57956
rect 267182 57944 267188 57956
rect 267240 57944 267246 57996
rect 293954 57944 293960 57996
rect 294012 57984 294018 57996
rect 294138 57984 294144 57996
rect 294012 57956 294144 57984
rect 294012 57944 294018 57956
rect 294138 57944 294144 57956
rect 294196 57944 294202 57996
rect 295518 57944 295524 57996
rect 295576 57944 295582 57996
rect 308030 57984 308036 57996
rect 307991 57956 308036 57984
rect 308030 57944 308036 57956
rect 308088 57944 308094 57996
rect 347958 57944 347964 57996
rect 348016 57984 348022 57996
rect 348050 57984 348056 57996
rect 348016 57956 348056 57984
rect 348016 57944 348022 57956
rect 348050 57944 348056 57956
rect 348108 57944 348114 57996
rect 356422 57984 356428 57996
rect 356383 57956 356428 57984
rect 356422 57944 356428 57956
rect 356480 57944 356486 57996
rect 386598 57944 386604 57996
rect 386656 57984 386662 57996
rect 386690 57984 386696 57996
rect 386656 57956 386696 57984
rect 386656 57944 386662 57956
rect 386690 57944 386696 57956
rect 386748 57944 386754 57996
rect 393222 57984 393228 57996
rect 393183 57956 393228 57984
rect 393222 57944 393228 57956
rect 393280 57944 393286 57996
rect 397641 57987 397699 57993
rect 397641 57953 397653 57987
rect 397687 57984 397699 57987
rect 397730 57984 397736 57996
rect 397687 57956 397736 57984
rect 397687 57953 397699 57956
rect 397641 57947 397699 57953
rect 397730 57944 397736 57956
rect 397788 57944 397794 57996
rect 408770 57984 408776 57996
rect 408731 57956 408776 57984
rect 408770 57944 408776 57956
rect 408828 57944 408834 57996
rect 277578 57876 277584 57928
rect 277636 57876 277642 57928
rect 288529 57919 288587 57925
rect 288529 57885 288541 57919
rect 288575 57916 288587 57919
rect 288618 57916 288624 57928
rect 288575 57888 288624 57916
rect 288575 57885 288587 57888
rect 288529 57879 288587 57885
rect 288618 57876 288624 57888
rect 288676 57876 288682 57928
rect 277596 57848 277624 57876
rect 277670 57848 277676 57860
rect 277596 57820 277676 57848
rect 277670 57808 277676 57820
rect 277728 57808 277734 57860
rect 295536 57848 295564 57944
rect 324406 57916 324412 57928
rect 324367 57888 324412 57916
rect 324406 57876 324412 57888
rect 324464 57876 324470 57928
rect 376938 57876 376944 57928
rect 376996 57916 377002 57928
rect 377030 57916 377036 57928
rect 376996 57888 377036 57916
rect 376996 57876 377002 57888
rect 377030 57876 377036 57888
rect 377088 57876 377094 57928
rect 382369 57919 382427 57925
rect 382369 57885 382381 57919
rect 382415 57916 382427 57919
rect 382458 57916 382464 57928
rect 382415 57888 382464 57916
rect 382415 57885 382427 57888
rect 382369 57879 382427 57885
rect 382458 57876 382464 57888
rect 382516 57876 382522 57928
rect 416869 57919 416927 57925
rect 416869 57885 416881 57919
rect 416915 57916 416927 57919
rect 416958 57916 416964 57928
rect 416915 57888 416964 57916
rect 416915 57885 416927 57888
rect 416869 57879 416927 57885
rect 416958 57876 416964 57888
rect 417016 57876 417022 57928
rect 433613 57919 433671 57925
rect 433613 57885 433625 57919
rect 433659 57916 433671 57919
rect 433702 57916 433708 57928
rect 433659 57888 433708 57916
rect 433659 57885 433671 57888
rect 433613 57879 433671 57885
rect 433702 57876 433708 57888
rect 433760 57876 433766 57928
rect 472069 57919 472127 57925
rect 472069 57885 472081 57919
rect 472115 57916 472127 57919
rect 472158 57916 472164 57928
rect 472115 57888 472164 57916
rect 472115 57885 472127 57888
rect 472069 57879 472127 57885
rect 472158 57876 472164 57888
rect 472216 57876 472222 57928
rect 295610 57848 295616 57860
rect 295536 57820 295616 57848
rect 295610 57808 295616 57820
rect 295668 57808 295674 57860
rect 270589 57579 270647 57585
rect 270589 57545 270601 57579
rect 270635 57576 270647 57579
rect 270678 57576 270684 57588
rect 270635 57548 270684 57576
rect 270635 57545 270647 57548
rect 270589 57539 270647 57545
rect 270678 57536 270684 57548
rect 270736 57536 270742 57588
rect 371418 56692 371424 56704
rect 371379 56664 371424 56692
rect 371418 56652 371424 56664
rect 371476 56652 371482 56704
rect 281718 56624 281724 56636
rect 281679 56596 281724 56624
rect 281718 56584 281724 56596
rect 281776 56584 281782 56636
rect 387981 56627 388039 56633
rect 387981 56593 387993 56627
rect 388027 56624 388039 56627
rect 388070 56624 388076 56636
rect 388027 56596 388076 56624
rect 388027 56593 388039 56596
rect 387981 56587 388039 56593
rect 388070 56584 388076 56596
rect 388128 56584 388134 56636
rect 466457 56627 466515 56633
rect 466457 56593 466469 56627
rect 466503 56624 466515 56627
rect 466822 56624 466828 56636
rect 466503 56596 466828 56624
rect 466503 56593 466515 56596
rect 466457 56587 466515 56593
rect 466822 56584 466828 56596
rect 466880 56584 466886 56636
rect 244369 56559 244427 56565
rect 244369 56525 244381 56559
rect 244415 56556 244427 56559
rect 244458 56556 244464 56568
rect 244415 56528 244464 56556
rect 244415 56525 244427 56528
rect 244369 56519 244427 56525
rect 244458 56516 244464 56528
rect 244516 56516 244522 56568
rect 249978 56556 249984 56568
rect 249939 56528 249984 56556
rect 249978 56516 249984 56528
rect 250036 56516 250042 56568
rect 255409 56559 255467 56565
rect 255409 56525 255421 56559
rect 255455 56556 255467 56559
rect 255498 56556 255504 56568
rect 255455 56528 255504 56556
rect 255455 56525 255467 56528
rect 255409 56519 255467 56525
rect 255498 56516 255504 56528
rect 255556 56516 255562 56568
rect 277486 56516 277492 56568
rect 277544 56556 277550 56568
rect 277670 56556 277676 56568
rect 277544 56528 277676 56556
rect 277544 56516 277550 56528
rect 277670 56516 277676 56528
rect 277728 56516 277734 56568
rect 282917 56559 282975 56565
rect 282917 56525 282929 56559
rect 282963 56556 282975 56559
rect 283098 56556 283104 56568
rect 282963 56528 283104 56556
rect 282963 56525 282975 56528
rect 282917 56519 282975 56525
rect 283098 56516 283104 56528
rect 283156 56516 283162 56568
rect 298278 56556 298284 56568
rect 298239 56528 298284 56556
rect 298278 56516 298284 56528
rect 298336 56516 298342 56568
rect 336918 56556 336924 56568
rect 336879 56528 336924 56556
rect 336918 56516 336924 56528
rect 336976 56516 336982 56568
rect 371418 56516 371424 56568
rect 371476 56556 371482 56568
rect 392121 56559 392179 56565
rect 371476 56528 371521 56556
rect 371476 56516 371482 56528
rect 392121 56525 392133 56559
rect 392167 56556 392179 56559
rect 392302 56556 392308 56568
rect 392167 56528 392308 56556
rect 392167 56525 392179 56528
rect 392121 56519 392179 56525
rect 392302 56516 392308 56528
rect 392360 56516 392366 56568
rect 451642 56556 451648 56568
rect 451603 56528 451648 56556
rect 451642 56516 451648 56528
rect 451700 56516 451706 56568
rect 331398 55672 331404 55684
rect 331359 55644 331404 55672
rect 331398 55632 331404 55644
rect 331456 55632 331462 55684
rect 334342 55672 334348 55684
rect 334303 55644 334348 55672
rect 334342 55632 334348 55644
rect 334400 55632 334406 55684
rect 324409 55335 324467 55341
rect 324409 55301 324421 55335
rect 324455 55301 324467 55335
rect 324409 55295 324467 55301
rect 242986 55264 242992 55276
rect 242947 55236 242992 55264
rect 242986 55224 242992 55236
rect 243044 55224 243050 55276
rect 260834 55264 260840 55276
rect 260795 55236 260840 55264
rect 260834 55224 260840 55236
rect 260892 55224 260898 55276
rect 292758 55196 292764 55208
rect 292719 55168 292764 55196
rect 292758 55156 292764 55168
rect 292816 55156 292822 55208
rect 324424 55196 324452 55295
rect 324501 55199 324559 55205
rect 324501 55196 324513 55199
rect 324424 55168 324513 55196
rect 324501 55165 324513 55168
rect 324547 55165 324559 55199
rect 332870 55196 332876 55208
rect 332831 55168 332876 55196
rect 324501 55159 324559 55165
rect 332870 55156 332876 55168
rect 332928 55156 332934 55208
rect 329926 53836 329932 53848
rect 329887 53808 329932 53836
rect 329926 53796 329932 53808
rect 329984 53796 329990 53848
rect 352006 53836 352012 53848
rect 351967 53808 352012 53836
rect 352006 53796 352012 53808
rect 352064 53796 352070 53848
rect 359093 53839 359151 53845
rect 359093 53805 359105 53839
rect 359139 53836 359151 53839
rect 359182 53836 359188 53848
rect 359139 53808 359188 53836
rect 359139 53805 359151 53808
rect 359093 53799 359151 53805
rect 359182 53796 359188 53808
rect 359240 53796 359246 53848
rect 400401 51187 400459 51193
rect 400401 51153 400413 51187
rect 400447 51184 400459 51187
rect 400490 51184 400496 51196
rect 400447 51156 400496 51184
rect 400447 51153 400459 51156
rect 400401 51147 400459 51153
rect 400490 51144 400496 51156
rect 400548 51144 400554 51196
rect 408770 51184 408776 51196
rect 408731 51156 408776 51184
rect 408770 51144 408776 51156
rect 408828 51144 408834 51196
rect 342438 51076 342444 51128
rect 342496 51076 342502 51128
rect 342456 50992 342484 51076
rect 342438 50940 342444 50992
rect 342496 50940 342502 50992
rect 254118 48356 254124 48408
rect 254176 48356 254182 48408
rect 309410 48396 309416 48408
rect 309371 48368 309416 48396
rect 309410 48356 309416 48368
rect 309468 48356 309474 48408
rect 327258 48396 327264 48408
rect 327184 48368 327264 48396
rect 254136 48328 254164 48356
rect 327184 48340 327212 48368
rect 327258 48356 327264 48368
rect 327316 48356 327322 48408
rect 400398 48396 400404 48408
rect 400359 48368 400404 48396
rect 400398 48356 400404 48368
rect 400456 48356 400462 48408
rect 408678 48356 408684 48408
rect 408736 48396 408742 48408
rect 408773 48399 408831 48405
rect 408773 48396 408785 48399
rect 408736 48368 408785 48396
rect 408736 48356 408742 48368
rect 408773 48365 408785 48368
rect 408819 48365 408831 48399
rect 416866 48396 416872 48408
rect 416827 48368 416872 48396
rect 408773 48359 408831 48365
rect 416866 48356 416872 48368
rect 416924 48356 416930 48408
rect 254210 48328 254216 48340
rect 254136 48300 254216 48328
rect 254210 48288 254216 48300
rect 254268 48288 254274 48340
rect 259641 48331 259699 48337
rect 259641 48297 259653 48331
rect 259687 48328 259699 48331
rect 259730 48328 259736 48340
rect 259687 48300 259736 48328
rect 259687 48297 259699 48300
rect 259641 48291 259699 48297
rect 259730 48288 259736 48300
rect 259788 48288 259794 48340
rect 265158 48288 265164 48340
rect 265216 48328 265222 48340
rect 265342 48328 265348 48340
rect 265216 48300 265348 48328
rect 265216 48288 265222 48300
rect 265342 48288 265348 48300
rect 265400 48288 265406 48340
rect 281718 48288 281724 48340
rect 281776 48328 281782 48340
rect 281810 48328 281816 48340
rect 281776 48300 281816 48328
rect 281776 48288 281782 48300
rect 281810 48288 281816 48300
rect 281868 48288 281874 48340
rect 288526 48328 288532 48340
rect 288487 48300 288532 48328
rect 288526 48288 288532 48300
rect 288584 48288 288590 48340
rect 327166 48288 327172 48340
rect 327224 48288 327230 48340
rect 331401 48331 331459 48337
rect 331401 48297 331413 48331
rect 331447 48328 331459 48331
rect 331490 48328 331496 48340
rect 331447 48300 331496 48328
rect 331447 48297 331459 48300
rect 331401 48291 331459 48297
rect 331490 48288 331496 48300
rect 331548 48288 331554 48340
rect 334345 48331 334403 48337
rect 334345 48297 334357 48331
rect 334391 48328 334403 48331
rect 334434 48328 334440 48340
rect 334391 48300 334440 48328
rect 334391 48297 334403 48300
rect 334345 48291 334403 48297
rect 334434 48288 334440 48300
rect 334492 48288 334498 48340
rect 370041 48331 370099 48337
rect 370041 48297 370053 48331
rect 370087 48328 370099 48331
rect 370130 48328 370136 48340
rect 370087 48300 370136 48328
rect 370087 48297 370099 48300
rect 370041 48291 370099 48297
rect 370130 48288 370136 48300
rect 370188 48288 370194 48340
rect 375561 48331 375619 48337
rect 375561 48297 375573 48331
rect 375607 48328 375619 48331
rect 375650 48328 375656 48340
rect 375607 48300 375656 48328
rect 375607 48297 375619 48300
rect 375561 48291 375619 48297
rect 375650 48288 375656 48300
rect 375708 48288 375714 48340
rect 382366 48328 382372 48340
rect 382327 48300 382372 48328
rect 382366 48288 382372 48300
rect 382424 48288 382430 48340
rect 386598 48288 386604 48340
rect 386656 48328 386662 48340
rect 386690 48328 386696 48340
rect 386656 48300 386696 48328
rect 386656 48288 386662 48300
rect 386690 48288 386696 48300
rect 386748 48288 386754 48340
rect 387886 48288 387892 48340
rect 387944 48328 387950 48340
rect 388070 48328 388076 48340
rect 387944 48300 388076 48328
rect 387944 48288 387950 48300
rect 388070 48288 388076 48300
rect 388128 48288 388134 48340
rect 422386 48288 422392 48340
rect 422444 48328 422450 48340
rect 422478 48328 422484 48340
rect 422444 48300 422484 48328
rect 422444 48288 422450 48300
rect 422478 48288 422484 48300
rect 422536 48288 422542 48340
rect 433610 48328 433616 48340
rect 433571 48300 433616 48328
rect 433610 48288 433616 48300
rect 433668 48288 433674 48340
rect 466638 48288 466644 48340
rect 466696 48328 466702 48340
rect 466822 48328 466828 48340
rect 466696 48300 466828 48328
rect 466696 48288 466702 48300
rect 466822 48288 466828 48300
rect 466880 48288 466886 48340
rect 472066 48328 472072 48340
rect 472027 48300 472072 48328
rect 472066 48288 472072 48300
rect 472124 48288 472130 48340
rect 295610 48220 295616 48272
rect 295668 48260 295674 48272
rect 295702 48260 295708 48272
rect 295668 48232 295708 48260
rect 295668 48220 295674 48232
rect 295702 48220 295708 48232
rect 295760 48220 295766 48272
rect 308122 48260 308128 48272
rect 308083 48232 308128 48260
rect 308122 48220 308128 48232
rect 308180 48220 308186 48272
rect 381170 48220 381176 48272
rect 381228 48260 381234 48272
rect 381262 48260 381268 48272
rect 381228 48232 381268 48260
rect 381228 48220 381234 48232
rect 381262 48220 381268 48232
rect 381320 48220 381326 48272
rect 400398 48220 400404 48272
rect 400456 48260 400462 48272
rect 400766 48260 400772 48272
rect 400456 48232 400772 48260
rect 400456 48220 400462 48232
rect 400766 48220 400772 48232
rect 400824 48220 400830 48272
rect 416866 48220 416872 48272
rect 416924 48260 416930 48272
rect 417050 48260 417056 48272
rect 416924 48232 417056 48260
rect 416924 48220 416930 48232
rect 417050 48220 417056 48232
rect 417108 48220 417114 48272
rect 236270 46996 236276 47048
rect 236328 47036 236334 47048
rect 236365 47039 236423 47045
rect 236365 47036 236377 47039
rect 236328 47008 236377 47036
rect 236328 46996 236334 47008
rect 236365 47005 236377 47008
rect 236411 47005 236423 47039
rect 282914 47036 282920 47048
rect 282875 47008 282920 47036
rect 236365 46999 236423 47005
rect 282914 46996 282920 47008
rect 282972 46996 282978 47048
rect 371326 46996 371332 47048
rect 371384 47036 371390 47048
rect 371421 47039 371479 47045
rect 371421 47036 371433 47039
rect 371384 47008 371433 47036
rect 371384 46996 371390 47008
rect 371421 47005 371433 47008
rect 371467 47005 371479 47039
rect 392118 47036 392124 47048
rect 392079 47008 392124 47036
rect 371421 46999 371479 47005
rect 392118 46996 392124 47008
rect 392176 46996 392182 47048
rect 244366 46968 244372 46980
rect 244327 46940 244372 46968
rect 244366 46928 244372 46940
rect 244424 46928 244430 46980
rect 249978 46968 249984 46980
rect 249939 46940 249984 46968
rect 249978 46928 249984 46940
rect 250036 46928 250042 46980
rect 255406 46968 255412 46980
rect 255367 46940 255412 46968
rect 255406 46928 255412 46940
rect 255464 46928 255470 46980
rect 270586 46968 270592 46980
rect 270547 46940 270592 46968
rect 270586 46928 270592 46940
rect 270644 46928 270650 46980
rect 298281 46971 298339 46977
rect 298281 46937 298293 46971
rect 298327 46968 298339 46971
rect 298370 46968 298376 46980
rect 298327 46940 298376 46968
rect 298327 46937 298339 46940
rect 298281 46931 298339 46937
rect 298370 46928 298376 46940
rect 298428 46928 298434 46980
rect 318978 46968 318984 46980
rect 318939 46940 318984 46968
rect 318978 46928 318984 46940
rect 319036 46928 319042 46980
rect 332870 46928 332876 46980
rect 332928 46928 332934 46980
rect 336918 46968 336924 46980
rect 336879 46940 336924 46968
rect 336918 46928 336924 46940
rect 336976 46928 336982 46980
rect 451645 46971 451703 46977
rect 451645 46937 451657 46971
rect 451691 46968 451703 46971
rect 451826 46968 451832 46980
rect 451691 46940 451832 46968
rect 451691 46937 451703 46940
rect 451645 46931 451703 46937
rect 451826 46928 451832 46940
rect 451884 46928 451890 46980
rect 231854 46860 231860 46912
rect 231912 46900 231918 46912
rect 232038 46900 232044 46912
rect 231912 46872 232044 46900
rect 231912 46860 231918 46872
rect 232038 46860 232044 46872
rect 232096 46860 232102 46912
rect 236270 46860 236276 46912
rect 236328 46900 236334 46912
rect 236454 46900 236460 46912
rect 236328 46872 236460 46900
rect 236328 46860 236334 46872
rect 236454 46860 236460 46872
rect 236512 46860 236518 46912
rect 243170 46860 243176 46912
rect 243228 46900 243234 46912
rect 243262 46900 243268 46912
rect 243228 46872 243268 46900
rect 243228 46860 243234 46872
rect 243262 46860 243268 46872
rect 243320 46860 243326 46912
rect 266998 46860 267004 46912
rect 267056 46900 267062 46912
rect 267182 46900 267188 46912
rect 267056 46872 267188 46900
rect 267056 46860 267062 46872
rect 267182 46860 267188 46872
rect 267240 46860 267246 46912
rect 282914 46860 282920 46912
rect 282972 46900 282978 46912
rect 283098 46900 283104 46912
rect 282972 46872 283104 46900
rect 282972 46860 282978 46872
rect 283098 46860 283104 46872
rect 283156 46860 283162 46912
rect 310517 46903 310575 46909
rect 310517 46869 310529 46903
rect 310563 46900 310575 46903
rect 310606 46900 310612 46912
rect 310563 46872 310612 46900
rect 310563 46869 310575 46872
rect 310517 46863 310575 46869
rect 310606 46860 310612 46872
rect 310664 46860 310670 46912
rect 332888 46844 332916 46928
rect 342438 46900 342444 46912
rect 342399 46872 342444 46900
rect 342438 46860 342444 46872
rect 342496 46860 342502 46912
rect 358998 46860 359004 46912
rect 359056 46900 359062 46912
rect 359182 46900 359188 46912
rect 359056 46872 359188 46900
rect 359056 46860 359062 46872
rect 359182 46860 359188 46872
rect 359240 46860 359246 46912
rect 371326 46860 371332 46912
rect 371384 46860 371390 46912
rect 387886 46900 387892 46912
rect 387847 46872 387892 46900
rect 387886 46860 387892 46872
rect 387944 46860 387950 46912
rect 392118 46860 392124 46912
rect 392176 46860 392182 46912
rect 408770 46900 408776 46912
rect 408731 46872 408776 46900
rect 408770 46860 408776 46872
rect 408828 46860 408834 46912
rect 332870 46792 332876 46844
rect 332928 46792 332934 46844
rect 371344 46832 371372 46860
rect 371510 46832 371516 46844
rect 371344 46804 371516 46832
rect 371510 46792 371516 46804
rect 371568 46792 371574 46844
rect 392136 46776 392164 46860
rect 392118 46724 392124 46776
rect 392176 46724 392182 46776
rect 271969 45611 272027 45617
rect 271969 45577 271981 45611
rect 272015 45608 272027 45611
rect 272058 45608 272064 45620
rect 272015 45580 272064 45608
rect 272015 45577 272027 45580
rect 271969 45571 272027 45577
rect 272058 45568 272064 45580
rect 272116 45568 272122 45620
rect 292761 45611 292819 45617
rect 292761 45577 292773 45611
rect 292807 45608 292819 45611
rect 292942 45608 292948 45620
rect 292807 45580 292948 45608
rect 292807 45577 292819 45580
rect 292761 45571 292819 45577
rect 292942 45568 292948 45580
rect 293000 45568 293006 45620
rect 324498 45608 324504 45620
rect 324459 45580 324504 45608
rect 324498 45568 324504 45580
rect 324556 45568 324562 45620
rect 242989 45543 243047 45549
rect 242989 45509 243001 45543
rect 243035 45540 243047 45543
rect 243262 45540 243268 45552
rect 243035 45512 243268 45540
rect 243035 45509 243047 45512
rect 242989 45503 243047 45509
rect 243262 45500 243268 45512
rect 243320 45500 243326 45552
rect 267001 45543 267059 45549
rect 267001 45509 267013 45543
rect 267047 45540 267059 45543
rect 267182 45540 267188 45552
rect 267047 45512 267188 45540
rect 267047 45509 267059 45512
rect 267001 45503 267059 45509
rect 267182 45500 267188 45512
rect 267240 45500 267246 45552
rect 277578 45540 277584 45552
rect 277539 45512 277584 45540
rect 277578 45500 277584 45512
rect 277636 45500 277642 45552
rect 282917 45543 282975 45549
rect 282917 45509 282929 45543
rect 282963 45540 282975 45543
rect 283098 45540 283104 45552
rect 282963 45512 283104 45540
rect 282963 45509 282975 45512
rect 282917 45503 282975 45509
rect 283098 45500 283104 45512
rect 283156 45500 283162 45552
rect 332689 45543 332747 45549
rect 332689 45509 332701 45543
rect 332735 45540 332747 45543
rect 332870 45540 332876 45552
rect 332735 45512 332876 45540
rect 332735 45509 332747 45512
rect 332689 45503 332747 45509
rect 332870 45500 332876 45512
rect 332928 45500 332934 45552
rect 352006 45500 352012 45552
rect 352064 45540 352070 45552
rect 352374 45540 352380 45552
rect 352064 45512 352380 45540
rect 352064 45500 352070 45512
rect 352374 45500 352380 45512
rect 352432 45500 352438 45552
rect 358998 45540 359004 45552
rect 358959 45512 359004 45540
rect 358998 45500 359004 45512
rect 359056 45500 359062 45552
rect 255406 44820 255412 44872
rect 255464 44860 255470 44872
rect 255501 44863 255559 44869
rect 255501 44860 255513 44863
rect 255464 44832 255513 44860
rect 255464 44820 255470 44832
rect 255501 44829 255513 44832
rect 255547 44829 255559 44863
rect 255501 44823 255559 44829
rect 230658 43460 230664 43512
rect 230716 43500 230722 43512
rect 230842 43500 230848 43512
rect 230716 43472 230848 43500
rect 230716 43460 230722 43472
rect 230842 43460 230848 43472
rect 230900 43460 230906 43512
rect 298370 42072 298376 42084
rect 298331 42044 298376 42072
rect 298370 42032 298376 42044
rect 298428 42032 298434 42084
rect 309321 42075 309379 42081
rect 309321 42041 309333 42075
rect 309367 42072 309379 42075
rect 309410 42072 309416 42084
rect 309367 42044 309416 42072
rect 309367 42041 309379 42044
rect 309321 42035 309379 42041
rect 309410 42032 309416 42044
rect 309468 42032 309474 42084
rect 375469 41599 375527 41605
rect 375469 41565 375481 41599
rect 375515 41596 375527 41599
rect 375650 41596 375656 41608
rect 375515 41568 375656 41596
rect 375515 41565 375527 41568
rect 375469 41559 375527 41565
rect 375650 41556 375656 41568
rect 375708 41556 375714 41608
rect 369949 41463 370007 41469
rect 369949 41429 369961 41463
rect 369995 41460 370007 41463
rect 370130 41460 370136 41472
rect 369995 41432 370136 41460
rect 369995 41429 370007 41432
rect 369949 41423 370007 41429
rect 370130 41420 370136 41432
rect 370188 41420 370194 41472
rect 310517 41395 310575 41401
rect 310517 41361 310529 41395
rect 310563 41392 310575 41395
rect 310606 41392 310612 41404
rect 310563 41364 310612 41392
rect 310563 41361 310575 41364
rect 310517 41355 310575 41361
rect 310606 41352 310612 41364
rect 310664 41352 310670 41404
rect 471974 41352 471980 41404
rect 472032 41392 472038 41404
rect 472158 41392 472164 41404
rect 472032 41364 472164 41392
rect 472032 41352 472038 41364
rect 472158 41352 472164 41364
rect 472216 41352 472222 41404
rect 433610 41324 433616 41336
rect 433571 41296 433616 41324
rect 433610 41284 433616 41296
rect 433668 41284 433674 41336
rect 397638 40332 397644 40384
rect 397696 40372 397702 40384
rect 405642 40372 405648 40384
rect 397696 40344 405648 40372
rect 397696 40332 397702 40344
rect 405642 40332 405648 40344
rect 405700 40332 405706 40384
rect 475930 40196 475936 40248
rect 475988 40236 475994 40248
rect 478230 40236 478236 40248
rect 475988 40208 478236 40236
rect 475988 40196 475994 40208
rect 478230 40196 478236 40208
rect 478288 40196 478294 40248
rect 514570 40196 514576 40248
rect 514628 40236 514634 40248
rect 514846 40236 514852 40248
rect 514628 40208 514852 40236
rect 514628 40196 514634 40208
rect 514846 40196 514852 40208
rect 514904 40196 514910 40248
rect 540974 40060 540980 40112
rect 541032 40100 541038 40112
rect 545850 40100 545856 40112
rect 541032 40072 545856 40100
rect 541032 40060 541038 40072
rect 545850 40060 545856 40072
rect 545908 40060 545914 40112
rect 302142 39992 302148 40044
rect 302200 40032 302206 40044
rect 307294 40032 307300 40044
rect 302200 40004 307300 40032
rect 302200 39992 302206 40004
rect 307294 39992 307300 40004
rect 307352 39992 307358 40044
rect 272058 38740 272064 38752
rect 272019 38712 272064 38740
rect 272058 38700 272064 38712
rect 272116 38700 272122 38752
rect 382366 38700 382372 38752
rect 382424 38700 382430 38752
rect 281626 38632 281632 38684
rect 281684 38672 281690 38684
rect 281810 38672 281816 38684
rect 281684 38644 281816 38672
rect 281684 38632 281690 38644
rect 281810 38632 281816 38644
rect 281868 38632 281874 38684
rect 308122 38672 308128 38684
rect 308083 38644 308128 38672
rect 308122 38632 308128 38644
rect 308180 38632 308186 38684
rect 376938 38632 376944 38684
rect 376996 38672 377002 38684
rect 377030 38672 377036 38684
rect 376996 38644 377036 38672
rect 376996 38632 377002 38644
rect 377030 38632 377036 38644
rect 377088 38632 377094 38684
rect 382384 38616 382412 38700
rect 294138 38604 294144 38616
rect 294099 38576 294144 38604
rect 294138 38564 294144 38576
rect 294196 38564 294202 38616
rect 369946 38604 369952 38616
rect 369907 38576 369952 38604
rect 369946 38564 369952 38576
rect 370004 38564 370010 38616
rect 382366 38564 382372 38616
rect 382424 38564 382430 38616
rect 416869 38607 416927 38613
rect 416869 38573 416881 38607
rect 416915 38604 416927 38607
rect 416958 38604 416964 38616
rect 416915 38576 416964 38604
rect 416915 38573 416927 38576
rect 416869 38567 416927 38573
rect 416958 38564 416964 38576
rect 417016 38564 417022 38616
rect 422478 38604 422484 38616
rect 422439 38576 422484 38604
rect 422478 38564 422484 38576
rect 422536 38564 422542 38616
rect 472069 38607 472127 38613
rect 472069 38573 472081 38607
rect 472115 38604 472127 38607
rect 472158 38604 472164 38616
rect 472115 38576 472164 38604
rect 472115 38573 472127 38576
rect 472069 38567 472127 38573
rect 472158 38564 472164 38576
rect 472216 38564 472222 38616
rect 408773 38539 408831 38545
rect 408773 38505 408785 38539
rect 408819 38536 408831 38539
rect 408862 38536 408868 38548
rect 408819 38508 408868 38536
rect 408819 38505 408831 38508
rect 408773 38499 408831 38505
rect 408862 38496 408868 38508
rect 408920 38496 408926 38548
rect 295702 38292 295708 38344
rect 295760 38292 295766 38344
rect 295720 38208 295748 38292
rect 295702 38156 295708 38208
rect 295760 38156 295766 38208
rect 252738 37380 252744 37392
rect 252699 37352 252744 37380
rect 252738 37340 252744 37352
rect 252796 37340 252802 37392
rect 331490 37380 331496 37392
rect 331416 37352 331496 37380
rect 331416 37324 331444 37352
rect 331490 37340 331496 37352
rect 331548 37340 331554 37392
rect 334434 37380 334440 37392
rect 334360 37352 334440 37380
rect 334360 37324 334388 37352
rect 334434 37340 334440 37352
rect 334492 37340 334498 37392
rect 386690 37340 386696 37392
rect 386748 37340 386754 37392
rect 433518 37340 433524 37392
rect 433576 37380 433582 37392
rect 433613 37383 433671 37389
rect 433613 37380 433625 37383
rect 433576 37352 433625 37380
rect 433576 37340 433582 37352
rect 433613 37349 433625 37352
rect 433659 37349 433671 37383
rect 433613 37343 433671 37349
rect 331398 37272 331404 37324
rect 331456 37272 331462 37324
rect 334342 37272 334348 37324
rect 334400 37272 334406 37324
rect 342441 37315 342499 37321
rect 342441 37281 342453 37315
rect 342487 37312 342499 37315
rect 342530 37312 342536 37324
rect 342487 37284 342536 37312
rect 342487 37281 342499 37284
rect 342441 37275 342499 37281
rect 342530 37272 342536 37284
rect 342588 37272 342594 37324
rect 375466 37312 375472 37324
rect 375427 37284 375472 37312
rect 375466 37272 375472 37284
rect 375524 37272 375530 37324
rect 386708 37312 386736 37340
rect 386782 37312 386788 37324
rect 386708 37284 386788 37312
rect 386782 37272 386788 37284
rect 386840 37272 386846 37324
rect 387886 37312 387892 37324
rect 387847 37284 387892 37312
rect 387886 37272 387892 37284
rect 387944 37272 387950 37324
rect 230658 37204 230664 37256
rect 230716 37244 230722 37256
rect 230750 37244 230756 37256
rect 230716 37216 230756 37244
rect 230716 37204 230722 37216
rect 230750 37204 230756 37216
rect 230808 37204 230814 37256
rect 272058 37244 272064 37256
rect 272019 37216 272064 37244
rect 272058 37204 272064 37216
rect 272116 37204 272122 37256
rect 433610 37244 433616 37256
rect 433571 37216 433616 37244
rect 433610 37204 433616 37216
rect 433668 37204 433674 37256
rect 292761 37179 292819 37185
rect 292761 37145 292773 37179
rect 292807 37176 292819 37179
rect 292942 37176 292948 37188
rect 292807 37148 292948 37176
rect 292807 37145 292819 37148
rect 292761 37139 292819 37145
rect 292942 37136 292948 37148
rect 293000 37136 293006 37188
rect 242986 35952 242992 35964
rect 242947 35924 242992 35952
rect 242986 35912 242992 35924
rect 243044 35912 243050 35964
rect 266998 35952 267004 35964
rect 266959 35924 267004 35952
rect 266998 35912 267004 35924
rect 267056 35912 267062 35964
rect 277578 35952 277584 35964
rect 277539 35924 277584 35952
rect 277578 35912 277584 35924
rect 277636 35912 277642 35964
rect 292758 35952 292764 35964
rect 292719 35924 292764 35952
rect 292758 35912 292764 35924
rect 292816 35912 292822 35964
rect 332686 35952 332692 35964
rect 332647 35924 332692 35952
rect 332686 35912 332692 35924
rect 332744 35912 332750 35964
rect 358998 35952 359004 35964
rect 358959 35924 359004 35952
rect 358998 35912 359004 35924
rect 359056 35912 359062 35964
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 72418 35884 72424 35896
rect 3476 35856 72424 35884
rect 3476 35844 3482 35856
rect 72418 35844 72424 35856
rect 72476 35844 72482 35896
rect 334342 35884 334348 35896
rect 334303 35856 334348 35884
rect 334342 35844 334348 35856
rect 334400 35844 334406 35896
rect 369946 33804 369952 33856
rect 370004 33844 370010 33856
rect 370222 33844 370228 33856
rect 370004 33816 370228 33844
rect 370004 33804 370010 33816
rect 370222 33804 370228 33816
rect 370280 33804 370286 33856
rect 298186 32376 298192 32428
rect 298244 32416 298250 32428
rect 298373 32419 298431 32425
rect 298373 32416 298385 32419
rect 298244 32388 298385 32416
rect 298244 32376 298250 32388
rect 298373 32385 298385 32388
rect 298419 32385 298431 32419
rect 298373 32379 298431 32385
rect 319070 31764 319076 31816
rect 319128 31764 319134 31816
rect 346578 31804 346584 31816
rect 346504 31776 346584 31804
rect 233326 31696 233332 31748
rect 233384 31736 233390 31748
rect 233510 31736 233516 31748
rect 233384 31708 233516 31736
rect 233384 31696 233390 31708
rect 233510 31696 233516 31708
rect 233568 31696 233574 31748
rect 281626 31696 281632 31748
rect 281684 31736 281690 31748
rect 281810 31736 281816 31748
rect 281684 31708 281816 31736
rect 281684 31696 281690 31708
rect 281810 31696 281816 31708
rect 281868 31696 281874 31748
rect 319088 31680 319116 31764
rect 346504 31748 346532 31776
rect 346578 31764 346584 31776
rect 346636 31764 346642 31816
rect 400674 31804 400680 31816
rect 400635 31776 400680 31804
rect 400674 31764 400680 31776
rect 400732 31764 400738 31816
rect 427906 31804 427912 31816
rect 427832 31776 427912 31804
rect 427832 31748 427860 31776
rect 427906 31764 427912 31776
rect 427964 31764 427970 31816
rect 346486 31696 346492 31748
rect 346544 31696 346550 31748
rect 427814 31696 427820 31748
rect 427872 31696 427878 31748
rect 451642 31696 451648 31748
rect 451700 31736 451706 31748
rect 451826 31736 451832 31748
rect 451700 31708 451832 31736
rect 451700 31696 451706 31708
rect 451826 31696 451832 31708
rect 451884 31696 451890 31748
rect 319070 31628 319076 31680
rect 319128 31628 319134 31680
rect 270678 29044 270684 29096
rect 270736 29044 270742 29096
rect 294138 29084 294144 29096
rect 294099 29056 294144 29084
rect 294138 29044 294144 29056
rect 294196 29044 294202 29096
rect 400674 29084 400680 29096
rect 400635 29056 400680 29084
rect 400674 29044 400680 29056
rect 400732 29044 400738 29096
rect 236270 28976 236276 29028
rect 236328 29016 236334 29028
rect 236362 29016 236368 29028
rect 236328 28988 236368 29016
rect 236328 28976 236334 28988
rect 236362 28976 236368 28988
rect 236420 28976 236426 29028
rect 252741 29019 252799 29025
rect 252741 28985 252753 29019
rect 252787 29016 252799 29019
rect 252830 29016 252836 29028
rect 252787 28988 252836 29016
rect 252787 28985 252799 28988
rect 252741 28979 252799 28985
rect 252830 28976 252836 28988
rect 252888 28976 252894 29028
rect 270696 29016 270724 29044
rect 270770 29016 270776 29028
rect 270696 28988 270776 29016
rect 270770 28976 270776 28988
rect 270828 28976 270834 29028
rect 309318 29016 309324 29028
rect 309279 28988 309324 29016
rect 309318 28976 309324 28988
rect 309376 28976 309382 29028
rect 381170 28976 381176 29028
rect 381228 29016 381234 29028
rect 381262 29016 381268 29028
rect 381228 28988 381268 29016
rect 381228 28976 381234 28988
rect 381262 28976 381268 28988
rect 381320 28976 381326 29028
rect 386690 28976 386696 29028
rect 386748 29016 386754 29028
rect 416866 29016 416872 29028
rect 386748 28988 386828 29016
rect 416827 28988 416872 29016
rect 386748 28976 386754 28988
rect 231854 28908 231860 28960
rect 231912 28948 231918 28960
rect 232038 28948 232044 28960
rect 231912 28920 232044 28948
rect 231912 28908 231918 28920
rect 232038 28908 232044 28920
rect 232096 28908 232102 28960
rect 244458 28908 244464 28960
rect 244516 28948 244522 28960
rect 244550 28948 244556 28960
rect 244516 28920 244556 28948
rect 244516 28908 244522 28920
rect 244550 28908 244556 28920
rect 244608 28908 244614 28960
rect 254026 28908 254032 28960
rect 254084 28948 254090 28960
rect 254210 28948 254216 28960
rect 254084 28920 254216 28948
rect 254084 28908 254090 28920
rect 254210 28908 254216 28920
rect 254268 28908 254274 28960
rect 259730 28908 259736 28960
rect 259788 28948 259794 28960
rect 259822 28948 259828 28960
rect 259788 28920 259828 28948
rect 259788 28908 259794 28920
rect 259822 28908 259828 28920
rect 259880 28908 259886 28960
rect 265158 28908 265164 28960
rect 265216 28948 265222 28960
rect 265250 28948 265256 28960
rect 265216 28920 265256 28948
rect 265216 28908 265222 28920
rect 265250 28908 265256 28920
rect 265308 28908 265314 28960
rect 266354 28908 266360 28960
rect 266412 28948 266418 28960
rect 266538 28948 266544 28960
rect 266412 28920 266544 28948
rect 266412 28908 266418 28920
rect 266538 28908 266544 28920
rect 266596 28908 266602 28960
rect 292758 28908 292764 28960
rect 292816 28948 292822 28960
rect 292850 28948 292856 28960
rect 292816 28920 292856 28948
rect 292816 28908 292822 28920
rect 292850 28908 292856 28920
rect 292908 28908 292914 28960
rect 293954 28908 293960 28960
rect 294012 28948 294018 28960
rect 294138 28948 294144 28960
rect 294012 28920 294144 28948
rect 294012 28908 294018 28920
rect 294138 28908 294144 28920
rect 294196 28908 294202 28960
rect 295518 28908 295524 28960
rect 295576 28948 295582 28960
rect 295610 28948 295616 28960
rect 295576 28920 295616 28948
rect 295576 28908 295582 28920
rect 295610 28908 295616 28920
rect 295668 28908 295674 28960
rect 308033 28951 308091 28957
rect 308033 28917 308045 28951
rect 308079 28948 308091 28951
rect 308122 28948 308128 28960
rect 308079 28920 308128 28948
rect 308079 28917 308091 28920
rect 308033 28911 308091 28917
rect 308122 28908 308128 28920
rect 308180 28908 308186 28960
rect 348050 28908 348056 28960
rect 348108 28948 348114 28960
rect 348142 28948 348148 28960
rect 348108 28920 348148 28948
rect 348108 28908 348114 28920
rect 348142 28908 348148 28920
rect 348200 28908 348206 28960
rect 353570 28908 353576 28960
rect 353628 28948 353634 28960
rect 353662 28948 353668 28960
rect 353628 28920 353668 28948
rect 353628 28908 353634 28920
rect 353662 28908 353668 28920
rect 353720 28908 353726 28960
rect 356422 28908 356428 28960
rect 356480 28948 356486 28960
rect 356514 28948 356520 28960
rect 356480 28920 356520 28948
rect 356480 28908 356486 28920
rect 356514 28908 356520 28920
rect 356572 28908 356578 28960
rect 386800 28892 386828 28988
rect 416866 28976 416872 28988
rect 416924 28976 416930 29028
rect 466546 28976 466552 29028
rect 466604 29016 466610 29028
rect 466638 29016 466644 29028
rect 466604 28988 466644 29016
rect 466604 28976 466610 28988
rect 466638 28976 466644 28988
rect 466696 28976 466702 29028
rect 472066 29016 472072 29028
rect 472027 28988 472072 29016
rect 472066 28976 472072 28988
rect 472124 28976 472130 29028
rect 392026 28908 392032 28960
rect 392084 28948 392090 28960
rect 392210 28948 392216 28960
rect 392084 28920 392216 28948
rect 392084 28908 392090 28920
rect 392210 28908 392216 28920
rect 392268 28908 392274 28960
rect 393222 28948 393228 28960
rect 393183 28920 393228 28948
rect 393222 28908 393228 28920
rect 393280 28908 393286 28960
rect 451737 28951 451795 28957
rect 451737 28917 451749 28951
rect 451783 28948 451795 28951
rect 451826 28948 451832 28960
rect 451783 28920 451832 28948
rect 451783 28917 451795 28920
rect 451737 28911 451795 28917
rect 451826 28908 451832 28920
rect 451884 28908 451890 28960
rect 386782 28840 386788 28892
rect 386840 28840 386846 28892
rect 387797 27795 387855 27801
rect 387797 27761 387809 27795
rect 387843 27792 387855 27795
rect 387886 27792 387892 27804
rect 387843 27764 387892 27792
rect 387843 27761 387855 27764
rect 387797 27755 387855 27761
rect 387886 27752 387892 27764
rect 387944 27752 387950 27804
rect 277578 27684 277584 27736
rect 277636 27724 277642 27736
rect 277670 27724 277676 27736
rect 277636 27696 277676 27724
rect 277636 27684 277642 27696
rect 277670 27684 277676 27696
rect 277728 27684 277734 27736
rect 282914 27656 282920 27668
rect 282875 27628 282920 27656
rect 282914 27616 282920 27628
rect 282972 27616 282978 27668
rect 327166 27616 327172 27668
rect 327224 27656 327230 27668
rect 327258 27656 327264 27668
rect 327224 27628 327264 27656
rect 327224 27616 327230 27628
rect 327258 27616 327264 27628
rect 327316 27616 327322 27668
rect 387794 27656 387800 27668
rect 387755 27628 387800 27656
rect 387794 27616 387800 27628
rect 387852 27616 387858 27668
rect 422386 27616 422392 27668
rect 422444 27656 422450 27668
rect 422481 27659 422539 27665
rect 422481 27656 422493 27659
rect 422444 27628 422493 27656
rect 422444 27616 422450 27628
rect 422481 27625 422493 27628
rect 422527 27625 422539 27659
rect 422481 27619 422539 27625
rect 433613 27659 433671 27665
rect 433613 27625 433625 27659
rect 433659 27656 433671 27659
rect 433702 27656 433708 27668
rect 433659 27628 433708 27656
rect 433659 27625 433671 27628
rect 433613 27619 433671 27625
rect 433702 27616 433708 27628
rect 433760 27616 433766 27668
rect 230750 27548 230756 27600
rect 230808 27588 230814 27600
rect 230842 27588 230848 27600
rect 230808 27560 230848 27588
rect 230808 27548 230814 27560
rect 230842 27548 230848 27560
rect 230900 27548 230906 27600
rect 252830 27588 252836 27600
rect 252791 27560 252836 27588
rect 252830 27548 252836 27560
rect 252888 27548 252894 27600
rect 255314 27548 255320 27600
rect 255372 27588 255378 27600
rect 255501 27591 255559 27597
rect 255501 27588 255513 27591
rect 255372 27560 255513 27588
rect 255372 27548 255378 27560
rect 255501 27557 255513 27560
rect 255547 27557 255559 27591
rect 259822 27588 259828 27600
rect 259783 27560 259828 27588
rect 255501 27551 255559 27557
rect 259822 27548 259828 27560
rect 259880 27548 259886 27600
rect 266998 27548 267004 27600
rect 267056 27588 267062 27600
rect 267090 27588 267096 27600
rect 267056 27560 267096 27588
rect 267056 27548 267062 27560
rect 267090 27548 267096 27560
rect 267148 27548 267154 27600
rect 271969 27591 272027 27597
rect 271969 27557 271981 27591
rect 272015 27588 272027 27591
rect 272058 27588 272064 27600
rect 272015 27560 272064 27588
rect 272015 27557 272027 27560
rect 271969 27551 272027 27557
rect 272058 27548 272064 27560
rect 272116 27548 272122 27600
rect 293954 27588 293960 27600
rect 293915 27560 293960 27588
rect 293954 27548 293960 27560
rect 294012 27548 294018 27600
rect 321646 27588 321652 27600
rect 321607 27560 321652 27588
rect 321646 27548 321652 27560
rect 321704 27548 321710 27600
rect 336829 27591 336887 27597
rect 336829 27557 336841 27591
rect 336875 27588 336887 27591
rect 336918 27588 336924 27600
rect 336875 27560 336924 27588
rect 336875 27557 336887 27560
rect 336829 27551 336887 27557
rect 336918 27548 336924 27560
rect 336976 27548 336982 27600
rect 346397 27591 346455 27597
rect 346397 27557 346409 27591
rect 346443 27588 346455 27591
rect 346486 27588 346492 27600
rect 346443 27560 346492 27588
rect 346443 27557 346455 27560
rect 346397 27551 346455 27557
rect 346486 27548 346492 27560
rect 346544 27548 346550 27600
rect 353662 27588 353668 27600
rect 353623 27560 353668 27588
rect 353662 27548 353668 27560
rect 353720 27548 353726 27600
rect 358998 27588 359004 27600
rect 358959 27560 359004 27588
rect 358998 27548 359004 27560
rect 359056 27548 359062 27600
rect 400582 27588 400588 27600
rect 400543 27560 400588 27588
rect 400582 27548 400588 27560
rect 400640 27548 400646 27600
rect 324498 26364 324504 26376
rect 324424 26336 324504 26364
rect 324424 26308 324452 26336
rect 324498 26324 324504 26336
rect 324556 26324 324562 26376
rect 324406 26256 324412 26308
rect 324464 26256 324470 26308
rect 334345 26299 334403 26305
rect 334345 26265 334357 26299
rect 334391 26296 334403 26299
rect 334526 26296 334532 26308
rect 334391 26268 334532 26296
rect 334391 26265 334403 26268
rect 334345 26259 334403 26265
rect 334526 26256 334532 26268
rect 334584 26256 334590 26308
rect 230661 26231 230719 26237
rect 230661 26197 230673 26231
rect 230707 26228 230719 26231
rect 230750 26228 230756 26240
rect 230707 26200 230756 26228
rect 230707 26197 230719 26200
rect 230661 26191 230719 26197
rect 230750 26188 230756 26200
rect 230808 26188 230814 26240
rect 277489 26231 277547 26237
rect 277489 26197 277501 26231
rect 277535 26228 277547 26231
rect 277578 26228 277584 26240
rect 277535 26200 277584 26228
rect 277535 26197 277547 26200
rect 277489 26191 277547 26197
rect 277578 26188 277584 26200
rect 277636 26188 277642 26240
rect 334342 26120 334348 26172
rect 334400 26160 334406 26172
rect 334526 26160 334532 26172
rect 334400 26132 334532 26160
rect 334400 26120 334406 26132
rect 334526 26120 334532 26132
rect 334584 26120 334590 26172
rect 346397 22763 346455 22769
rect 346397 22729 346409 22763
rect 346443 22760 346455 22763
rect 346486 22760 346492 22772
rect 346443 22732 346492 22760
rect 346443 22729 346455 22732
rect 346397 22723 346455 22729
rect 346486 22720 346492 22732
rect 346544 22720 346550 22772
rect 347869 22763 347927 22769
rect 347869 22729 347881 22763
rect 347915 22760 347927 22763
rect 348142 22760 348148 22772
rect 347915 22732 348148 22760
rect 347915 22729 347927 22732
rect 347869 22723 347927 22729
rect 348142 22720 348148 22732
rect 348200 22720 348206 22772
rect 270681 22627 270739 22633
rect 270681 22593 270693 22627
rect 270727 22624 270739 22627
rect 270770 22624 270776 22636
rect 270727 22596 270776 22624
rect 270727 22593 270739 22596
rect 270681 22587 270739 22593
rect 270770 22584 270776 22596
rect 270828 22584 270834 22636
rect 305089 22219 305147 22225
rect 305089 22185 305101 22219
rect 305135 22216 305147 22219
rect 305270 22216 305276 22228
rect 305135 22188 305276 22216
rect 305135 22185 305147 22188
rect 305089 22179 305147 22185
rect 305270 22176 305276 22188
rect 305328 22176 305334 22228
rect 281810 22148 281816 22160
rect 281736 22120 281816 22148
rect 281736 22092 281764 22120
rect 281810 22108 281816 22120
rect 281868 22108 281874 22160
rect 364518 22108 364524 22160
rect 364576 22108 364582 22160
rect 408770 22148 408776 22160
rect 408696 22120 408776 22148
rect 281718 22040 281724 22092
rect 281776 22040 281782 22092
rect 364536 22024 364564 22108
rect 408696 22092 408724 22120
rect 408770 22108 408776 22120
rect 408828 22108 408834 22160
rect 408678 22040 408684 22092
rect 408736 22040 408742 22092
rect 416774 22040 416780 22092
rect 416832 22080 416838 22092
rect 416958 22080 416964 22092
rect 416832 22052 416964 22080
rect 416832 22040 416838 22052
rect 416958 22040 416964 22052
rect 417016 22040 417022 22092
rect 364518 21972 364524 22024
rect 364576 21972 364582 22024
rect 236270 19320 236276 19372
rect 236328 19320 236334 19372
rect 260926 19320 260932 19372
rect 260984 19360 260990 19372
rect 261018 19360 261024 19372
rect 260984 19332 261024 19360
rect 260984 19320 260990 19332
rect 261018 19320 261024 19332
rect 261076 19320 261082 19372
rect 282914 19320 282920 19372
rect 282972 19360 282978 19372
rect 283190 19360 283196 19372
rect 282972 19332 283196 19360
rect 282972 19320 282978 19332
rect 283190 19320 283196 19332
rect 283248 19320 283254 19372
rect 288434 19320 288440 19372
rect 288492 19360 288498 19372
rect 288618 19360 288624 19372
rect 288492 19332 288624 19360
rect 288492 19320 288498 19332
rect 288618 19320 288624 19332
rect 288676 19320 288682 19372
rect 305086 19360 305092 19372
rect 305047 19332 305092 19360
rect 305086 19320 305092 19332
rect 305144 19320 305150 19372
rect 308030 19360 308036 19372
rect 307991 19332 308036 19360
rect 308030 19320 308036 19332
rect 308088 19320 308094 19372
rect 310422 19320 310428 19372
rect 310480 19360 310486 19372
rect 310698 19360 310704 19372
rect 310480 19332 310704 19360
rect 310480 19320 310486 19332
rect 310698 19320 310704 19332
rect 310756 19320 310762 19372
rect 324406 19320 324412 19372
rect 324464 19360 324470 19372
rect 324498 19360 324504 19372
rect 324464 19332 324504 19360
rect 324464 19320 324470 19332
rect 324498 19320 324504 19332
rect 324556 19320 324562 19372
rect 352006 19320 352012 19372
rect 352064 19360 352070 19372
rect 352190 19360 352196 19372
rect 352064 19332 352196 19360
rect 352064 19320 352070 19332
rect 352190 19320 352196 19332
rect 352248 19320 352254 19372
rect 357526 19320 357532 19372
rect 357584 19360 357590 19372
rect 357618 19360 357624 19372
rect 357584 19332 357624 19360
rect 357584 19320 357590 19332
rect 357618 19320 357624 19332
rect 357676 19320 357682 19372
rect 370038 19320 370044 19372
rect 370096 19360 370102 19372
rect 370222 19360 370228 19372
rect 370096 19332 370228 19360
rect 370096 19320 370102 19332
rect 370222 19320 370228 19332
rect 370280 19320 370286 19372
rect 371326 19320 371332 19372
rect 371384 19360 371390 19372
rect 371510 19360 371516 19372
rect 371384 19332 371516 19360
rect 371384 19320 371390 19332
rect 371510 19320 371516 19332
rect 371568 19320 371574 19372
rect 375558 19320 375564 19372
rect 375616 19360 375622 19372
rect 375742 19360 375748 19372
rect 375616 19332 375748 19360
rect 375616 19320 375622 19332
rect 375742 19320 375748 19332
rect 375800 19320 375806 19372
rect 381078 19320 381084 19372
rect 381136 19360 381142 19372
rect 381262 19360 381268 19372
rect 381136 19332 381268 19360
rect 381136 19320 381142 19332
rect 381262 19320 381268 19332
rect 381320 19320 381326 19372
rect 382274 19320 382280 19372
rect 382332 19360 382338 19372
rect 382458 19360 382464 19372
rect 382332 19332 382464 19360
rect 382332 19320 382338 19332
rect 382458 19320 382464 19332
rect 382516 19320 382522 19372
rect 393222 19360 393228 19372
rect 393183 19332 393228 19360
rect 393222 19320 393228 19332
rect 393280 19320 393286 19372
rect 451734 19360 451740 19372
rect 451695 19332 451740 19360
rect 451734 19320 451740 19332
rect 451792 19320 451798 19372
rect 231854 19252 231860 19304
rect 231912 19252 231918 19304
rect 233326 19252 233332 19304
rect 233384 19292 233390 19304
rect 233418 19292 233424 19304
rect 233384 19264 233424 19292
rect 233384 19252 233390 19264
rect 233418 19252 233424 19264
rect 233476 19252 233482 19304
rect 231872 19224 231900 19252
rect 231946 19224 231952 19236
rect 231872 19196 231952 19224
rect 231946 19184 231952 19196
rect 232004 19184 232010 19236
rect 236288 19224 236316 19320
rect 353662 19292 353668 19304
rect 353623 19264 353668 19292
rect 353662 19252 353668 19264
rect 353720 19252 353726 19304
rect 416958 19292 416964 19304
rect 416919 19264 416964 19292
rect 416958 19252 416964 19264
rect 417016 19252 417022 19304
rect 236362 19224 236368 19236
rect 236288 19196 236368 19224
rect 236362 19184 236368 19196
rect 236420 19184 236426 19236
rect 422110 19184 422116 19236
rect 422168 19224 422174 19236
rect 422478 19224 422484 19236
rect 422168 19196 422484 19224
rect 422168 19184 422174 19196
rect 422478 19184 422484 19196
rect 422536 19184 422542 19236
rect 386782 18980 386788 19032
rect 386840 18980 386846 19032
rect 386800 18896 386828 18980
rect 386782 18844 386788 18896
rect 386840 18844 386846 18896
rect 252830 18000 252836 18012
rect 252791 17972 252836 18000
rect 252830 17960 252836 17972
rect 252888 17960 252894 18012
rect 259822 18000 259828 18012
rect 259783 17972 259828 18000
rect 259822 17960 259828 17972
rect 259880 17960 259886 18012
rect 271966 18000 271972 18012
rect 271927 17972 271972 18000
rect 271966 17960 271972 17972
rect 272024 17960 272030 18012
rect 293954 18000 293960 18012
rect 293915 17972 293960 18000
rect 293954 17960 293960 17972
rect 294012 17960 294018 18012
rect 321649 18003 321707 18009
rect 321649 17969 321661 18003
rect 321695 18000 321707 18003
rect 321738 18000 321744 18012
rect 321695 17972 321744 18000
rect 321695 17969 321707 17972
rect 321649 17963 321707 17969
rect 321738 17960 321744 17972
rect 321796 17960 321802 18012
rect 336826 18000 336832 18012
rect 336787 17972 336832 18000
rect 336826 17960 336832 17972
rect 336884 17960 336890 18012
rect 358998 18000 359004 18012
rect 358959 17972 359004 18000
rect 358998 17960 359004 17972
rect 359056 17960 359062 18012
rect 400582 18000 400588 18012
rect 400543 17972 400588 18000
rect 400582 17960 400588 17972
rect 400640 17960 400646 18012
rect 380989 17935 381047 17941
rect 380989 17901 381001 17935
rect 381035 17932 381047 17935
rect 381078 17932 381084 17944
rect 381035 17904 381084 17932
rect 381035 17901 381047 17904
rect 380989 17895 381047 17901
rect 381078 17892 381084 17904
rect 381136 17892 381142 17944
rect 382369 17935 382427 17941
rect 382369 17901 382381 17935
rect 382415 17932 382427 17935
rect 382458 17932 382464 17944
rect 382415 17904 382464 17932
rect 382415 17901 382427 17904
rect 382369 17895 382427 17901
rect 382458 17892 382464 17904
rect 382516 17892 382522 17944
rect 400401 17867 400459 17873
rect 400401 17833 400413 17867
rect 400447 17864 400459 17867
rect 400582 17864 400588 17876
rect 400447 17836 400588 17864
rect 400447 17833 400459 17836
rect 400401 17827 400459 17833
rect 400582 17824 400588 17836
rect 400640 17824 400646 17876
rect 278774 16872 278780 16924
rect 278832 16912 278838 16924
rect 288342 16912 288348 16924
rect 278832 16884 288348 16912
rect 278832 16872 278838 16884
rect 288342 16872 288348 16884
rect 288400 16872 288406 16924
rect 408402 16804 408408 16856
rect 408460 16844 408466 16856
rect 410702 16844 410708 16856
rect 408460 16816 410708 16844
rect 408460 16804 408466 16816
rect 410702 16804 410708 16816
rect 410760 16804 410766 16856
rect 475930 16804 475936 16856
rect 475988 16844 475994 16856
rect 477494 16844 477500 16856
rect 475988 16816 477500 16844
rect 475988 16804 475994 16816
rect 477494 16804 477500 16816
rect 477552 16804 477558 16856
rect 347682 16668 347688 16720
rect 347740 16708 347746 16720
rect 355962 16708 355968 16720
rect 347740 16680 355968 16708
rect 347740 16668 347746 16680
rect 355962 16668 355968 16680
rect 356020 16668 356026 16720
rect 521654 16668 521660 16720
rect 521712 16708 521718 16720
rect 524506 16708 524512 16720
rect 521712 16680 524512 16708
rect 521712 16668 521718 16680
rect 524506 16668 524512 16680
rect 524564 16668 524570 16720
rect 277486 16640 277492 16652
rect 277447 16612 277492 16640
rect 277486 16600 277492 16612
rect 277544 16600 277550 16652
rect 125410 16328 125416 16380
rect 125468 16368 125474 16380
rect 292758 16368 292764 16380
rect 125468 16340 292764 16368
rect 125468 16328 125474 16340
rect 292758 16328 292764 16340
rect 292816 16328 292822 16380
rect 121362 16260 121368 16312
rect 121420 16300 121426 16312
rect 291286 16300 291292 16312
rect 121420 16272 291292 16300
rect 121420 16260 121426 16272
rect 291286 16260 291292 16272
rect 291344 16260 291350 16312
rect 114462 16192 114468 16244
rect 114520 16232 114526 16244
rect 287238 16232 287244 16244
rect 114520 16204 287244 16232
rect 114520 16192 114526 16204
rect 287238 16192 287244 16204
rect 287296 16192 287302 16244
rect 110322 16124 110328 16176
rect 110380 16164 110386 16176
rect 285766 16164 285772 16176
rect 110380 16136 285772 16164
rect 110380 16124 110386 16136
rect 285766 16124 285772 16136
rect 285824 16124 285830 16176
rect 107562 16056 107568 16108
rect 107620 16096 107626 16108
rect 284386 16096 284392 16108
rect 107620 16068 284392 16096
rect 107620 16056 107626 16068
rect 284386 16056 284392 16068
rect 284444 16056 284450 16108
rect 103422 15988 103428 16040
rect 103480 16028 103486 16040
rect 281718 16028 281724 16040
rect 103480 16000 281724 16028
rect 103480 15988 103486 16000
rect 281718 15988 281724 16000
rect 281776 15988 281782 16040
rect 28902 15920 28908 15972
rect 28960 15960 28966 15972
rect 243078 15960 243084 15972
rect 28960 15932 243084 15960
rect 28960 15920 28966 15932
rect 243078 15920 243084 15932
rect 243136 15920 243142 15972
rect 31662 15852 31668 15904
rect 31720 15892 31726 15904
rect 245746 15892 245752 15904
rect 31720 15864 245752 15892
rect 31720 15852 31726 15864
rect 245746 15852 245752 15864
rect 245804 15852 245810 15904
rect 129642 15104 129648 15156
rect 129700 15144 129706 15156
rect 295518 15144 295524 15156
rect 129700 15116 295524 15144
rect 129700 15104 129706 15116
rect 295518 15104 295524 15116
rect 295576 15104 295582 15156
rect 99282 15036 99288 15088
rect 99340 15076 99346 15088
rect 280246 15076 280252 15088
rect 99340 15048 280252 15076
rect 99340 15036 99346 15048
rect 280246 15036 280252 15048
rect 280304 15036 280310 15088
rect 96522 14968 96528 15020
rect 96580 15008 96586 15020
rect 278866 15008 278872 15020
rect 96580 14980 278872 15008
rect 96580 14968 96586 14980
rect 278866 14968 278872 14980
rect 278924 14968 278930 15020
rect 92382 14900 92388 14952
rect 92440 14940 92446 14952
rect 276106 14940 276112 14952
rect 92440 14912 276112 14940
rect 92440 14900 92446 14912
rect 276106 14900 276112 14912
rect 276164 14900 276170 14952
rect 89622 14832 89628 14884
rect 89680 14872 89686 14884
rect 274726 14872 274732 14884
rect 89680 14844 274732 14872
rect 89680 14832 89686 14844
rect 274726 14832 274732 14844
rect 274784 14832 274790 14884
rect 85482 14764 85488 14816
rect 85540 14804 85546 14816
rect 273346 14804 273352 14816
rect 85540 14776 273352 14804
rect 85540 14764 85546 14776
rect 273346 14764 273352 14776
rect 273404 14764 273410 14816
rect 82722 14696 82728 14748
rect 82780 14736 82786 14748
rect 270681 14739 270739 14745
rect 270681 14736 270693 14739
rect 82780 14708 270693 14736
rect 82780 14696 82786 14708
rect 270681 14705 270693 14708
rect 270727 14705 270739 14739
rect 270681 14699 270739 14705
rect 78582 14628 78588 14680
rect 78640 14668 78646 14680
rect 269206 14668 269212 14680
rect 78640 14640 269212 14668
rect 78640 14628 78646 14640
rect 269206 14628 269212 14640
rect 269264 14628 269270 14680
rect 74442 14560 74448 14612
rect 74500 14600 74506 14612
rect 267826 14600 267832 14612
rect 74500 14572 267832 14600
rect 74500 14560 74506 14572
rect 267826 14560 267832 14572
rect 267884 14560 267890 14612
rect 71682 14492 71688 14544
rect 71740 14532 71746 14544
rect 265158 14532 265164 14544
rect 71740 14504 265164 14532
rect 71740 14492 71746 14504
rect 265158 14492 265164 14504
rect 265216 14492 265222 14544
rect 329926 14492 329932 14544
rect 329984 14532 329990 14544
rect 330110 14532 330116 14544
rect 329984 14504 330116 14532
rect 329984 14492 329990 14504
rect 330110 14492 330116 14504
rect 330168 14492 330174 14544
rect 23382 14424 23388 14476
rect 23440 14464 23446 14476
rect 241698 14464 241704 14476
rect 23440 14436 241704 14464
rect 23440 14424 23446 14436
rect 241698 14424 241704 14436
rect 241756 14424 241762 14476
rect 244182 14424 244188 14476
rect 244240 14464 244246 14476
rect 354766 14464 354772 14476
rect 244240 14436 354772 14464
rect 244240 14424 244246 14436
rect 354766 14424 354772 14436
rect 354824 14424 354830 14476
rect 160002 14356 160008 14408
rect 160060 14396 160066 14408
rect 311986 14396 311992 14408
rect 160060 14368 311992 14396
rect 160060 14356 160066 14368
rect 311986 14356 311992 14368
rect 312044 14356 312050 14408
rect 157242 14288 157248 14340
rect 157300 14328 157306 14340
rect 309410 14328 309416 14340
rect 157300 14300 309416 14328
rect 157300 14288 157306 14300
rect 309410 14288 309416 14300
rect 309468 14288 309474 14340
rect 165522 14220 165528 14272
rect 165580 14260 165586 14272
rect 313458 14260 313464 14272
rect 165580 14232 313464 14260
rect 165580 14220 165586 14232
rect 313458 14220 313464 14232
rect 313516 14220 313522 14272
rect 168282 14152 168288 14204
rect 168340 14192 168346 14204
rect 316126 14192 316132 14204
rect 168340 14164 316132 14192
rect 168340 14152 168346 14164
rect 316126 14152 316132 14164
rect 316184 14152 316190 14204
rect 117222 14084 117228 14136
rect 117280 14124 117286 14136
rect 246298 14124 246304 14136
rect 117280 14096 246304 14124
rect 117280 14084 117286 14096
rect 246298 14084 246304 14096
rect 246356 14084 246362 14136
rect 240042 14016 240048 14068
rect 240100 14056 240106 14068
rect 352006 14056 352012 14068
rect 240100 14028 352012 14056
rect 240100 14016 240106 14028
rect 352006 14016 352012 14028
rect 352064 14016 352070 14068
rect 202782 13744 202788 13796
rect 202840 13784 202846 13796
rect 334158 13784 334164 13796
rect 202840 13756 334164 13784
rect 202840 13744 202846 13756
rect 334158 13744 334164 13756
rect 334216 13744 334222 13796
rect 159910 13676 159916 13728
rect 159968 13716 159974 13728
rect 310698 13716 310704 13728
rect 159968 13688 310704 13716
rect 159968 13676 159974 13688
rect 310698 13676 310704 13688
rect 310756 13676 310762 13728
rect 155862 13608 155868 13660
rect 155920 13648 155926 13660
rect 309134 13648 309140 13660
rect 155920 13620 309140 13648
rect 155920 13608 155926 13620
rect 309134 13608 309140 13620
rect 309192 13608 309198 13660
rect 153102 13540 153108 13592
rect 153160 13580 153166 13592
rect 307846 13580 307852 13592
rect 153160 13552 307852 13580
rect 153160 13540 153166 13552
rect 307846 13540 307852 13552
rect 307904 13540 307910 13592
rect 148962 13472 148968 13524
rect 149020 13512 149026 13524
rect 305086 13512 305092 13524
rect 149020 13484 305092 13512
rect 149020 13472 149026 13484
rect 305086 13472 305092 13484
rect 305144 13472 305150 13524
rect 150342 13404 150348 13456
rect 150400 13444 150406 13456
rect 306466 13444 306472 13456
rect 150400 13416 306472 13444
rect 150400 13404 150406 13416
rect 306466 13404 306472 13416
rect 306524 13404 306530 13456
rect 151722 13336 151728 13388
rect 151780 13376 151786 13388
rect 307938 13376 307944 13388
rect 151780 13348 307944 13376
rect 151780 13336 151786 13348
rect 307938 13336 307944 13348
rect 307996 13336 308002 13388
rect 146202 13268 146208 13320
rect 146260 13308 146266 13320
rect 303614 13308 303620 13320
rect 146260 13280 303620 13308
rect 146260 13268 146266 13280
rect 303614 13268 303620 13280
rect 303672 13268 303678 13320
rect 144822 13200 144828 13252
rect 144880 13240 144886 13252
rect 303706 13240 303712 13252
rect 144880 13212 303712 13240
rect 144880 13200 144886 13212
rect 303706 13200 303712 13212
rect 303764 13200 303770 13252
rect 132402 13132 132408 13184
rect 132460 13172 132466 13184
rect 296898 13172 296904 13184
rect 132460 13144 296904 13172
rect 132460 13132 132466 13144
rect 296898 13132 296904 13144
rect 296956 13132 296962 13184
rect 19242 13064 19248 13116
rect 19300 13104 19306 13116
rect 238846 13104 238852 13116
rect 19300 13076 238852 13104
rect 19300 13064 19306 13076
rect 238846 13064 238852 13076
rect 238904 13064 238910 13116
rect 200022 12996 200028 13048
rect 200080 13036 200086 13048
rect 331398 13036 331404 13048
rect 200080 13008 331404 13036
rect 200080 12996 200086 13008
rect 331398 12996 331404 13008
rect 331456 12996 331462 13048
rect 206922 12928 206928 12980
rect 206980 12968 206986 12980
rect 335446 12968 335452 12980
rect 206980 12940 335452 12968
rect 206980 12928 206986 12940
rect 335446 12928 335452 12940
rect 335504 12928 335510 12980
rect 213822 12860 213828 12912
rect 213880 12900 213886 12912
rect 339678 12900 339684 12912
rect 213880 12872 339684 12900
rect 213880 12860 213886 12872
rect 339678 12860 339684 12872
rect 339736 12860 339742 12912
rect 211062 12792 211068 12844
rect 211120 12832 211126 12844
rect 336826 12832 336832 12844
rect 211120 12804 336832 12832
rect 211120 12792 211126 12804
rect 336826 12792 336832 12804
rect 336884 12792 336890 12844
rect 217962 12724 217968 12776
rect 218020 12764 218026 12776
rect 340966 12764 340972 12776
rect 218020 12736 340972 12764
rect 218020 12724 218026 12736
rect 340966 12724 340972 12736
rect 341024 12724 341030 12776
rect 220722 12656 220728 12708
rect 220780 12696 220786 12708
rect 342346 12696 342352 12708
rect 220780 12668 342352 12696
rect 220780 12656 220786 12668
rect 342346 12656 342352 12668
rect 342404 12656 342410 12708
rect 260929 12563 260987 12569
rect 260929 12529 260941 12563
rect 260975 12560 260987 12563
rect 261018 12560 261024 12572
rect 260975 12532 261024 12560
rect 260975 12529 260987 12532
rect 260929 12523 260987 12529
rect 261018 12520 261024 12532
rect 261076 12520 261082 12572
rect 232777 12495 232835 12501
rect 232777 12461 232789 12495
rect 232823 12492 232835 12495
rect 236178 12492 236184 12504
rect 232823 12464 236184 12492
rect 232823 12461 232835 12464
rect 232777 12455 232835 12461
rect 236178 12452 236184 12464
rect 236236 12452 236242 12504
rect 293954 12492 293960 12504
rect 293915 12464 293960 12492
rect 293954 12452 293960 12464
rect 294012 12452 294018 12504
rect 397638 12492 397644 12504
rect 397564 12464 397644 12492
rect 397564 12436 397592 12464
rect 397638 12452 397644 12464
rect 397696 12452 397702 12504
rect 184842 12384 184848 12436
rect 184900 12424 184906 12436
rect 323118 12424 323124 12436
rect 184900 12396 323124 12424
rect 184900 12384 184906 12396
rect 323118 12384 323124 12396
rect 323176 12384 323182 12436
rect 347866 12424 347872 12436
rect 347827 12396 347872 12424
rect 347866 12384 347872 12396
rect 347924 12384 347930 12436
rect 397546 12384 397552 12436
rect 397604 12384 397610 12436
rect 180702 12316 180708 12368
rect 180760 12356 180766 12368
rect 321738 12356 321744 12368
rect 180760 12328 321744 12356
rect 180760 12316 180766 12328
rect 321738 12316 321744 12328
rect 321796 12316 321802 12368
rect 427906 12316 427912 12368
rect 427964 12356 427970 12368
rect 428090 12356 428096 12368
rect 427964 12328 428096 12356
rect 427964 12316 427970 12328
rect 428090 12316 428096 12328
rect 428148 12316 428154 12368
rect 176562 12248 176568 12300
rect 176620 12288 176626 12300
rect 320266 12288 320272 12300
rect 176620 12260 320272 12288
rect 176620 12248 176626 12260
rect 320266 12248 320272 12260
rect 320324 12248 320330 12300
rect 416958 12288 416964 12300
rect 416919 12260 416964 12288
rect 416958 12248 416964 12260
rect 417016 12248 417022 12300
rect 173802 12180 173808 12232
rect 173860 12220 173866 12232
rect 317598 12220 317604 12232
rect 173860 12192 317604 12220
rect 173860 12180 173866 12192
rect 317598 12180 317604 12192
rect 317656 12180 317662 12232
rect 169662 12112 169668 12164
rect 169720 12152 169726 12164
rect 316034 12152 316040 12164
rect 169720 12124 316040 12152
rect 169720 12112 169726 12124
rect 316034 12112 316040 12124
rect 316092 12112 316098 12164
rect 166902 12044 166908 12096
rect 166960 12084 166966 12096
rect 314746 12084 314752 12096
rect 166960 12056 314752 12084
rect 166960 12044 166966 12056
rect 314746 12044 314752 12056
rect 314804 12044 314810 12096
rect 162762 11976 162768 12028
rect 162820 12016 162826 12028
rect 313366 12016 313372 12028
rect 162820 11988 313372 12016
rect 162820 11976 162826 11988
rect 313366 11976 313372 11988
rect 313424 11976 313430 12028
rect 142062 11908 142068 11960
rect 142120 11948 142126 11960
rect 302418 11948 302424 11960
rect 142120 11920 302424 11948
rect 142120 11908 142126 11920
rect 302418 11908 302424 11920
rect 302476 11908 302482 11960
rect 126882 11840 126888 11892
rect 126940 11880 126946 11892
rect 293957 11883 294015 11889
rect 293957 11880 293969 11883
rect 126940 11852 293969 11880
rect 126940 11840 126946 11852
rect 293957 11849 293969 11852
rect 294003 11849 294015 11883
rect 293957 11843 294015 11849
rect 128262 11772 128268 11824
rect 128320 11812 128326 11824
rect 295334 11812 295340 11824
rect 128320 11784 295340 11812
rect 128320 11772 128326 11784
rect 295334 11772 295340 11784
rect 295392 11772 295398 11824
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 232777 11747 232835 11753
rect 232777 11744 232789 11747
rect 13688 11716 232789 11744
rect 13688 11704 13694 11716
rect 232777 11713 232789 11716
rect 232823 11713 232835 11747
rect 260926 11744 260932 11756
rect 260887 11716 260932 11744
rect 232777 11707 232835 11713
rect 260926 11704 260932 11716
rect 260984 11704 260990 11756
rect 187602 11636 187608 11688
rect 187660 11676 187666 11688
rect 325786 11676 325792 11688
rect 187660 11648 325792 11676
rect 187660 11636 187666 11648
rect 325786 11636 325792 11648
rect 325844 11636 325850 11688
rect 191742 11568 191748 11620
rect 191800 11608 191806 11620
rect 327258 11608 327264 11620
rect 191800 11580 327264 11608
rect 191800 11568 191806 11580
rect 327258 11568 327264 11580
rect 327316 11568 327322 11620
rect 194502 11500 194508 11552
rect 194560 11540 194566 11552
rect 328638 11540 328644 11552
rect 194560 11512 328644 11540
rect 194560 11500 194566 11512
rect 328638 11500 328644 11512
rect 328696 11500 328702 11552
rect 198642 11432 198648 11484
rect 198700 11472 198706 11484
rect 331214 11472 331220 11484
rect 198700 11444 331220 11472
rect 198700 11432 198706 11444
rect 331214 11432 331220 11444
rect 331272 11432 331278 11484
rect 201494 11364 201500 11416
rect 201552 11404 201558 11416
rect 332778 11404 332784 11416
rect 201552 11376 332784 11404
rect 201552 11364 201558 11376
rect 332778 11364 332784 11376
rect 332836 11364 332842 11416
rect 205542 11296 205548 11348
rect 205600 11336 205606 11348
rect 334434 11336 334440 11348
rect 205600 11308 334440 11336
rect 205600 11296 205606 11308
rect 334434 11296 334440 11308
rect 334492 11296 334498 11348
rect 143442 10956 143448 11008
rect 143500 10996 143506 11008
rect 302326 10996 302332 11008
rect 143500 10968 302332 10996
rect 143500 10956 143506 10968
rect 302326 10956 302332 10968
rect 302384 10956 302390 11008
rect 140682 10888 140688 10940
rect 140740 10928 140746 10940
rect 301038 10928 301044 10940
rect 140740 10900 301044 10928
rect 140740 10888 140746 10900
rect 301038 10888 301044 10900
rect 301096 10888 301102 10940
rect 124122 10820 124128 10872
rect 124180 10860 124186 10872
rect 292574 10860 292580 10872
rect 124180 10832 292580 10860
rect 124180 10820 124186 10832
rect 292574 10820 292580 10832
rect 292632 10820 292638 10872
rect 119982 10752 119988 10804
rect 120040 10792 120046 10804
rect 291194 10792 291200 10804
rect 120040 10764 291200 10792
rect 120040 10752 120046 10764
rect 291194 10752 291200 10764
rect 291252 10752 291258 10804
rect 117130 10684 117136 10736
rect 117188 10724 117194 10736
rect 288342 10724 288348 10736
rect 117188 10696 288348 10724
rect 117188 10684 117194 10696
rect 288342 10684 288348 10696
rect 288400 10684 288406 10736
rect 113082 10616 113088 10668
rect 113140 10656 113146 10668
rect 287054 10656 287060 10668
rect 113140 10628 287060 10656
rect 113140 10616 113146 10628
rect 287054 10616 287060 10628
rect 287112 10616 287118 10668
rect 289814 10616 289820 10668
rect 289872 10656 289878 10668
rect 367186 10656 367192 10668
rect 289872 10628 367192 10656
rect 289872 10616 289878 10628
rect 367186 10616 367192 10628
rect 367244 10616 367250 10668
rect 108758 10548 108764 10600
rect 108816 10588 108822 10600
rect 285674 10588 285680 10600
rect 108816 10560 285680 10588
rect 108816 10548 108822 10560
rect 285674 10548 285680 10560
rect 285732 10548 285738 10600
rect 289906 10548 289912 10600
rect 289964 10588 289970 10600
rect 367278 10588 367284 10600
rect 289964 10560 367284 10588
rect 289964 10548 289970 10560
rect 367278 10548 367284 10560
rect 367336 10548 367342 10600
rect 105170 10480 105176 10532
rect 105228 10520 105234 10532
rect 283190 10520 283196 10532
rect 105228 10492 283196 10520
rect 105228 10480 105234 10492
rect 283190 10480 283196 10492
rect 283248 10480 283254 10532
rect 287606 10480 287612 10532
rect 287664 10520 287670 10532
rect 365622 10520 365628 10532
rect 287664 10492 365628 10520
rect 287664 10480 287670 10492
rect 365622 10480 365628 10492
rect 365680 10480 365686 10532
rect 101582 10412 101588 10464
rect 101640 10452 101646 10464
rect 281534 10452 281540 10464
rect 101640 10424 281540 10452
rect 101640 10412 101646 10424
rect 281534 10412 281540 10424
rect 281592 10412 281598 10464
rect 299658 10412 299664 10464
rect 299716 10452 299722 10464
rect 379606 10452 379612 10464
rect 299716 10424 379612 10452
rect 299716 10412 299722 10424
rect 379606 10412 379612 10424
rect 379664 10412 379670 10464
rect 99190 10344 99196 10396
rect 99248 10384 99254 10396
rect 280154 10384 280160 10396
rect 99248 10356 280160 10384
rect 99248 10344 99254 10356
rect 280154 10344 280160 10356
rect 280212 10344 280218 10396
rect 300946 10344 300952 10396
rect 301004 10384 301010 10396
rect 383746 10384 383752 10396
rect 301004 10356 383752 10384
rect 301004 10344 301010 10356
rect 383746 10344 383752 10356
rect 383804 10344 383810 10396
rect 64782 10276 64788 10328
rect 64840 10316 64846 10328
rect 262306 10316 262312 10328
rect 64840 10288 262312 10316
rect 64840 10276 64846 10288
rect 262306 10276 262312 10288
rect 262364 10276 262370 10328
rect 292942 10276 292948 10328
rect 293000 10316 293006 10328
rect 378318 10316 378324 10328
rect 293000 10288 378324 10316
rect 293000 10276 293006 10288
rect 378318 10276 378324 10288
rect 378376 10276 378382 10328
rect 147582 10208 147588 10260
rect 147640 10248 147646 10260
rect 304994 10248 305000 10260
rect 147640 10220 305000 10248
rect 147640 10208 147646 10220
rect 304994 10208 305000 10220
rect 305052 10208 305058 10260
rect 151630 10140 151636 10192
rect 151688 10180 151694 10192
rect 306374 10180 306380 10192
rect 151688 10152 306380 10180
rect 151688 10140 151694 10152
rect 306374 10140 306380 10152
rect 306432 10140 306438 10192
rect 154482 10072 154488 10124
rect 154540 10112 154546 10124
rect 307846 10112 307852 10124
rect 154540 10084 307852 10112
rect 154540 10072 154546 10084
rect 307846 10072 307852 10084
rect 307904 10072 307910 10124
rect 158622 10004 158628 10056
rect 158680 10044 158686 10056
rect 310514 10044 310520 10056
rect 158680 10016 310520 10044
rect 158680 10004 158686 10016
rect 310514 10004 310520 10016
rect 310572 10004 310578 10056
rect 161382 9936 161388 9988
rect 161440 9976 161446 9988
rect 311894 9976 311900 9988
rect 161440 9948 311900 9976
rect 161440 9936 161446 9948
rect 311894 9936 311900 9948
rect 311952 9936 311958 9988
rect 246758 9868 246764 9920
rect 246816 9908 246822 9920
rect 356238 9908 356244 9920
rect 246816 9880 356244 9908
rect 246816 9868 246822 9880
rect 356238 9868 356244 9880
rect 356296 9868 356302 9920
rect 250346 9800 250352 9852
rect 250404 9840 250410 9852
rect 357618 9840 357624 9852
rect 250404 9812 357624 9840
rect 250404 9800 250410 9812
rect 357618 9800 357624 9812
rect 357676 9800 357682 9852
rect 253842 9732 253848 9784
rect 253900 9772 253906 9784
rect 360286 9772 360292 9784
rect 253900 9744 360292 9772
rect 253900 9732 253906 9744
rect 360286 9732 360292 9744
rect 360344 9732 360350 9784
rect 244274 9664 244280 9716
rect 244332 9704 244338 9716
rect 244550 9704 244556 9716
rect 244332 9676 244556 9704
rect 244332 9664 244338 9676
rect 244550 9664 244556 9676
rect 244608 9664 244614 9716
rect 249978 9664 249984 9716
rect 250036 9704 250042 9716
rect 250070 9704 250076 9716
rect 250036 9676 250076 9704
rect 250036 9664 250042 9676
rect 250070 9664 250076 9676
rect 250128 9664 250134 9716
rect 257430 9664 257436 9716
rect 257488 9704 257494 9716
rect 361758 9704 361764 9716
rect 257488 9676 361764 9704
rect 257488 9664 257494 9676
rect 361758 9664 361764 9676
rect 361816 9664 361822 9716
rect 386506 9664 386512 9716
rect 386564 9704 386570 9716
rect 386782 9704 386788 9716
rect 386564 9676 386788 9704
rect 386564 9664 386570 9676
rect 386782 9664 386788 9676
rect 386840 9664 386846 9716
rect 387886 9664 387892 9716
rect 387944 9704 387950 9716
rect 388070 9704 388076 9716
rect 387944 9676 388076 9704
rect 387944 9664 387950 9676
rect 388070 9664 388076 9676
rect 388128 9664 388134 9716
rect 422294 9664 422300 9716
rect 422352 9704 422358 9716
rect 422478 9704 422484 9716
rect 422352 9676 422484 9704
rect 422352 9664 422358 9676
rect 422478 9664 422484 9676
rect 422536 9664 422542 9716
rect 203886 9596 203892 9648
rect 203944 9636 203950 9648
rect 333974 9636 333980 9648
rect 203944 9608 333980 9636
rect 203944 9596 203950 9608
rect 333974 9596 333980 9608
rect 334032 9596 334038 9648
rect 346486 9636 346492 9648
rect 346447 9608 346492 9636
rect 346486 9596 346492 9608
rect 346544 9596 346550 9648
rect 393038 9636 393044 9648
rect 392999 9608 393044 9636
rect 393038 9596 393044 9608
rect 393096 9596 393102 9648
rect 200390 9528 200396 9580
rect 200448 9568 200454 9580
rect 332594 9568 332600 9580
rect 200448 9540 332600 9568
rect 200448 9528 200454 9540
rect 332594 9528 332600 9540
rect 332652 9528 332658 9580
rect 196802 9460 196808 9512
rect 196860 9500 196866 9512
rect 330018 9500 330024 9512
rect 196860 9472 330024 9500
rect 196860 9460 196866 9472
rect 330018 9460 330024 9472
rect 330076 9460 330082 9512
rect 193214 9392 193220 9444
rect 193272 9432 193278 9444
rect 328730 9432 328736 9444
rect 193272 9404 328736 9432
rect 193272 9392 193278 9404
rect 328730 9392 328736 9404
rect 328788 9392 328794 9444
rect 189626 9324 189632 9376
rect 189684 9364 189690 9376
rect 327074 9364 327080 9376
rect 189684 9336 327080 9364
rect 189684 9324 189690 9336
rect 327074 9324 327080 9336
rect 327132 9324 327138 9376
rect 186038 9256 186044 9308
rect 186096 9296 186102 9308
rect 324406 9296 324412 9308
rect 186096 9268 324412 9296
rect 186096 9256 186102 9268
rect 324406 9256 324412 9268
rect 324464 9256 324470 9308
rect 361666 9296 361672 9308
rect 325344 9268 361672 9296
rect 182542 9188 182548 9240
rect 182600 9228 182606 9240
rect 323210 9228 323216 9240
rect 182600 9200 323216 9228
rect 182600 9188 182606 9200
rect 323210 9188 323216 9200
rect 323268 9188 323274 9240
rect 178954 9120 178960 9172
rect 179012 9160 179018 9172
rect 321554 9160 321560 9172
rect 179012 9132 321560 9160
rect 179012 9120 179018 9132
rect 321554 9120 321560 9132
rect 321612 9120 321618 9172
rect 322566 9120 322572 9172
rect 322624 9160 322630 9172
rect 325344 9160 325372 9268
rect 361666 9256 361672 9268
rect 361724 9256 361730 9308
rect 327074 9188 327080 9240
rect 327132 9228 327138 9240
rect 392026 9228 392032 9240
rect 327132 9200 392032 9228
rect 327132 9188 327138 9200
rect 392026 9188 392032 9200
rect 392084 9188 392090 9240
rect 322624 9132 325372 9160
rect 322624 9120 322630 9132
rect 325510 9120 325516 9172
rect 325568 9160 325574 9172
rect 390646 9160 390652 9172
rect 325568 9132 390652 9160
rect 325568 9120 325574 9132
rect 390646 9120 390652 9132
rect 390704 9120 390710 9172
rect 175366 9052 175372 9104
rect 175424 9092 175430 9104
rect 318886 9092 318892 9104
rect 175424 9064 318892 9092
rect 175424 9052 175430 9064
rect 318886 9052 318892 9064
rect 318944 9052 318950 9104
rect 328546 9052 328552 9104
rect 328604 9092 328610 9104
rect 394786 9092 394792 9104
rect 328604 9064 394792 9092
rect 328604 9052 328610 9064
rect 394786 9052 394792 9064
rect 394844 9052 394850 9104
rect 171778 8984 171784 9036
rect 171836 9024 171842 9036
rect 317690 9024 317696 9036
rect 171836 8996 317696 9024
rect 171836 8984 171842 8996
rect 317690 8984 317696 8996
rect 317748 8984 317754 9036
rect 323578 8984 323584 9036
rect 323636 9024 323642 9036
rect 389266 9024 389272 9036
rect 323636 8996 389272 9024
rect 323636 8984 323642 8996
rect 389266 8984 389272 8996
rect 389324 8984 389330 9036
rect 132586 8916 132592 8968
rect 132644 8956 132650 8968
rect 296806 8956 296812 8968
rect 132644 8928 296812 8956
rect 132644 8916 132650 8928
rect 296806 8916 296812 8928
rect 296864 8916 296870 8968
rect 334710 8916 334716 8968
rect 334768 8956 334774 8968
rect 401686 8956 401692 8968
rect 334768 8928 401692 8956
rect 334768 8916 334774 8928
rect 401686 8916 401692 8928
rect 401744 8916 401750 8968
rect 210970 8848 210976 8900
rect 211028 8888 211034 8900
rect 338206 8888 338212 8900
rect 211028 8860 338212 8888
rect 211028 8848 211034 8860
rect 338206 8848 338212 8860
rect 338264 8848 338270 8900
rect 207474 8780 207480 8832
rect 207532 8820 207538 8832
rect 335354 8820 335360 8832
rect 207532 8792 335360 8820
rect 207532 8780 207538 8792
rect 335354 8780 335360 8792
rect 335412 8780 335418 8832
rect 214650 8712 214656 8764
rect 214708 8752 214714 8764
rect 339770 8752 339776 8764
rect 214708 8724 339776 8752
rect 214708 8712 214714 8724
rect 339770 8712 339776 8724
rect 339828 8712 339834 8764
rect 221734 8644 221740 8696
rect 221792 8684 221798 8696
rect 343726 8684 343732 8696
rect 221792 8656 343732 8684
rect 221792 8644 221798 8656
rect 343726 8644 343732 8656
rect 343784 8644 343790 8696
rect 218146 8576 218152 8628
rect 218204 8616 218210 8628
rect 340874 8616 340880 8628
rect 218204 8588 340880 8616
rect 218204 8576 218210 8588
rect 340874 8576 340880 8588
rect 340932 8576 340938 8628
rect 225322 8508 225328 8560
rect 225380 8548 225386 8560
rect 345198 8548 345204 8560
rect 225380 8520 345204 8548
rect 225380 8508 225386 8520
rect 345198 8508 345204 8520
rect 345256 8508 345262 8560
rect 228910 8440 228916 8492
rect 228968 8480 228974 8492
rect 346489 8483 346547 8489
rect 346489 8480 346501 8483
rect 228968 8452 346501 8480
rect 228968 8440 228974 8452
rect 346489 8449 346501 8452
rect 346535 8449 346547 8483
rect 346489 8443 346547 8449
rect 232498 8372 232504 8424
rect 232556 8412 232562 8424
rect 349246 8412 349252 8424
rect 232556 8384 349252 8412
rect 232556 8372 232562 8384
rect 349246 8372 349252 8384
rect 349304 8372 349310 8424
rect 230658 8344 230664 8356
rect 230619 8316 230664 8344
rect 230658 8304 230664 8316
rect 230716 8304 230722 8356
rect 235994 8304 236000 8356
rect 236052 8344 236058 8356
rect 350718 8344 350724 8356
rect 236052 8316 350724 8344
rect 236052 8304 236058 8316
rect 350718 8304 350724 8316
rect 350776 8304 350782 8356
rect 380986 8344 380992 8356
rect 380947 8316 380992 8344
rect 380986 8304 380992 8316
rect 381044 8304 381050 8356
rect 382366 8344 382372 8356
rect 382327 8316 382372 8344
rect 382366 8304 382372 8316
rect 382424 8304 382430 8356
rect 400398 8344 400404 8356
rect 400359 8316 400404 8344
rect 400398 8304 400404 8316
rect 400456 8304 400462 8356
rect 56410 8236 56416 8288
rect 56468 8276 56474 8288
rect 258350 8276 258356 8288
rect 56468 8248 258356 8276
rect 56468 8236 56474 8248
rect 258350 8236 258356 8248
rect 258408 8236 258414 8288
rect 274082 8236 274088 8288
rect 274140 8276 274146 8288
rect 370130 8276 370136 8288
rect 274140 8248 370136 8276
rect 274140 8236 274146 8248
rect 370130 8236 370136 8248
rect 370188 8236 370194 8288
rect 52822 8168 52828 8220
rect 52880 8208 52886 8220
rect 256786 8208 256792 8220
rect 52880 8180 256792 8208
rect 52880 8168 52886 8180
rect 256786 8168 256792 8180
rect 256844 8168 256850 8220
rect 270494 8168 270500 8220
rect 270552 8208 270558 8220
rect 368566 8208 368572 8220
rect 270552 8180 368572 8208
rect 270552 8168 270558 8180
rect 368566 8168 368572 8180
rect 368624 8168 368630 8220
rect 49326 8100 49332 8152
rect 49384 8140 49390 8152
rect 254026 8140 254032 8152
rect 49384 8112 254032 8140
rect 49384 8100 49390 8112
rect 254026 8100 254032 8112
rect 254084 8100 254090 8152
rect 266998 8100 267004 8152
rect 267056 8140 267062 8152
rect 367094 8140 367100 8152
rect 267056 8112 367100 8140
rect 267056 8100 267062 8112
rect 367094 8100 367100 8112
rect 367152 8100 367158 8152
rect 44542 8032 44548 8084
rect 44600 8072 44606 8084
rect 252646 8072 252652 8084
rect 44600 8044 252652 8072
rect 44600 8032 44606 8044
rect 252646 8032 252652 8044
rect 252704 8032 252710 8084
rect 263410 8032 263416 8084
rect 263468 8072 263474 8084
rect 364518 8072 364524 8084
rect 263468 8044 364524 8072
rect 263468 8032 263474 8044
rect 364518 8032 364524 8044
rect 364576 8032 364582 8084
rect 40954 7964 40960 8016
rect 41012 8004 41018 8016
rect 249978 8004 249984 8016
rect 41012 7976 249984 8004
rect 41012 7964 41018 7976
rect 249978 7964 249984 7976
rect 250036 7964 250042 8016
rect 259822 7964 259828 8016
rect 259880 8004 259886 8016
rect 363046 8004 363052 8016
rect 259880 7976 363052 8004
rect 259880 7964 259886 7976
rect 363046 7964 363052 7976
rect 363104 7964 363110 8016
rect 37366 7896 37372 7948
rect 37424 7936 37430 7948
rect 248506 7936 248512 7948
rect 37424 7908 248512 7936
rect 37424 7896 37430 7908
rect 248506 7896 248512 7908
rect 248564 7896 248570 7948
rect 256234 7896 256240 7948
rect 256292 7936 256298 7948
rect 361574 7936 361580 7948
rect 256292 7908 361580 7936
rect 256292 7896 256298 7908
rect 361574 7896 361580 7908
rect 361632 7896 361638 7948
rect 33870 7828 33876 7880
rect 33928 7868 33934 7880
rect 247218 7868 247224 7880
rect 33928 7840 247224 7868
rect 33928 7828 33934 7840
rect 247218 7828 247224 7840
rect 247276 7828 247282 7880
rect 252646 7828 252652 7880
rect 252704 7868 252710 7880
rect 358998 7868 359004 7880
rect 252704 7840 359004 7868
rect 252704 7828 252710 7840
rect 358998 7828 359004 7840
rect 359056 7828 359062 7880
rect 30282 7760 30288 7812
rect 30340 7800 30346 7812
rect 244274 7800 244280 7812
rect 30340 7772 244280 7800
rect 30340 7760 30346 7772
rect 244274 7760 244280 7772
rect 244332 7760 244338 7812
rect 249150 7760 249156 7812
rect 249208 7800 249214 7812
rect 357434 7800 357440 7812
rect 249208 7772 357440 7800
rect 249208 7760 249214 7772
rect 357434 7760 357440 7772
rect 357492 7760 357498 7812
rect 26694 7692 26700 7744
rect 26752 7732 26758 7744
rect 242894 7732 242900 7744
rect 26752 7704 242900 7732
rect 26752 7692 26758 7704
rect 242894 7692 242900 7704
rect 242952 7692 242958 7744
rect 245562 7692 245568 7744
rect 245620 7732 245626 7744
rect 356146 7732 356152 7744
rect 245620 7704 356152 7732
rect 245620 7692 245626 7704
rect 356146 7692 356152 7704
rect 356204 7692 356210 7744
rect 8846 7624 8852 7676
rect 8904 7664 8910 7676
rect 233326 7664 233332 7676
rect 8904 7636 233332 7664
rect 8904 7624 8910 7636
rect 233326 7624 233332 7636
rect 233384 7624 233390 7676
rect 234798 7624 234804 7676
rect 234856 7664 234862 7676
rect 350626 7664 350632 7676
rect 234856 7636 350632 7664
rect 234856 7624 234862 7636
rect 350626 7624 350632 7636
rect 350684 7624 350690 7676
rect 3970 7556 3976 7608
rect 4028 7596 4034 7608
rect 230658 7596 230664 7608
rect 4028 7568 230664 7596
rect 4028 7556 4034 7568
rect 230658 7556 230664 7568
rect 230716 7556 230722 7608
rect 231302 7556 231308 7608
rect 231360 7596 231366 7608
rect 347866 7596 347872 7608
rect 231360 7568 347872 7596
rect 231360 7556 231366 7568
rect 347866 7556 347872 7568
rect 347924 7556 347930 7608
rect 351822 7556 351828 7608
rect 351880 7596 351886 7608
rect 405826 7596 405832 7608
rect 351880 7568 405832 7596
rect 351880 7556 351886 7568
rect 405826 7556 405832 7568
rect 405884 7556 405890 7608
rect 87322 7488 87328 7540
rect 87380 7528 87386 7540
rect 274634 7528 274640 7540
rect 87380 7500 274640 7528
rect 87380 7488 87386 7500
rect 274634 7488 274640 7500
rect 274692 7488 274698 7540
rect 277670 7488 277676 7540
rect 277728 7528 277734 7540
rect 372706 7528 372712 7540
rect 277728 7500 372712 7528
rect 277728 7488 277734 7500
rect 372706 7488 372712 7500
rect 372764 7488 372770 7540
rect 90910 7420 90916 7472
rect 90968 7460 90974 7472
rect 276014 7460 276020 7472
rect 90968 7432 276020 7460
rect 90968 7420 90974 7432
rect 276014 7420 276020 7432
rect 276072 7420 276078 7472
rect 281258 7420 281264 7472
rect 281316 7460 281322 7472
rect 374086 7460 374092 7472
rect 281316 7432 374092 7460
rect 281316 7420 281322 7432
rect 374086 7420 374092 7432
rect 374144 7420 374150 7472
rect 94498 7352 94504 7404
rect 94556 7392 94562 7404
rect 277578 7392 277584 7404
rect 94556 7364 277584 7392
rect 94556 7352 94562 7364
rect 277578 7352 277584 7364
rect 277636 7352 277642 7404
rect 284754 7352 284760 7404
rect 284812 7392 284818 7404
rect 375558 7392 375564 7404
rect 284812 7364 375564 7392
rect 284812 7352 284818 7364
rect 375558 7352 375564 7364
rect 375616 7352 375622 7404
rect 138474 7284 138480 7336
rect 138532 7324 138538 7336
rect 300854 7324 300860 7336
rect 138532 7296 300860 7324
rect 138532 7284 138538 7296
rect 300854 7284 300860 7296
rect 300912 7284 300918 7336
rect 347958 7284 347964 7336
rect 348016 7324 348022 7336
rect 397546 7324 397552 7336
rect 348016 7296 397552 7324
rect 348016 7284 348022 7296
rect 397546 7284 397552 7296
rect 397604 7284 397610 7336
rect 141970 7216 141976 7268
rect 142028 7256 142034 7268
rect 302510 7256 302516 7268
rect 142028 7228 302516 7256
rect 142028 7216 142034 7228
rect 302510 7216 302516 7228
rect 302568 7216 302574 7268
rect 346486 7216 346492 7268
rect 346544 7256 346550 7268
rect 396166 7256 396172 7268
rect 346544 7228 396172 7256
rect 346544 7216 346550 7228
rect 396166 7216 396172 7228
rect 396224 7216 396230 7268
rect 224126 7148 224132 7200
rect 224184 7188 224190 7200
rect 345106 7188 345112 7200
rect 224184 7160 345112 7188
rect 224184 7148 224190 7160
rect 345106 7148 345112 7160
rect 345164 7148 345170 7200
rect 227714 7080 227720 7132
rect 227772 7120 227778 7132
rect 346394 7120 346400 7132
rect 227772 7092 346400 7120
rect 227772 7080 227778 7092
rect 346394 7080 346400 7092
rect 346452 7080 346458 7132
rect 238386 7012 238392 7064
rect 238444 7052 238450 7064
rect 351914 7052 351920 7064
rect 238444 7024 351920 7052
rect 238444 7012 238450 7024
rect 351914 7012 351920 7024
rect 351972 7012 351978 7064
rect 241974 6944 241980 6996
rect 242032 6984 242038 6996
rect 353386 6984 353392 6996
rect 242032 6956 353392 6984
rect 242032 6944 242038 6956
rect 353386 6944 353392 6956
rect 353444 6944 353450 6996
rect 163498 6808 163504 6860
rect 163556 6848 163562 6860
rect 313550 6848 313556 6860
rect 163556 6820 313556 6848
rect 163556 6808 163562 6820
rect 313550 6808 313556 6820
rect 313608 6808 313614 6860
rect 349062 6808 349068 6860
rect 349120 6848 349126 6860
rect 408770 6848 408776 6860
rect 349120 6820 408776 6848
rect 349120 6808 349126 6820
rect 408770 6808 408776 6820
rect 408828 6808 408834 6860
rect 83826 6740 83832 6792
rect 83884 6780 83890 6792
rect 271874 6780 271880 6792
rect 83884 6752 271880 6780
rect 83884 6740 83890 6752
rect 271874 6740 271880 6752
rect 271932 6740 271938 6792
rect 315209 6783 315267 6789
rect 315209 6749 315221 6783
rect 315255 6780 315267 6783
rect 320174 6780 320180 6792
rect 315255 6752 320180 6780
rect 315255 6749 315267 6752
rect 315209 6743 315267 6749
rect 320174 6740 320180 6752
rect 320232 6740 320238 6792
rect 325602 6740 325608 6792
rect 325660 6780 325666 6792
rect 386506 6780 386512 6792
rect 325660 6752 386512 6780
rect 325660 6740 325666 6752
rect 386506 6740 386512 6752
rect 386564 6740 386570 6792
rect 80238 6672 80244 6724
rect 80296 6712 80302 6724
rect 270586 6712 270592 6724
rect 80296 6684 270592 6712
rect 80296 6672 80302 6684
rect 270586 6672 270592 6684
rect 270644 6672 270650 6724
rect 318794 6672 318800 6724
rect 318852 6712 318858 6724
rect 380986 6712 380992 6724
rect 318852 6684 380992 6712
rect 318852 6672 318858 6684
rect 380986 6672 380992 6684
rect 381044 6672 381050 6724
rect 76650 6604 76656 6656
rect 76708 6644 76714 6656
rect 269114 6644 269120 6656
rect 76708 6616 269120 6644
rect 76708 6604 76714 6616
rect 269114 6604 269120 6616
rect 269172 6604 269178 6656
rect 320174 6604 320180 6656
rect 320232 6644 320238 6656
rect 385126 6644 385132 6656
rect 320232 6616 385132 6644
rect 320232 6604 320238 6616
rect 385126 6604 385132 6616
rect 385184 6604 385190 6656
rect 73062 6536 73068 6588
rect 73120 6576 73126 6588
rect 266354 6576 266360 6588
rect 73120 6548 266360 6576
rect 73120 6536 73126 6548
rect 266354 6536 266360 6548
rect 266412 6536 266418 6588
rect 312170 6536 312176 6588
rect 312228 6576 312234 6588
rect 389358 6576 389364 6588
rect 312228 6548 389364 6576
rect 312228 6536 312234 6548
rect 389358 6536 389364 6548
rect 389416 6536 389422 6588
rect 69474 6468 69480 6520
rect 69532 6508 69538 6520
rect 264974 6508 264980 6520
rect 69532 6480 264980 6508
rect 69532 6468 69538 6480
rect 264974 6468 264980 6480
rect 265032 6468 265038 6520
rect 308582 6468 308588 6520
rect 308640 6508 308646 6520
rect 387886 6508 387892 6520
rect 308640 6480 387892 6508
rect 308640 6468 308646 6480
rect 387886 6468 387892 6480
rect 387944 6468 387950 6520
rect 62390 6400 62396 6452
rect 62448 6440 62454 6452
rect 260926 6440 260932 6452
rect 62448 6412 260932 6440
rect 62448 6400 62454 6412
rect 260926 6400 260932 6412
rect 260984 6400 260990 6452
rect 304994 6400 305000 6452
rect 305052 6440 305058 6452
rect 386414 6440 386420 6452
rect 305052 6412 386420 6440
rect 305052 6400 305058 6412
rect 386414 6400 386420 6412
rect 386472 6400 386478 6452
rect 65978 6332 65984 6384
rect 66036 6372 66042 6384
rect 263686 6372 263692 6384
rect 66036 6344 263692 6372
rect 66036 6332 66042 6344
rect 263686 6332 263692 6344
rect 263744 6332 263750 6384
rect 290734 6332 290740 6384
rect 290792 6372 290798 6384
rect 378226 6372 378232 6384
rect 290792 6344 378232 6372
rect 290792 6332 290798 6344
rect 378226 6332 378232 6344
rect 378284 6332 378290 6384
rect 58802 6264 58808 6316
rect 58860 6304 58866 6316
rect 259454 6304 259460 6316
rect 58860 6276 259460 6304
rect 58860 6264 58866 6276
rect 259454 6264 259460 6276
rect 259512 6264 259518 6316
rect 287146 6264 287152 6316
rect 287204 6304 287210 6316
rect 376938 6304 376944 6316
rect 287204 6276 376944 6304
rect 287204 6264 287210 6276
rect 376938 6264 376944 6276
rect 376996 6264 377002 6316
rect 55214 6196 55220 6248
rect 55272 6236 55278 6248
rect 258258 6236 258264 6248
rect 55272 6208 258264 6236
rect 55272 6196 55278 6208
rect 258258 6196 258264 6208
rect 258316 6196 258322 6248
rect 283650 6196 283656 6248
rect 283708 6236 283714 6248
rect 375374 6236 375380 6248
rect 283708 6208 375380 6236
rect 283708 6196 283714 6208
rect 375374 6196 375380 6208
rect 375432 6196 375438 6248
rect 379974 6196 379980 6248
rect 380032 6236 380038 6248
rect 425146 6236 425152 6248
rect 380032 6208 425152 6236
rect 380032 6196 380038 6208
rect 425146 6196 425152 6208
rect 425204 6196 425210 6248
rect 51626 6128 51632 6180
rect 51684 6168 51690 6180
rect 255314 6168 255320 6180
rect 51684 6140 255320 6168
rect 51684 6128 51690 6140
rect 255314 6128 255320 6140
rect 255372 6128 255378 6180
rect 279970 6128 279976 6180
rect 280028 6168 280034 6180
rect 372798 6168 372804 6180
rect 280028 6140 372804 6168
rect 280028 6128 280034 6140
rect 372798 6128 372804 6140
rect 372856 6128 372862 6180
rect 372890 6128 372896 6180
rect 372948 6168 372954 6180
rect 421098 6168 421104 6180
rect 372948 6140 421104 6168
rect 372948 6128 372954 6140
rect 421098 6128 421104 6140
rect 421156 6128 421162 6180
rect 167086 6060 167092 6112
rect 167144 6100 167150 6112
rect 314562 6100 314568 6112
rect 167144 6072 314568 6100
rect 167144 6060 167150 6072
rect 314562 6060 314568 6072
rect 314620 6060 314626 6112
rect 314654 6060 314660 6112
rect 314712 6100 314718 6112
rect 371326 6100 371332 6112
rect 314712 6072 371332 6100
rect 314712 6060 314718 6072
rect 371326 6060 371332 6072
rect 371384 6060 371390 6112
rect 170582 5992 170588 6044
rect 170640 6032 170646 6044
rect 317414 6032 317420 6044
rect 170640 6004 317420 6032
rect 170640 5992 170646 6004
rect 317414 5992 317420 6004
rect 317472 5992 317478 6044
rect 322201 6035 322259 6041
rect 322201 6001 322213 6035
rect 322247 6032 322259 6035
rect 322934 6032 322940 6044
rect 322247 6004 322940 6032
rect 322247 6001 322259 6004
rect 322201 5995 322259 6001
rect 322934 5992 322940 6004
rect 322992 5992 322998 6044
rect 354950 5992 354956 6044
rect 355008 6032 355014 6044
rect 411346 6032 411352 6044
rect 355008 6004 411352 6032
rect 355008 5992 355014 6004
rect 411346 5992 411352 6004
rect 411404 5992 411410 6044
rect 174170 5924 174176 5976
rect 174228 5964 174234 5976
rect 174228 5936 315344 5964
rect 174228 5924 174234 5936
rect 177758 5856 177764 5908
rect 177816 5896 177822 5908
rect 315209 5899 315267 5905
rect 315209 5896 315221 5899
rect 177816 5868 315221 5896
rect 177816 5856 177822 5868
rect 315209 5865 315221 5868
rect 315255 5865 315267 5899
rect 315316 5896 315344 5936
rect 316586 5924 316592 5976
rect 316644 5964 316650 5976
rect 369854 5964 369860 5976
rect 316644 5936 369860 5964
rect 316644 5924 316650 5936
rect 369854 5924 369860 5936
rect 369912 5924 369918 5976
rect 318886 5896 318892 5908
rect 315316 5868 318892 5896
rect 315209 5859 315267 5865
rect 318886 5856 318892 5868
rect 318944 5856 318950 5908
rect 325326 5856 325332 5908
rect 325384 5896 325390 5908
rect 360194 5896 360200 5908
rect 325384 5868 360200 5896
rect 325384 5856 325390 5868
rect 360194 5856 360200 5868
rect 360252 5856 360258 5908
rect 362126 5856 362132 5908
rect 362184 5896 362190 5908
rect 415578 5896 415584 5908
rect 362184 5868 415584 5896
rect 362184 5856 362190 5868
rect 415578 5856 415584 5868
rect 415636 5856 415642 5908
rect 181346 5788 181352 5840
rect 181404 5828 181410 5840
rect 322201 5831 322259 5837
rect 322201 5828 322213 5831
rect 181404 5800 322213 5828
rect 181404 5788 181410 5800
rect 322201 5797 322213 5800
rect 322247 5797 322259 5831
rect 322201 5791 322259 5797
rect 322658 5788 322664 5840
rect 322716 5828 322722 5840
rect 364334 5828 364340 5840
rect 322716 5800 364340 5828
rect 322716 5788 322722 5800
rect 364334 5788 364340 5800
rect 364392 5788 364398 5840
rect 369210 5788 369216 5840
rect 369268 5828 369274 5840
rect 419626 5828 419632 5840
rect 369268 5800 419632 5828
rect 369268 5788 369274 5800
rect 419626 5788 419632 5800
rect 419684 5788 419690 5840
rect 184842 5720 184848 5772
rect 184900 5760 184906 5772
rect 324314 5760 324320 5772
rect 184900 5732 324320 5760
rect 184900 5720 184906 5732
rect 324314 5720 324320 5732
rect 324372 5720 324378 5772
rect 188430 5652 188436 5704
rect 188488 5692 188494 5704
rect 325694 5692 325700 5704
rect 188488 5664 325700 5692
rect 188488 5652 188494 5664
rect 325694 5652 325700 5664
rect 325752 5652 325758 5704
rect 192018 5584 192024 5636
rect 192076 5624 192082 5636
rect 328454 5624 328460 5636
rect 192076 5596 328460 5624
rect 192076 5584 192082 5596
rect 328454 5584 328460 5596
rect 328512 5584 328518 5636
rect 195606 5516 195612 5568
rect 195664 5556 195670 5568
rect 329834 5556 329840 5568
rect 195664 5528 329840 5556
rect 195664 5516 195670 5528
rect 329834 5516 329840 5528
rect 329892 5516 329898 5568
rect 137278 5448 137284 5500
rect 137336 5488 137342 5500
rect 299474 5488 299480 5500
rect 137336 5460 299480 5488
rect 137336 5448 137342 5460
rect 299474 5448 299480 5460
rect 299532 5448 299538 5500
rect 315758 5448 315764 5500
rect 315816 5488 315822 5500
rect 391934 5488 391940 5500
rect 315816 5460 391940 5488
rect 315816 5448 315822 5460
rect 391934 5448 391940 5460
rect 391992 5448 391998 5500
rect 401318 5448 401324 5500
rect 401376 5488 401382 5500
rect 436186 5488 436192 5500
rect 401376 5460 436192 5488
rect 401376 5448 401382 5460
rect 436186 5448 436192 5460
rect 436244 5448 436250 5500
rect 133782 5380 133788 5432
rect 133840 5420 133846 5432
rect 298094 5420 298100 5432
rect 133840 5392 298100 5420
rect 133840 5380 133846 5392
rect 298094 5380 298100 5392
rect 298152 5380 298158 5432
rect 301406 5380 301412 5432
rect 301464 5420 301470 5432
rect 383838 5420 383844 5432
rect 301464 5392 383844 5420
rect 301464 5380 301470 5392
rect 383838 5380 383844 5392
rect 383896 5380 383902 5432
rect 397822 5380 397828 5432
rect 397880 5420 397886 5432
rect 433610 5420 433616 5432
rect 397880 5392 433616 5420
rect 397880 5380 397886 5392
rect 433610 5380 433616 5392
rect 433668 5380 433674 5432
rect 130194 5312 130200 5364
rect 130252 5352 130258 5364
rect 296714 5352 296720 5364
rect 130252 5324 296720 5352
rect 130252 5312 130258 5324
rect 296714 5312 296720 5324
rect 296772 5312 296778 5364
rect 297910 5312 297916 5364
rect 297968 5352 297974 5364
rect 382366 5352 382372 5364
rect 297968 5324 382372 5352
rect 297968 5312 297974 5324
rect 382366 5312 382372 5324
rect 382424 5312 382430 5364
rect 394234 5312 394240 5364
rect 394292 5352 394298 5364
rect 432138 5352 432144 5364
rect 394292 5324 432144 5352
rect 394292 5312 394298 5324
rect 432138 5312 432144 5324
rect 432196 5312 432202 5364
rect 67174 5244 67180 5296
rect 67232 5284 67238 5296
rect 263778 5284 263784 5296
rect 67232 5256 263784 5284
rect 67232 5244 67238 5256
rect 263778 5244 263784 5256
rect 263836 5244 263842 5296
rect 294322 5244 294328 5296
rect 294380 5284 294386 5296
rect 380894 5284 380900 5296
rect 294380 5256 380900 5284
rect 294380 5244 294386 5256
rect 380894 5244 380900 5256
rect 380952 5244 380958 5296
rect 390646 5244 390652 5296
rect 390704 5284 390710 5296
rect 430666 5284 430672 5296
rect 390704 5256 430672 5284
rect 390704 5244 390710 5256
rect 430666 5244 430672 5256
rect 430724 5244 430730 5296
rect 21910 5176 21916 5228
rect 21968 5216 21974 5228
rect 240226 5216 240232 5228
rect 21968 5188 240232 5216
rect 21968 5176 21974 5188
rect 240226 5176 240232 5188
rect 240284 5176 240290 5228
rect 251450 5176 251456 5228
rect 251508 5216 251514 5228
rect 358814 5216 358820 5228
rect 251508 5188 358820 5216
rect 251508 5176 251514 5188
rect 358814 5176 358820 5188
rect 358872 5176 358878 5228
rect 387058 5176 387064 5228
rect 387116 5216 387122 5228
rect 427906 5216 427912 5228
rect 387116 5188 427912 5216
rect 387116 5176 387122 5188
rect 427906 5176 427912 5188
rect 427964 5176 427970 5228
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 237466 5148 237472 5160
rect 17368 5120 237472 5148
rect 17368 5108 17374 5120
rect 237466 5108 237472 5120
rect 237524 5108 237530 5160
rect 247954 5108 247960 5160
rect 248012 5148 248018 5160
rect 356422 5148 356428 5160
rect 248012 5120 356428 5148
rect 248012 5108 248018 5120
rect 356422 5108 356428 5120
rect 356480 5108 356486 5160
rect 383562 5108 383568 5160
rect 383620 5148 383626 5160
rect 426710 5148 426716 5160
rect 383620 5120 426716 5148
rect 383620 5108 383626 5120
rect 426710 5108 426716 5120
rect 426768 5108 426774 5160
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 236086 5080 236092 5092
rect 12492 5052 236092 5080
rect 12492 5040 12498 5052
rect 236086 5040 236092 5052
rect 236144 5040 236150 5092
rect 244366 5040 244372 5092
rect 244424 5080 244430 5092
rect 354674 5080 354680 5092
rect 244424 5052 354680 5080
rect 244424 5040 244430 5052
rect 354674 5040 354680 5052
rect 354732 5040 354738 5092
rect 376386 5040 376392 5092
rect 376444 5080 376450 5092
rect 422294 5080 422300 5092
rect 376444 5052 422300 5080
rect 376444 5040 376450 5052
rect 422294 5040 422300 5052
rect 422352 5040 422358 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 233234 5012 233240 5024
rect 7708 4984 233240 5012
rect 7708 4972 7714 4984
rect 233234 4972 233240 4984
rect 233292 4972 233298 5024
rect 240778 4972 240784 5024
rect 240836 5012 240842 5024
rect 353294 5012 353300 5024
rect 240836 4984 353300 5012
rect 240836 4972 240842 4984
rect 353294 4972 353300 4984
rect 353352 4972 353358 5024
rect 365714 4972 365720 5024
rect 365772 5012 365778 5024
rect 416958 5012 416964 5024
rect 365772 4984 416964 5012
rect 365772 4972 365778 4984
rect 416958 4972 416964 4984
rect 417016 4972 417022 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 230474 4944 230480 4956
rect 2924 4916 230480 4944
rect 2924 4904 2930 4916
rect 230474 4904 230480 4916
rect 230532 4904 230538 4956
rect 237190 4904 237196 4956
rect 237248 4944 237254 4956
rect 350534 4944 350540 4956
rect 237248 4916 350540 4944
rect 237248 4904 237254 4916
rect 350534 4904 350540 4916
rect 350592 4904 350598 4956
rect 358538 4904 358544 4956
rect 358596 4944 358602 4956
rect 414106 4944 414112 4956
rect 358596 4916 414112 4944
rect 358596 4904 358602 4916
rect 414106 4904 414112 4916
rect 414164 4904 414170 4956
rect 503530 4904 503536 4956
rect 503588 4944 503594 4956
rect 529658 4944 529664 4956
rect 503588 4916 529664 4944
rect 503588 4904 503594 4916
rect 529658 4904 529664 4916
rect 529716 4904 529722 4956
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 229094 4876 229100 4888
rect 624 4848 229100 4876
rect 624 4836 630 4848
rect 229094 4836 229100 4848
rect 229152 4836 229158 4888
rect 230106 4836 230112 4888
rect 230164 4876 230170 4888
rect 347774 4876 347780 4888
rect 230164 4848 347780 4876
rect 230164 4836 230170 4848
rect 347774 4836 347780 4848
rect 347832 4836 347838 4888
rect 347866 4836 347872 4888
rect 347924 4876 347930 4888
rect 408494 4876 408500 4888
rect 347924 4848 408500 4876
rect 347924 4836 347930 4848
rect 408494 4836 408500 4848
rect 408552 4836 408558 4888
rect 509142 4836 509148 4888
rect 509200 4876 509206 4888
rect 540514 4876 540520 4888
rect 509200 4848 540520 4876
rect 509200 4836 509206 4848
rect 540514 4836 540520 4848
rect 540572 4836 540578 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 230566 4808 230572 4820
rect 1728 4780 230572 4808
rect 1728 4768 1734 4780
rect 230566 4768 230572 4780
rect 230624 4768 230630 4820
rect 233694 4768 233700 4820
rect 233752 4808 233758 4820
rect 349154 4808 349160 4820
rect 233752 4780 349160 4808
rect 233752 4768 233758 4780
rect 349154 4768 349160 4780
rect 349212 4768 349218 4820
rect 351362 4768 351368 4820
rect 351420 4808 351426 4820
rect 410058 4808 410064 4820
rect 351420 4780 410064 4808
rect 351420 4768 351426 4780
rect 410058 4768 410064 4780
rect 410116 4768 410122 4820
rect 506290 4768 506296 4820
rect 506348 4808 506354 4820
rect 536926 4808 536932 4820
rect 506348 4780 536932 4808
rect 506348 4768 506354 4780
rect 536926 4768 536932 4780
rect 536984 4768 536990 4820
rect 215846 4700 215852 4752
rect 215904 4740 215910 4752
rect 339494 4740 339500 4752
rect 215904 4712 339500 4740
rect 215904 4700 215910 4712
rect 339494 4700 339500 4712
rect 339552 4700 339558 4752
rect 340690 4700 340696 4752
rect 340748 4740 340754 4752
rect 404538 4740 404544 4752
rect 340748 4712 404544 4740
rect 340748 4700 340754 4712
rect 404538 4700 404544 4712
rect 404596 4700 404602 4752
rect 404906 4700 404912 4752
rect 404964 4740 404970 4752
rect 437750 4740 437756 4752
rect 404964 4712 437756 4740
rect 404964 4700 404970 4712
rect 437750 4700 437756 4712
rect 437808 4700 437814 4752
rect 222930 4632 222936 4684
rect 222988 4672 222994 4684
rect 343634 4672 343640 4684
rect 222988 4644 343640 4672
rect 222988 4632 222994 4644
rect 343634 4632 343640 4644
rect 343692 4632 343698 4684
rect 344278 4632 344284 4684
rect 344336 4672 344342 4684
rect 405918 4672 405924 4684
rect 344336 4644 405924 4672
rect 344336 4632 344342 4644
rect 405918 4632 405924 4644
rect 405976 4632 405982 4684
rect 226518 4564 226524 4616
rect 226576 4604 226582 4616
rect 345014 4604 345020 4616
rect 226576 4576 345020 4604
rect 226576 4564 226582 4576
rect 345014 4564 345020 4576
rect 345072 4564 345078 4616
rect 356054 4564 356060 4616
rect 356112 4604 356118 4616
rect 362954 4604 362960 4616
rect 356112 4576 362960 4604
rect 356112 4564 356118 4576
rect 362954 4564 362960 4576
rect 363012 4564 363018 4616
rect 208670 4496 208676 4548
rect 208728 4536 208734 4548
rect 283558 4536 283564 4548
rect 208728 4508 283564 4536
rect 208728 4496 208734 4508
rect 283558 4496 283564 4508
rect 283616 4496 283622 4548
rect 319254 4496 319260 4548
rect 319312 4536 319318 4548
rect 393498 4536 393504 4548
rect 319312 4508 393504 4536
rect 319312 4496 319318 4508
rect 393498 4496 393504 4508
rect 393556 4496 393562 4548
rect 212258 4428 212264 4480
rect 212316 4468 212322 4480
rect 284938 4468 284944 4480
rect 212316 4440 284944 4468
rect 212316 4428 212322 4440
rect 284938 4428 284944 4440
rect 284996 4428 285002 4480
rect 322842 4428 322848 4480
rect 322900 4468 322906 4480
rect 394878 4468 394884 4480
rect 322900 4440 394884 4468
rect 322900 4428 322906 4440
rect 394878 4428 394884 4440
rect 394936 4428 394942 4480
rect 326430 4360 326436 4412
rect 326488 4400 326494 4412
rect 397454 4400 397460 4412
rect 326488 4372 397460 4400
rect 326488 4360 326494 4372
rect 397454 4360 397460 4372
rect 397512 4360 397518 4412
rect 330018 4292 330024 4344
rect 330076 4332 330082 4344
rect 399018 4332 399024 4344
rect 330076 4304 399024 4332
rect 330076 4292 330082 4304
rect 399018 4292 399024 4304
rect 399076 4292 399082 4344
rect 403253 4335 403311 4341
rect 403253 4301 403265 4335
rect 403299 4332 403311 4335
rect 408405 4335 408463 4341
rect 408405 4332 408417 4335
rect 403299 4304 408417 4332
rect 403299 4301 403311 4304
rect 403253 4295 403311 4301
rect 408405 4301 408417 4304
rect 408451 4301 408463 4335
rect 408405 4295 408463 4301
rect 333606 4224 333612 4276
rect 333664 4264 333670 4276
rect 400398 4264 400404 4276
rect 333664 4236 400404 4264
rect 333664 4224 333670 4236
rect 400398 4224 400404 4236
rect 400456 4224 400462 4276
rect 408221 4267 408279 4273
rect 408221 4233 408233 4267
rect 408267 4264 408279 4267
rect 408678 4264 408684 4276
rect 408267 4236 408684 4264
rect 408267 4233 408279 4236
rect 408221 4227 408279 4233
rect 408678 4224 408684 4236
rect 408736 4224 408742 4276
rect 124214 4156 124220 4208
rect 124272 4196 124278 4208
rect 125410 4196 125416 4208
rect 124272 4168 125416 4196
rect 124272 4156 124278 4168
rect 125410 4156 125416 4168
rect 125468 4156 125474 4208
rect 140866 4156 140872 4208
rect 140924 4196 140930 4208
rect 142062 4196 142068 4208
rect 140924 4168 142068 4196
rect 140924 4156 140930 4168
rect 142062 4156 142068 4168
rect 142120 4156 142126 4208
rect 150434 4156 150440 4208
rect 150492 4196 150498 4208
rect 151630 4196 151636 4208
rect 150492 4168 151636 4196
rect 150492 4156 150498 4168
rect 151630 4156 151636 4168
rect 151688 4156 151694 4208
rect 158714 4156 158720 4208
rect 158772 4196 158778 4208
rect 159910 4196 159916 4208
rect 158772 4168 159916 4196
rect 158772 4156 158778 4168
rect 159910 4156 159916 4168
rect 159968 4156 159974 4208
rect 209866 4156 209872 4208
rect 209924 4196 209930 4208
rect 211062 4196 211068 4208
rect 209924 4168 211068 4196
rect 209924 4156 209930 4168
rect 211062 4156 211068 4168
rect 211120 4156 211126 4208
rect 314654 4196 314660 4208
rect 314488 4168 314660 4196
rect 42150 4088 42156 4140
rect 42208 4128 42214 4140
rect 50338 4128 50344 4140
rect 42208 4100 50344 4128
rect 42208 4088 42214 4100
rect 50338 4088 50344 4100
rect 50396 4088 50402 4140
rect 57606 4088 57612 4140
rect 57664 4128 57670 4140
rect 255958 4128 255964 4140
rect 57664 4100 255964 4128
rect 57664 4088 57670 4100
rect 255958 4088 255964 4100
rect 256016 4088 256022 4140
rect 275278 4088 275284 4140
rect 275336 4128 275342 4140
rect 276658 4128 276664 4140
rect 275336 4100 276664 4128
rect 275336 4088 275342 4100
rect 276658 4088 276664 4100
rect 276716 4088 276722 4140
rect 278866 4088 278872 4140
rect 278924 4128 278930 4140
rect 280062 4128 280068 4140
rect 278924 4100 280068 4128
rect 278924 4088 278930 4100
rect 280062 4088 280068 4100
rect 280120 4088 280126 4140
rect 280157 4131 280215 4137
rect 280157 4097 280169 4131
rect 280203 4128 280215 4131
rect 314488 4128 314516 4168
rect 314654 4156 314660 4168
rect 314712 4156 314718 4208
rect 337102 4156 337108 4208
rect 337160 4196 337166 4208
rect 403066 4196 403072 4208
rect 337160 4168 403072 4196
rect 337160 4156 337166 4168
rect 403066 4156 403072 4168
rect 403124 4156 403130 4208
rect 403345 4199 403403 4205
rect 403345 4165 403357 4199
rect 403391 4196 403403 4199
rect 404998 4196 405004 4208
rect 403391 4168 405004 4196
rect 403391 4165 403403 4168
rect 403345 4159 403403 4165
rect 404998 4156 405004 4168
rect 405056 4156 405062 4208
rect 408313 4199 408371 4205
rect 408313 4165 408325 4199
rect 408359 4196 408371 4199
rect 408359 4168 408540 4196
rect 408359 4165 408371 4168
rect 408313 4159 408371 4165
rect 280203 4100 314516 4128
rect 280203 4097 280215 4100
rect 280157 4091 280215 4097
rect 314562 4088 314568 4140
rect 314620 4128 314626 4140
rect 316678 4128 316684 4140
rect 314620 4100 316684 4128
rect 314620 4088 314626 4100
rect 316678 4088 316684 4100
rect 316736 4088 316742 4140
rect 321646 4088 321652 4140
rect 321704 4128 321710 4140
rect 322750 4128 322756 4140
rect 321704 4100 322756 4128
rect 321704 4088 321710 4100
rect 322750 4088 322756 4100
rect 322808 4088 322814 4140
rect 331214 4088 331220 4140
rect 331272 4128 331278 4140
rect 332502 4128 332508 4140
rect 331272 4100 332508 4128
rect 331272 4088 331278 4100
rect 332502 4088 332508 4100
rect 332560 4088 332566 4140
rect 346670 4088 346676 4140
rect 346728 4128 346734 4140
rect 391201 4131 391259 4137
rect 391201 4128 391213 4131
rect 346728 4100 391213 4128
rect 346728 4088 346734 4100
rect 391201 4097 391213 4100
rect 391247 4097 391259 4131
rect 391201 4091 391259 4097
rect 393869 4131 393927 4137
rect 393869 4097 393881 4131
rect 393915 4128 393927 4131
rect 393915 4100 400168 4128
rect 393915 4097 393927 4100
rect 393869 4091 393927 4097
rect 50522 4020 50528 4072
rect 50580 4060 50586 4072
rect 253198 4060 253204 4072
rect 50580 4032 253204 4060
rect 50580 4020 50586 4032
rect 253198 4020 253204 4032
rect 253256 4020 253262 4072
rect 262214 4020 262220 4072
rect 262272 4060 262278 4072
rect 322658 4060 322664 4072
rect 262272 4032 322664 4060
rect 262272 4020 262278 4032
rect 322658 4020 322664 4032
rect 322716 4020 322722 4072
rect 339494 4020 339500 4072
rect 339552 4060 339558 4072
rect 392949 4063 393007 4069
rect 392949 4060 392961 4063
rect 339552 4032 392961 4060
rect 339552 4020 339558 4032
rect 392949 4029 392961 4032
rect 392995 4029 393007 4063
rect 392949 4023 393007 4029
rect 393961 4063 394019 4069
rect 393961 4029 393973 4063
rect 394007 4060 394019 4063
rect 400033 4063 400091 4069
rect 400033 4060 400045 4063
rect 394007 4032 400045 4060
rect 394007 4029 394019 4032
rect 393961 4023 394019 4029
rect 400033 4029 400045 4032
rect 400079 4029 400091 4063
rect 400140 4060 400168 4100
rect 400214 4088 400220 4140
rect 400272 4128 400278 4140
rect 408402 4128 408408 4140
rect 400272 4100 408408 4128
rect 400272 4088 400278 4100
rect 408402 4088 408408 4100
rect 408460 4088 408466 4140
rect 408512 4128 408540 4168
rect 408586 4156 408592 4208
rect 408644 4196 408650 4208
rect 408644 4168 412680 4196
rect 408644 4156 408650 4168
rect 410518 4128 410524 4140
rect 408512 4100 410524 4128
rect 410518 4088 410524 4100
rect 410576 4088 410582 4140
rect 411898 4128 411904 4140
rect 410628 4100 411904 4128
rect 403526 4060 403532 4072
rect 400140 4032 403532 4060
rect 400033 4023 400091 4029
rect 403526 4020 403532 4032
rect 403584 4020 403590 4072
rect 408497 4063 408555 4069
rect 408497 4060 408509 4063
rect 403636 4032 408509 4060
rect 34974 3952 34980 4004
rect 35032 3992 35038 4004
rect 46198 3992 46204 4004
rect 35032 3964 46204 3992
rect 35032 3952 35038 3964
rect 46198 3952 46204 3964
rect 46256 3952 46262 4004
rect 46934 3952 46940 4004
rect 46992 3992 46998 4004
rect 252738 3992 252744 4004
rect 46992 3964 252744 3992
rect 46992 3952 46998 3964
rect 252738 3952 252744 3964
rect 252796 3952 252802 4004
rect 271690 3952 271696 4004
rect 271748 3992 271754 4004
rect 277949 3995 278007 4001
rect 277949 3992 277961 3995
rect 271748 3964 277961 3992
rect 271748 3952 271754 3964
rect 277949 3961 277961 3964
rect 277995 3961 278007 3995
rect 277949 3955 278007 3961
rect 278041 3995 278099 4001
rect 278041 3961 278053 3995
rect 278087 3992 278099 3995
rect 283466 3992 283472 4004
rect 278087 3964 283472 3992
rect 278087 3961 278099 3964
rect 278041 3955 278099 3961
rect 283466 3952 283472 3964
rect 283524 3952 283530 4004
rect 300302 3952 300308 4004
rect 300360 3992 300366 4004
rect 363598 3992 363604 4004
rect 300360 3964 363604 3992
rect 300360 3952 300366 3964
rect 363598 3952 363604 3964
rect 363656 3952 363662 4004
rect 364518 3952 364524 4004
rect 364576 3992 364582 4004
rect 366358 3992 366364 4004
rect 364576 3964 366364 3992
rect 364576 3952 364582 3964
rect 366358 3952 366364 3964
rect 366416 3952 366422 4004
rect 371602 3952 371608 4004
rect 371660 3992 371666 4004
rect 372522 3992 372528 4004
rect 371660 3964 372528 3992
rect 371660 3952 371666 3964
rect 372522 3952 372528 3964
rect 372580 3952 372586 4004
rect 384301 3995 384359 4001
rect 384301 3961 384313 3995
rect 384347 3992 384359 3995
rect 403636 3992 403664 4032
rect 408497 4029 408509 4032
rect 408543 4029 408555 4063
rect 409138 4060 409144 4072
rect 408497 4023 408555 4029
rect 408604 4032 409144 4060
rect 384347 3964 403664 3992
rect 403713 3995 403771 4001
rect 384347 3961 384359 3964
rect 384301 3955 384359 3961
rect 403713 3961 403725 3995
rect 403759 3992 403771 3995
rect 408313 3995 408371 4001
rect 408313 3992 408325 3995
rect 403759 3964 408325 3992
rect 403759 3961 403771 3964
rect 403713 3955 403771 3961
rect 408313 3961 408325 3964
rect 408359 3961 408371 3995
rect 408313 3955 408371 3961
rect 408405 3995 408463 4001
rect 408405 3961 408417 3995
rect 408451 3992 408463 3995
rect 408604 3992 408632 4032
rect 409138 4020 409144 4032
rect 409196 4020 409202 4072
rect 409233 4063 409291 4069
rect 409233 4029 409245 4063
rect 409279 4060 409291 4063
rect 410628 4060 410656 4100
rect 411898 4088 411904 4100
rect 411956 4088 411962 4140
rect 412082 4088 412088 4140
rect 412140 4128 412146 4140
rect 412542 4128 412548 4140
rect 412140 4100 412548 4128
rect 412140 4088 412146 4100
rect 412542 4088 412548 4100
rect 412600 4088 412606 4140
rect 412652 4128 412680 4168
rect 413649 4131 413707 4137
rect 413649 4128 413661 4131
rect 412652 4100 413661 4128
rect 413649 4097 413661 4100
rect 413695 4097 413707 4131
rect 413649 4091 413707 4097
rect 414474 4088 414480 4140
rect 414532 4128 414538 4140
rect 416038 4128 416044 4140
rect 414532 4100 416044 4128
rect 414532 4088 414538 4100
rect 416038 4088 416044 4100
rect 416096 4088 416102 4140
rect 416133 4131 416191 4137
rect 416133 4097 416145 4131
rect 416179 4128 416191 4131
rect 419077 4131 419135 4137
rect 419077 4128 419089 4131
rect 416179 4100 419089 4128
rect 416179 4097 416191 4100
rect 416133 4091 416191 4097
rect 419077 4097 419089 4100
rect 419123 4097 419135 4131
rect 419077 4091 419135 4097
rect 419166 4088 419172 4140
rect 419224 4128 419230 4140
rect 420178 4128 420184 4140
rect 419224 4100 420184 4128
rect 419224 4088 419230 4100
rect 420178 4088 420184 4100
rect 420236 4088 420242 4140
rect 420362 4088 420368 4140
rect 420420 4128 420426 4140
rect 420822 4128 420828 4140
rect 420420 4100 420828 4128
rect 420420 4088 420426 4100
rect 420822 4088 420828 4100
rect 420880 4088 420886 4140
rect 422754 4088 422760 4140
rect 422812 4128 422818 4140
rect 423582 4128 423588 4140
rect 422812 4100 423588 4128
rect 422812 4088 422818 4100
rect 423582 4088 423588 4100
rect 423640 4088 423646 4140
rect 423950 4088 423956 4140
rect 424008 4128 424014 4140
rect 424962 4128 424968 4140
rect 424008 4100 424968 4128
rect 424008 4088 424014 4100
rect 424962 4088 424968 4100
rect 425020 4088 425026 4140
rect 425057 4131 425115 4137
rect 425057 4097 425069 4131
rect 425103 4128 425115 4131
rect 429286 4128 429292 4140
rect 425103 4100 429292 4128
rect 425103 4097 425115 4100
rect 425057 4091 425115 4097
rect 429286 4088 429292 4100
rect 429344 4088 429350 4140
rect 429930 4088 429936 4140
rect 429988 4128 429994 4140
rect 430482 4128 430488 4140
rect 429988 4100 430488 4128
rect 429988 4088 429994 4100
rect 430482 4088 430488 4100
rect 430540 4088 430546 4140
rect 431126 4088 431132 4140
rect 431184 4128 431190 4140
rect 431862 4128 431868 4140
rect 431184 4100 431868 4128
rect 431184 4088 431190 4100
rect 431862 4088 431868 4100
rect 431920 4088 431926 4140
rect 433518 4088 433524 4140
rect 433576 4128 433582 4140
rect 434622 4128 434628 4140
rect 433576 4100 434628 4128
rect 433576 4088 433582 4100
rect 434622 4088 434628 4100
rect 434680 4088 434686 4140
rect 437014 4088 437020 4140
rect 437072 4128 437078 4140
rect 442350 4128 442356 4140
rect 437072 4100 442356 4128
rect 437072 4088 437078 4100
rect 442350 4088 442356 4100
rect 442408 4088 442414 4140
rect 451274 4088 451280 4140
rect 451332 4128 451338 4140
rect 453298 4128 453304 4140
rect 451332 4100 453304 4128
rect 451332 4088 451338 4100
rect 453298 4088 453304 4100
rect 453356 4088 453362 4140
rect 454862 4088 454868 4140
rect 454920 4128 454926 4140
rect 456058 4128 456064 4140
rect 454920 4100 456064 4128
rect 454920 4088 454926 4100
rect 456058 4088 456064 4100
rect 456116 4088 456122 4140
rect 469122 4088 469128 4140
rect 469180 4128 469186 4140
rect 469858 4128 469864 4140
rect 469180 4100 469864 4128
rect 469180 4088 469186 4100
rect 469858 4088 469864 4100
rect 469916 4088 469922 4140
rect 472158 4088 472164 4140
rect 472216 4128 472222 4140
rect 472710 4128 472716 4140
rect 472216 4100 472716 4128
rect 472216 4088 472222 4100
rect 472710 4088 472716 4100
rect 472768 4088 472774 4140
rect 473354 4088 473360 4140
rect 473412 4128 473418 4140
rect 473906 4128 473912 4140
rect 473412 4100 473912 4128
rect 473412 4088 473418 4100
rect 473906 4088 473912 4100
rect 473964 4088 473970 4140
rect 474642 4088 474648 4140
rect 474700 4128 474706 4140
rect 475102 4128 475108 4140
rect 474700 4100 475108 4128
rect 474700 4088 474706 4100
rect 475102 4088 475108 4100
rect 475160 4088 475166 4140
rect 493962 4088 493968 4140
rect 494020 4128 494026 4140
rect 511994 4128 512000 4140
rect 494020 4100 512000 4128
rect 494020 4088 494026 4100
rect 511994 4088 512000 4100
rect 512052 4088 512058 4140
rect 518802 4088 518808 4140
rect 518860 4128 518866 4140
rect 559558 4128 559564 4140
rect 518860 4100 559564 4128
rect 518860 4088 518866 4100
rect 559558 4088 559564 4100
rect 559616 4088 559622 4140
rect 409279 4032 410656 4060
rect 409279 4029 409291 4032
rect 409233 4023 409291 4029
rect 410886 4020 410892 4072
rect 410944 4060 410950 4072
rect 413278 4060 413284 4072
rect 410944 4032 413284 4060
rect 410944 4020 410950 4032
rect 413278 4020 413284 4032
rect 413336 4020 413342 4072
rect 413373 4063 413431 4069
rect 413373 4029 413385 4063
rect 413419 4060 413431 4063
rect 438946 4060 438952 4072
rect 413419 4032 438952 4060
rect 413419 4029 413431 4032
rect 413373 4023 413431 4029
rect 438946 4020 438952 4032
rect 439004 4020 439010 4072
rect 440602 4020 440608 4072
rect 440660 4060 440666 4072
rect 445018 4060 445024 4072
rect 440660 4032 445024 4060
rect 440660 4020 440666 4032
rect 445018 4020 445024 4032
rect 445076 4020 445082 4072
rect 492490 4020 492496 4072
rect 492548 4060 492554 4072
rect 509602 4060 509608 4072
rect 492548 4032 509608 4060
rect 492548 4020 492554 4032
rect 509602 4020 509608 4032
rect 509660 4020 509666 4072
rect 520090 4020 520096 4072
rect 520148 4060 520154 4072
rect 561950 4060 561956 4072
rect 520148 4032 561956 4060
rect 520148 4020 520154 4032
rect 561950 4020 561956 4032
rect 562008 4020 562014 4072
rect 408451 3964 408632 3992
rect 408451 3961 408463 3964
rect 408405 3955 408463 3961
rect 408678 3952 408684 4004
rect 408736 3992 408742 4004
rect 418985 3995 419043 4001
rect 418985 3992 418997 3995
rect 408736 3964 418997 3992
rect 408736 3952 408742 3964
rect 418985 3961 418997 3964
rect 419031 3961 419043 3995
rect 418985 3955 419043 3961
rect 419077 3995 419135 4001
rect 419077 3961 419089 3995
rect 419123 3992 419135 3995
rect 420270 3992 420276 4004
rect 419123 3964 420276 3992
rect 419123 3961 419135 3964
rect 419077 3955 419135 3961
rect 420270 3952 420276 3964
rect 420328 3952 420334 4004
rect 421285 3995 421343 4001
rect 421285 3961 421297 3995
rect 421331 3992 421343 3995
rect 424410 3992 424416 4004
rect 421331 3964 424416 3992
rect 421331 3961 421343 3964
rect 421285 3955 421343 3961
rect 424410 3952 424416 3964
rect 424468 3952 424474 4004
rect 427538 3952 427544 4004
rect 427596 3992 427602 4004
rect 432601 3995 432659 4001
rect 432601 3992 432613 3995
rect 427596 3964 432613 3992
rect 427596 3952 427602 3964
rect 432601 3961 432613 3964
rect 432647 3961 432659 3995
rect 448514 3992 448520 4004
rect 432601 3955 432659 3961
rect 432708 3964 448520 3992
rect 45738 3884 45744 3936
rect 45796 3924 45802 3936
rect 251818 3924 251824 3936
rect 45796 3896 251824 3924
rect 45796 3884 45802 3896
rect 251818 3884 251824 3896
rect 251876 3884 251882 3936
rect 258626 3884 258632 3936
rect 258684 3924 258690 3936
rect 322566 3924 322572 3936
rect 258684 3896 322572 3924
rect 258684 3884 258690 3896
rect 322566 3884 322572 3896
rect 322624 3884 322630 3936
rect 325234 3884 325240 3936
rect 325292 3924 325298 3936
rect 391106 3924 391112 3936
rect 325292 3896 391112 3924
rect 325292 3884 325298 3896
rect 391106 3884 391112 3896
rect 391164 3884 391170 3936
rect 391201 3927 391259 3933
rect 391201 3893 391213 3927
rect 391247 3924 391259 3927
rect 400858 3924 400864 3936
rect 391247 3896 400864 3924
rect 391247 3893 391259 3896
rect 391201 3887 391259 3893
rect 400858 3884 400864 3896
rect 400916 3884 400922 3936
rect 408586 3884 408592 3936
rect 408644 3924 408650 3936
rect 423033 3927 423091 3933
rect 423033 3924 423045 3927
rect 408644 3896 423045 3924
rect 408644 3884 408650 3896
rect 423033 3893 423045 3896
rect 423079 3893 423091 3927
rect 423033 3887 423091 3893
rect 425146 3884 425152 3936
rect 425204 3924 425210 3936
rect 432708 3924 432736 3964
rect 448514 3952 448520 3964
rect 448572 3952 448578 4004
rect 458450 3952 458456 4004
rect 458508 3992 458514 4004
rect 464430 3992 464436 4004
rect 458508 3964 464436 3992
rect 458508 3952 458514 3964
rect 464430 3952 464436 3964
rect 464488 3952 464494 4004
rect 493870 3952 493876 4004
rect 493928 3992 493934 4004
rect 513190 3992 513196 4004
rect 493928 3964 513196 3992
rect 493928 3952 493934 3964
rect 513190 3952 513196 3964
rect 513248 3952 513254 4004
rect 520182 3952 520188 4004
rect 520240 3992 520246 4004
rect 564342 3992 564348 4004
rect 520240 3964 564348 3992
rect 520240 3952 520246 3964
rect 564342 3952 564348 3964
rect 564400 3952 564406 4004
rect 565078 3952 565084 4004
rect 565136 3992 565142 4004
rect 579798 3992 579804 4004
rect 565136 3964 579804 3992
rect 565136 3952 565142 3964
rect 579798 3952 579804 3964
rect 579856 3952 579862 4004
rect 425204 3896 432736 3924
rect 432785 3927 432843 3933
rect 425204 3884 425210 3896
rect 432785 3893 432797 3927
rect 432831 3924 432843 3927
rect 442258 3924 442264 3936
rect 432831 3896 442264 3924
rect 432831 3893 432843 3896
rect 432785 3887 432843 3893
rect 442258 3884 442264 3896
rect 442316 3884 442322 3936
rect 496078 3884 496084 3936
rect 496136 3924 496142 3936
rect 496136 3896 509832 3924
rect 496136 3884 496142 3896
rect 39758 3816 39764 3868
rect 39816 3856 39822 3868
rect 249794 3856 249800 3868
rect 39816 3828 249800 3856
rect 39816 3816 39822 3828
rect 249794 3816 249800 3828
rect 249852 3816 249858 3868
rect 255038 3816 255044 3868
rect 255096 3856 255102 3868
rect 255096 3828 316724 3856
rect 255096 3816 255102 3828
rect 38562 3748 38568 3800
rect 38620 3788 38626 3800
rect 248414 3788 248420 3800
rect 38620 3760 248420 3788
rect 38620 3748 38626 3760
rect 248414 3748 248420 3760
rect 248472 3748 248478 3800
rect 272886 3748 272892 3800
rect 272944 3788 272950 3800
rect 316586 3788 316592 3800
rect 272944 3760 316592 3788
rect 272944 3748 272950 3760
rect 316586 3748 316592 3760
rect 316644 3748 316650 3800
rect 32674 3680 32680 3732
rect 32732 3720 32738 3732
rect 245654 3720 245660 3732
rect 32732 3692 245660 3720
rect 32732 3680 32738 3692
rect 245654 3680 245660 3692
rect 245712 3680 245718 3732
rect 264606 3680 264612 3732
rect 264664 3720 264670 3732
rect 278041 3723 278099 3729
rect 278041 3720 278053 3723
rect 264664 3692 278053 3720
rect 264664 3680 264670 3692
rect 278041 3689 278053 3692
rect 278087 3689 278099 3723
rect 278041 3683 278099 3689
rect 278133 3723 278191 3729
rect 278133 3689 278145 3723
rect 278179 3720 278191 3723
rect 287698 3720 287704 3732
rect 278179 3692 287704 3720
rect 278179 3689 278191 3692
rect 278133 3683 278191 3689
rect 287698 3680 287704 3692
rect 287756 3680 287762 3732
rect 299106 3680 299112 3732
rect 299164 3720 299170 3732
rect 300946 3720 300952 3732
rect 299164 3692 300952 3720
rect 299164 3680 299170 3692
rect 300946 3680 300952 3692
rect 301004 3680 301010 3732
rect 307386 3680 307392 3732
rect 307444 3720 307450 3732
rect 309778 3720 309784 3732
rect 307444 3692 309784 3720
rect 307444 3680 307450 3692
rect 309778 3680 309784 3692
rect 309836 3680 309842 3732
rect 316696 3720 316724 3828
rect 316954 3816 316960 3868
rect 317012 3856 317018 3868
rect 327074 3856 327080 3868
rect 317012 3828 327080 3856
rect 317012 3816 317018 3828
rect 327074 3816 327080 3828
rect 327132 3816 327138 3868
rect 332410 3816 332416 3868
rect 332468 3856 332474 3868
rect 392949 3859 393007 3865
rect 332468 3828 392256 3856
rect 332468 3816 332474 3828
rect 318058 3748 318064 3800
rect 318116 3788 318122 3800
rect 389818 3788 389824 3800
rect 318116 3760 389824 3788
rect 318116 3748 318122 3760
rect 389818 3748 389824 3760
rect 389876 3748 389882 3800
rect 392228 3788 392256 3828
rect 392949 3825 392961 3859
rect 392995 3856 393007 3859
rect 396718 3856 396724 3868
rect 392995 3828 396724 3856
rect 392995 3825 393007 3828
rect 392949 3819 393007 3825
rect 396718 3816 396724 3828
rect 396776 3816 396782 3868
rect 400033 3859 400091 3865
rect 400033 3825 400045 3859
rect 400079 3856 400091 3859
rect 403345 3859 403403 3865
rect 403345 3856 403357 3859
rect 400079 3828 403357 3856
rect 400079 3825 400091 3828
rect 400033 3819 400091 3825
rect 403345 3825 403357 3828
rect 403391 3825 403403 3859
rect 403345 3819 403403 3825
rect 403710 3816 403716 3868
rect 403768 3856 403774 3868
rect 437658 3856 437664 3868
rect 403768 3828 437664 3856
rect 403768 3816 403774 3828
rect 437658 3816 437664 3828
rect 437716 3816 437722 3868
rect 448974 3816 448980 3868
rect 449032 3856 449038 3868
rect 453390 3856 453396 3868
rect 449032 3828 453396 3856
rect 449032 3816 449038 3828
rect 453390 3816 453396 3828
rect 453448 3816 453454 3868
rect 482922 3816 482928 3868
rect 482980 3856 482986 3868
rect 490558 3856 490564 3868
rect 482980 3828 490564 3856
rect 482980 3816 482986 3828
rect 490558 3816 490564 3828
rect 490616 3816 490622 3868
rect 496722 3816 496728 3868
rect 496780 3856 496786 3868
rect 509697 3859 509755 3865
rect 509697 3856 509709 3859
rect 496780 3828 509709 3856
rect 496780 3816 496786 3828
rect 509697 3825 509709 3828
rect 509743 3825 509755 3859
rect 509804 3856 509832 3896
rect 509878 3884 509884 3936
rect 509936 3924 509942 3936
rect 520274 3924 520280 3936
rect 509936 3896 520280 3924
rect 509936 3884 509942 3896
rect 520274 3884 520280 3896
rect 520332 3884 520338 3936
rect 521562 3884 521568 3936
rect 521620 3924 521626 3936
rect 566734 3924 566740 3936
rect 521620 3896 566740 3924
rect 521620 3884 521626 3896
rect 566734 3884 566740 3896
rect 566792 3884 566798 3936
rect 515582 3856 515588 3868
rect 509804 3828 515588 3856
rect 509697 3819 509755 3825
rect 515582 3816 515588 3828
rect 515640 3816 515646 3868
rect 516778 3816 516784 3868
rect 516836 3856 516842 3868
rect 523037 3859 523095 3865
rect 516836 3828 522896 3856
rect 516836 3816 516842 3828
rect 395338 3788 395344 3800
rect 392228 3760 395344 3788
rect 395338 3748 395344 3760
rect 395396 3748 395402 3800
rect 399018 3748 399024 3800
rect 399076 3788 399082 3800
rect 434806 3788 434812 3800
rect 399076 3760 434812 3788
rect 399076 3748 399082 3760
rect 434806 3748 434812 3760
rect 434864 3748 434870 3800
rect 438210 3748 438216 3800
rect 438268 3788 438274 3800
rect 447778 3788 447784 3800
rect 438268 3760 447784 3788
rect 438268 3748 438274 3760
rect 447778 3748 447784 3760
rect 447836 3748 447842 3800
rect 455598 3788 455604 3800
rect 447888 3760 455604 3788
rect 325326 3720 325332 3732
rect 316696 3692 325332 3720
rect 325326 3680 325332 3692
rect 325384 3680 325390 3732
rect 352558 3680 352564 3732
rect 352616 3720 352622 3732
rect 353202 3720 353208 3732
rect 352616 3692 353208 3720
rect 352616 3680 352622 3692
rect 353202 3680 353208 3692
rect 353260 3680 353266 3732
rect 374641 3723 374699 3729
rect 374641 3689 374653 3723
rect 374687 3720 374699 3723
rect 384301 3723 384359 3729
rect 384301 3720 384313 3723
rect 374687 3692 384313 3720
rect 374687 3689 374699 3692
rect 374641 3683 374699 3689
rect 384301 3689 384313 3692
rect 384347 3689 384359 3723
rect 384301 3683 384359 3689
rect 385862 3680 385868 3732
rect 385920 3720 385926 3732
rect 403253 3723 403311 3729
rect 403253 3720 403265 3723
rect 385920 3692 403265 3720
rect 385920 3680 385926 3692
rect 403253 3689 403265 3692
rect 403299 3689 403311 3723
rect 403253 3683 403311 3689
rect 403713 3723 403771 3729
rect 403713 3689 403725 3723
rect 403759 3720 403771 3723
rect 408221 3723 408279 3729
rect 408221 3720 408233 3723
rect 403759 3692 408233 3720
rect 403759 3689 403771 3692
rect 403713 3683 403771 3689
rect 408221 3689 408233 3692
rect 408267 3689 408279 3723
rect 408221 3683 408279 3689
rect 418065 3723 418123 3729
rect 418065 3689 418077 3723
rect 418111 3720 418123 3723
rect 418111 3692 422984 3720
rect 418111 3689 418123 3692
rect 418065 3683 418123 3689
rect 25498 3612 25504 3664
rect 25556 3652 25562 3664
rect 238205 3655 238263 3661
rect 238205 3652 238217 3655
rect 25556 3624 238217 3652
rect 25556 3612 25562 3624
rect 238205 3621 238217 3624
rect 238251 3621 238263 3655
rect 238205 3615 238263 3621
rect 239582 3612 239588 3664
rect 239640 3652 239646 3664
rect 240042 3652 240048 3664
rect 239640 3624 240048 3652
rect 239640 3612 239646 3624
rect 240042 3612 240048 3624
rect 240100 3612 240106 3664
rect 243170 3612 243176 3664
rect 243228 3652 243234 3664
rect 244182 3652 244188 3664
rect 243228 3624 244188 3652
rect 243228 3612 243234 3624
rect 244182 3612 244188 3624
rect 244240 3612 244246 3664
rect 269298 3612 269304 3664
rect 269356 3652 269362 3664
rect 289814 3652 289820 3664
rect 269356 3624 289820 3652
rect 269356 3612 269362 3624
rect 289814 3612 289820 3624
rect 289872 3612 289878 3664
rect 291930 3612 291936 3664
rect 291988 3652 291994 3664
rect 299658 3652 299664 3664
rect 291988 3624 299664 3652
rect 291988 3612 291994 3624
rect 299658 3612 299664 3624
rect 299716 3612 299722 3664
rect 303798 3612 303804 3664
rect 303856 3652 303862 3664
rect 382918 3652 382924 3664
rect 303856 3624 382924 3652
rect 303856 3612 303862 3624
rect 382918 3612 382924 3624
rect 382976 3612 382982 3664
rect 388254 3612 388260 3664
rect 388312 3652 388318 3664
rect 389082 3652 389088 3664
rect 388312 3624 389088 3652
rect 388312 3612 388318 3624
rect 389082 3612 389088 3624
rect 389140 3612 389146 3664
rect 391842 3612 391848 3664
rect 391900 3652 391906 3664
rect 408310 3652 408316 3664
rect 391900 3624 408316 3652
rect 391900 3612 391906 3624
rect 408310 3612 408316 3624
rect 408368 3612 408374 3664
rect 408405 3655 408463 3661
rect 408405 3621 408417 3655
rect 408451 3652 408463 3655
rect 408494 3652 408500 3664
rect 408451 3624 408500 3652
rect 408451 3621 408463 3624
rect 408405 3615 408463 3621
rect 408494 3612 408500 3624
rect 408552 3612 408558 3664
rect 408586 3612 408592 3664
rect 408644 3652 408650 3664
rect 422849 3655 422907 3661
rect 422849 3652 422861 3655
rect 408644 3624 422861 3652
rect 408644 3612 408650 3624
rect 422849 3621 422861 3624
rect 422895 3621 422907 3655
rect 422849 3615 422907 3621
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 19242 3584 19248 3596
rect 18380 3556 19248 3584
rect 18380 3544 18386 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 24118 3584 24124 3596
rect 19576 3556 24124 3584
rect 19576 3544 19582 3556
rect 24118 3544 24124 3556
rect 24176 3544 24182 3596
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 241514 3584 241520 3596
rect 24360 3556 241520 3584
rect 24360 3544 24366 3556
rect 241514 3544 241520 3556
rect 241572 3544 241578 3596
rect 278041 3587 278099 3593
rect 278041 3553 278053 3587
rect 278087 3584 278099 3587
rect 278087 3556 287744 3584
rect 278087 3553 278099 3556
rect 278041 3547 278099 3553
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 236362 3516 236368 3528
rect 14884 3488 236368 3516
rect 14884 3476 14890 3488
rect 236362 3476 236368 3488
rect 236420 3476 236426 3528
rect 238205 3519 238263 3525
rect 238205 3485 238217 3519
rect 238251 3516 238263 3519
rect 241790 3516 241796 3528
rect 238251 3488 241796 3516
rect 238251 3485 238263 3488
rect 238205 3479 238263 3485
rect 241790 3476 241796 3488
rect 241848 3476 241854 3528
rect 265802 3476 265808 3528
rect 265860 3516 265866 3528
rect 287606 3516 287612 3528
rect 265860 3488 287612 3516
rect 265860 3476 265866 3488
rect 287606 3476 287612 3488
rect 287664 3476 287670 3528
rect 287716 3516 287744 3556
rect 289538 3544 289544 3596
rect 289596 3584 289602 3596
rect 292577 3587 292635 3593
rect 292577 3584 292589 3587
rect 289596 3556 292589 3584
rect 289596 3544 289602 3556
rect 292577 3553 292589 3556
rect 292623 3553 292635 3587
rect 292577 3547 292635 3553
rect 296714 3544 296720 3596
rect 296772 3584 296778 3596
rect 381538 3584 381544 3596
rect 296772 3556 381544 3584
rect 296772 3544 296778 3556
rect 381538 3544 381544 3556
rect 381596 3544 381602 3596
rect 389450 3544 389456 3596
rect 389508 3584 389514 3596
rect 422956 3584 422984 3692
rect 434530 3680 434536 3732
rect 434588 3720 434594 3732
rect 446490 3720 446496 3732
rect 434588 3692 446496 3720
rect 434588 3680 434594 3692
rect 446490 3680 446496 3692
rect 446548 3680 446554 3732
rect 447689 3723 447747 3729
rect 447689 3689 447701 3723
rect 447735 3720 447747 3723
rect 447888 3720 447916 3760
rect 455598 3748 455604 3760
rect 455656 3748 455662 3800
rect 489178 3748 489184 3800
rect 489236 3788 489242 3800
rect 497734 3788 497740 3800
rect 489236 3760 497740 3788
rect 489236 3748 489242 3760
rect 497734 3748 497740 3760
rect 497792 3748 497798 3800
rect 498838 3748 498844 3800
rect 498896 3788 498902 3800
rect 519078 3788 519084 3800
rect 498896 3760 519084 3788
rect 498896 3748 498902 3760
rect 519078 3748 519084 3760
rect 519136 3748 519142 3800
rect 447735 3692 447916 3720
rect 447735 3689 447747 3692
rect 447689 3683 447747 3689
rect 450170 3680 450176 3732
rect 450228 3720 450234 3732
rect 451182 3720 451188 3732
rect 450228 3692 451188 3720
rect 450228 3680 450234 3692
rect 451182 3680 451188 3692
rect 451240 3680 451246 3732
rect 457254 3680 457260 3732
rect 457312 3720 457318 3732
rect 465350 3720 465356 3732
rect 457312 3692 465356 3720
rect 457312 3680 457318 3692
rect 465350 3680 465356 3692
rect 465408 3680 465414 3732
rect 466822 3680 466828 3732
rect 466880 3720 466886 3732
rect 467742 3720 467748 3732
rect 466880 3692 467748 3720
rect 466880 3680 466886 3692
rect 467742 3680 467748 3692
rect 467800 3680 467806 3732
rect 485682 3680 485688 3732
rect 485740 3720 485746 3732
rect 495342 3720 495348 3732
rect 485740 3692 495348 3720
rect 485740 3680 485746 3692
rect 495342 3680 495348 3692
rect 495400 3680 495406 3732
rect 499482 3680 499488 3732
rect 499540 3720 499546 3732
rect 522666 3720 522672 3732
rect 499540 3692 522672 3720
rect 499540 3680 499546 3692
rect 522666 3680 522672 3692
rect 522724 3680 522730 3732
rect 522868 3720 522896 3828
rect 523037 3825 523049 3859
rect 523083 3856 523095 3859
rect 525058 3856 525064 3868
rect 523083 3828 525064 3856
rect 523083 3825 523095 3828
rect 523037 3819 523095 3825
rect 525058 3816 525064 3828
rect 525116 3816 525122 3868
rect 525610 3816 525616 3868
rect 525668 3856 525674 3868
rect 572622 3856 572628 3868
rect 525668 3828 572628 3856
rect 525668 3816 525674 3828
rect 572622 3816 572628 3828
rect 572680 3816 572686 3868
rect 522942 3748 522948 3800
rect 523000 3788 523006 3800
rect 569034 3788 569040 3800
rect 523000 3760 569040 3788
rect 523000 3748 523006 3760
rect 569034 3748 569040 3760
rect 569092 3748 569098 3800
rect 522868 3692 524000 3720
rect 423033 3655 423091 3661
rect 423033 3621 423045 3655
rect 423079 3652 423091 3655
rect 432598 3652 432604 3664
rect 423079 3624 432604 3652
rect 423079 3621 423091 3624
rect 423033 3615 423091 3621
rect 432598 3612 432604 3624
rect 432656 3612 432662 3664
rect 442994 3612 443000 3664
rect 443052 3652 443058 3664
rect 456886 3652 456892 3664
rect 443052 3624 456892 3652
rect 443052 3612 443058 3624
rect 456886 3612 456892 3624
rect 456944 3612 456950 3664
rect 478782 3612 478788 3664
rect 478840 3652 478846 3664
rect 482278 3652 482284 3664
rect 478840 3624 482284 3652
rect 478840 3612 478846 3624
rect 482278 3612 482284 3624
rect 482336 3612 482342 3664
rect 484210 3612 484216 3664
rect 484268 3652 484274 3664
rect 492950 3652 492956 3664
rect 484268 3624 492956 3652
rect 484268 3612 484274 3624
rect 492950 3612 492956 3624
rect 493008 3612 493014 3664
rect 500770 3612 500776 3664
rect 500828 3652 500834 3664
rect 523037 3655 523095 3661
rect 523037 3652 523049 3655
rect 500828 3624 523049 3652
rect 500828 3612 500834 3624
rect 523037 3621 523049 3624
rect 523083 3621 523095 3655
rect 523037 3615 523095 3621
rect 433334 3584 433340 3596
rect 389508 3556 422892 3584
rect 422956 3556 433340 3584
rect 389508 3544 389514 3556
rect 289906 3516 289912 3528
rect 287716 3488 289912 3516
rect 289906 3476 289912 3488
rect 289964 3476 289970 3528
rect 302145 3519 302203 3525
rect 302145 3485 302157 3519
rect 302191 3516 302203 3519
rect 378410 3516 378416 3528
rect 302191 3488 378416 3516
rect 302191 3485 302203 3488
rect 302145 3479 302203 3485
rect 378410 3476 378416 3488
rect 378468 3476 378474 3528
rect 382366 3476 382372 3528
rect 382424 3516 382430 3528
rect 418893 3519 418951 3525
rect 418893 3516 418905 3519
rect 382424 3488 418905 3516
rect 382424 3476 382430 3488
rect 418893 3485 418905 3488
rect 418939 3485 418951 3519
rect 418893 3479 418951 3485
rect 418985 3519 419043 3525
rect 418985 3485 418997 3519
rect 419031 3516 419043 3519
rect 421285 3519 421343 3525
rect 421285 3516 421297 3519
rect 419031 3488 421297 3516
rect 419031 3485 419043 3488
rect 418985 3479 419043 3485
rect 421285 3485 421297 3488
rect 421331 3485 421343 3519
rect 422864 3516 422892 3556
rect 433334 3544 433340 3556
rect 433392 3544 433398 3596
rect 439406 3544 439412 3596
rect 439464 3584 439470 3596
rect 447689 3587 447747 3593
rect 447689 3584 447701 3587
rect 439464 3556 447701 3584
rect 439464 3544 439470 3556
rect 447689 3553 447701 3556
rect 447735 3553 447747 3587
rect 447689 3547 447747 3553
rect 447778 3544 447784 3596
rect 447836 3584 447842 3596
rect 448422 3584 448428 3596
rect 447836 3556 448428 3584
rect 447836 3544 447842 3556
rect 448422 3544 448428 3556
rect 448480 3544 448486 3596
rect 467926 3544 467932 3596
rect 467984 3584 467990 3596
rect 470778 3584 470784 3596
rect 467984 3556 470784 3584
rect 467984 3544 467990 3556
rect 470778 3544 470784 3556
rect 470836 3544 470842 3596
rect 484302 3544 484308 3596
rect 484360 3584 484366 3596
rect 494146 3584 494152 3596
rect 484360 3556 494152 3584
rect 484360 3544 484366 3556
rect 494146 3544 494152 3556
rect 494204 3544 494210 3596
rect 499390 3544 499396 3596
rect 499448 3584 499454 3596
rect 523862 3584 523868 3596
rect 499448 3556 523868 3584
rect 499448 3544 499454 3556
rect 523862 3544 523868 3556
rect 523920 3544 523926 3596
rect 523972 3584 524000 3692
rect 524322 3680 524328 3732
rect 524380 3720 524386 3732
rect 571426 3720 571432 3732
rect 524380 3692 571432 3720
rect 524380 3680 524386 3692
rect 571426 3680 571432 3692
rect 571484 3680 571490 3732
rect 525518 3612 525524 3664
rect 525576 3652 525582 3664
rect 573818 3652 573824 3664
rect 525576 3624 573824 3652
rect 525576 3612 525582 3624
rect 573818 3612 573824 3624
rect 573876 3612 573882 3664
rect 527450 3584 527456 3596
rect 523972 3556 527456 3584
rect 527450 3544 527456 3556
rect 527508 3544 527514 3596
rect 529842 3544 529848 3596
rect 529900 3584 529906 3596
rect 582190 3584 582196 3596
rect 529900 3556 582196 3584
rect 529900 3544 529906 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 425057 3519 425115 3525
rect 425057 3516 425069 3519
rect 422864 3488 425069 3516
rect 421285 3479 421343 3485
rect 425057 3485 425069 3488
rect 425103 3485 425115 3519
rect 425057 3479 425115 3485
rect 426342 3476 426348 3528
rect 426400 3516 426406 3528
rect 428458 3516 428464 3528
rect 426400 3488 428464 3516
rect 426400 3476 426406 3488
rect 428458 3476 428464 3488
rect 428516 3476 428522 3528
rect 432322 3476 432328 3528
rect 432380 3516 432386 3528
rect 451550 3516 451556 3528
rect 432380 3488 451556 3516
rect 432380 3476 432386 3488
rect 451550 3476 451556 3488
rect 451608 3476 451614 3528
rect 459738 3516 459744 3528
rect 451936 3488 459744 3516
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 16022 3408 16028 3460
rect 16080 3448 16086 3460
rect 237558 3448 237564 3460
rect 16080 3420 237564 3448
rect 16080 3408 16086 3420
rect 237558 3408 237564 3420
rect 237616 3408 237622 3460
rect 261018 3408 261024 3460
rect 261076 3448 261082 3460
rect 356054 3448 356060 3460
rect 261076 3420 356060 3448
rect 261076 3408 261082 3420
rect 356054 3408 356060 3420
rect 356112 3408 356118 3460
rect 368014 3408 368020 3460
rect 368072 3448 368078 3460
rect 374641 3451 374699 3457
rect 374641 3448 374653 3451
rect 368072 3420 374653 3448
rect 368072 3408 368078 3420
rect 374641 3417 374653 3420
rect 374687 3417 374699 3451
rect 374641 3411 374699 3417
rect 374733 3451 374791 3457
rect 374733 3417 374745 3451
rect 374779 3448 374791 3451
rect 402425 3451 402483 3457
rect 402425 3448 402437 3451
rect 374779 3420 402437 3448
rect 374779 3417 374791 3420
rect 374733 3411 374791 3417
rect 402425 3417 402437 3420
rect 402471 3417 402483 3451
rect 402425 3411 402483 3417
rect 402514 3408 402520 3460
rect 402572 3448 402578 3460
rect 403529 3451 403587 3457
rect 403529 3448 403541 3451
rect 402572 3420 403541 3448
rect 402572 3408 402578 3420
rect 403529 3417 403541 3420
rect 403575 3417 403587 3451
rect 408405 3451 408463 3457
rect 408405 3448 408417 3451
rect 403529 3411 403587 3417
rect 403636 3420 408417 3448
rect 36170 3340 36176 3392
rect 36228 3380 36234 3392
rect 39298 3380 39304 3392
rect 36228 3352 39304 3380
rect 36228 3340 36234 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 50356 3352 58296 3380
rect 11238 3272 11244 3324
rect 11296 3312 11302 3324
rect 17218 3312 17224 3324
rect 11296 3284 17224 3312
rect 11296 3272 11302 3284
rect 17218 3272 17224 3284
rect 17276 3272 17282 3324
rect 20714 3272 20720 3324
rect 20772 3312 20778 3324
rect 28258 3312 28264 3324
rect 20772 3284 28264 3312
rect 20772 3272 20778 3284
rect 28258 3272 28264 3284
rect 28316 3272 28322 3324
rect 43346 3204 43352 3256
rect 43404 3244 43410 3256
rect 50356 3244 50384 3352
rect 54018 3272 54024 3324
rect 54076 3312 54082 3324
rect 57238 3312 57244 3324
rect 54076 3284 57244 3312
rect 54076 3272 54082 3284
rect 57238 3272 57244 3284
rect 57296 3272 57302 3324
rect 58268 3312 58296 3352
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64782 3380 64788 3392
rect 63644 3352 64788 3380
rect 63644 3340 63650 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 257338 3380 257344 3392
rect 71792 3352 257344 3380
rect 61378 3312 61384 3324
rect 58268 3284 61384 3312
rect 61378 3272 61384 3284
rect 61436 3272 61442 3324
rect 43404 3216 50384 3244
rect 43404 3204 43410 3216
rect 64782 3204 64788 3256
rect 64840 3244 64846 3256
rect 71792 3244 71820 3352
rect 257338 3340 257344 3352
rect 257396 3340 257402 3392
rect 268102 3340 268108 3392
rect 268160 3380 268166 3392
rect 278041 3383 278099 3389
rect 278041 3380 278053 3383
rect 268160 3352 278053 3380
rect 268160 3340 268166 3352
rect 278041 3349 278053 3352
rect 278087 3349 278099 3383
rect 278041 3343 278099 3349
rect 282454 3340 282460 3392
rect 282512 3380 282518 3392
rect 294598 3380 294604 3392
rect 282512 3352 294604 3380
rect 282512 3340 282518 3352
rect 294598 3340 294604 3352
rect 294656 3340 294662 3392
rect 295518 3340 295524 3392
rect 295576 3380 295582 3392
rect 318794 3380 318800 3392
rect 295576 3352 318800 3380
rect 295576 3340 295582 3352
rect 318794 3340 318800 3352
rect 318852 3340 318858 3392
rect 324038 3340 324044 3392
rect 324096 3380 324102 3392
rect 346486 3380 346492 3392
rect 324096 3352 346492 3380
rect 324096 3340 324102 3352
rect 346486 3340 346492 3352
rect 346544 3340 346550 3392
rect 353754 3340 353760 3392
rect 353812 3380 353818 3392
rect 393961 3383 394019 3389
rect 393961 3380 393973 3383
rect 353812 3352 393973 3380
rect 353812 3340 353818 3352
rect 393961 3349 393973 3352
rect 394007 3349 394019 3383
rect 393961 3343 394019 3349
rect 396626 3340 396632 3392
rect 396684 3380 396690 3392
rect 403636 3380 403664 3420
rect 408405 3417 408417 3420
rect 408451 3417 408463 3451
rect 408405 3411 408463 3417
rect 408494 3408 408500 3460
rect 408552 3448 408558 3460
rect 409782 3448 409788 3460
rect 408552 3420 409788 3448
rect 408552 3408 408558 3420
rect 409782 3408 409788 3420
rect 409840 3408 409846 3460
rect 409877 3451 409935 3457
rect 409877 3417 409889 3451
rect 409923 3448 409935 3451
rect 412545 3451 412603 3457
rect 412545 3448 412557 3451
rect 409923 3420 412557 3448
rect 409923 3417 409935 3420
rect 409877 3411 409935 3417
rect 412545 3417 412557 3420
rect 412591 3417 412603 3451
rect 412545 3411 412603 3417
rect 412634 3408 412640 3460
rect 412692 3448 412698 3460
rect 413462 3448 413468 3460
rect 412692 3420 413468 3448
rect 412692 3408 412698 3420
rect 413462 3408 413468 3420
rect 413520 3408 413526 3460
rect 413649 3451 413707 3457
rect 413649 3417 413661 3451
rect 413695 3448 413707 3451
rect 418065 3451 418123 3457
rect 418065 3448 418077 3451
rect 413695 3420 418077 3448
rect 413695 3417 413707 3420
rect 413649 3411 413707 3417
rect 418065 3417 418077 3420
rect 418111 3417 418123 3451
rect 418065 3411 418123 3417
rect 427725 3451 427783 3457
rect 427725 3417 427737 3451
rect 427771 3448 427783 3451
rect 427771 3420 443132 3448
rect 427771 3417 427783 3420
rect 427725 3411 427783 3417
rect 409509 3383 409567 3389
rect 409509 3380 409521 3383
rect 396684 3352 403664 3380
rect 403728 3352 409521 3380
rect 396684 3340 396690 3352
rect 71866 3272 71872 3324
rect 71924 3312 71930 3324
rect 258718 3312 258724 3324
rect 71924 3284 258724 3312
rect 71924 3272 71930 3284
rect 258718 3272 258724 3284
rect 258776 3272 258782 3324
rect 276474 3272 276480 3324
rect 276532 3312 276538 3324
rect 280157 3315 280215 3321
rect 280157 3312 280169 3315
rect 276532 3284 280169 3312
rect 276532 3272 276538 3284
rect 280157 3281 280169 3284
rect 280203 3281 280215 3315
rect 280157 3275 280215 3281
rect 292577 3315 292635 3321
rect 292577 3281 292589 3315
rect 292623 3312 292635 3315
rect 302145 3315 302203 3321
rect 302145 3312 302157 3315
rect 292623 3284 302157 3312
rect 292623 3281 292635 3284
rect 292577 3275 292635 3281
rect 302145 3281 302157 3284
rect 302191 3281 302203 3315
rect 302145 3275 302203 3281
rect 306190 3272 306196 3324
rect 306248 3312 306254 3324
rect 325602 3312 325608 3324
rect 306248 3284 325608 3312
rect 306248 3272 306254 3284
rect 325602 3272 325608 3284
rect 325660 3272 325666 3324
rect 335173 3315 335231 3321
rect 335173 3281 335185 3315
rect 335219 3312 335231 3315
rect 347958 3312 347964 3324
rect 335219 3284 347964 3312
rect 335219 3281 335231 3284
rect 335173 3275 335231 3281
rect 347958 3272 347964 3284
rect 348016 3272 348022 3324
rect 363233 3315 363291 3321
rect 363233 3281 363245 3315
rect 363279 3312 363291 3315
rect 366450 3312 366456 3324
rect 363279 3284 366456 3312
rect 363279 3281 363291 3284
rect 363233 3275 363291 3281
rect 366450 3272 366456 3284
rect 366508 3272 366514 3324
rect 403437 3315 403495 3321
rect 403437 3312 403449 3315
rect 370332 3284 403449 3312
rect 64840 3216 71820 3244
rect 64840 3204 64846 3216
rect 77846 3204 77852 3256
rect 77904 3244 77910 3256
rect 78582 3244 78588 3256
rect 77904 3216 78588 3244
rect 77904 3204 77910 3216
rect 78582 3204 78588 3216
rect 78640 3204 78646 3256
rect 81434 3204 81440 3256
rect 81492 3244 81498 3256
rect 82722 3244 82728 3256
rect 81492 3216 82728 3244
rect 81492 3204 81498 3216
rect 82722 3204 82728 3216
rect 82780 3204 82786 3256
rect 84838 3244 84844 3256
rect 82832 3216 84844 3244
rect 27890 3136 27896 3188
rect 27948 3176 27954 3188
rect 28902 3176 28908 3188
rect 27948 3148 28908 3176
rect 27948 3136 27954 3148
rect 28902 3136 28908 3148
rect 28960 3136 28966 3188
rect 29086 3136 29092 3188
rect 29144 3176 29150 3188
rect 32398 3176 32404 3188
rect 29144 3148 32404 3176
rect 29144 3136 29150 3148
rect 32398 3136 32404 3148
rect 32456 3136 32462 3188
rect 61194 3136 61200 3188
rect 61252 3176 61258 3188
rect 66898 3176 66904 3188
rect 61252 3148 66904 3176
rect 61252 3136 61258 3148
rect 66898 3136 66904 3148
rect 66956 3136 66962 3188
rect 82630 3136 82636 3188
rect 82688 3176 82694 3188
rect 82832 3176 82860 3216
rect 84838 3204 84844 3216
rect 84896 3204 84902 3256
rect 84930 3204 84936 3256
rect 84988 3244 84994 3256
rect 85482 3244 85488 3256
rect 84988 3216 85488 3244
rect 84988 3204 84994 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 88518 3204 88524 3256
rect 88576 3244 88582 3256
rect 89622 3244 89628 3256
rect 88576 3216 89628 3244
rect 88576 3204 88582 3216
rect 89622 3204 89628 3216
rect 89680 3204 89686 3256
rect 261478 3244 261484 3256
rect 89732 3216 261484 3244
rect 82688 3148 82860 3176
rect 82909 3179 82967 3185
rect 82688 3136 82694 3148
rect 82909 3145 82921 3179
rect 82955 3176 82967 3179
rect 89732 3176 89760 3216
rect 261478 3204 261484 3216
rect 261536 3204 261542 3256
rect 288342 3204 288348 3256
rect 288400 3244 288406 3256
rect 292942 3244 292948 3256
rect 288400 3216 292948 3244
rect 288400 3204 288406 3216
rect 292942 3204 292948 3216
rect 293000 3204 293006 3256
rect 302602 3204 302608 3256
rect 302660 3244 302666 3256
rect 320174 3244 320180 3256
rect 302660 3216 320180 3244
rect 302660 3204 302666 3216
rect 320174 3204 320180 3216
rect 320232 3204 320238 3256
rect 328822 3204 328828 3256
rect 328880 3244 328886 3256
rect 363690 3244 363696 3256
rect 328880 3216 363696 3244
rect 328880 3204 328886 3216
rect 363690 3204 363696 3216
rect 363748 3204 363754 3256
rect 82955 3148 89760 3176
rect 82955 3145 82967 3148
rect 82909 3139 82967 3145
rect 89806 3136 89812 3188
rect 89864 3176 89870 3188
rect 262858 3176 262864 3188
rect 89864 3148 262864 3176
rect 89864 3136 89870 3148
rect 262858 3136 262864 3148
rect 262916 3136 262922 3188
rect 285950 3136 285956 3188
rect 286008 3176 286014 3188
rect 286962 3176 286968 3188
rect 286008 3148 286968 3176
rect 286008 3136 286014 3148
rect 286962 3136 286968 3148
rect 287020 3136 287026 3188
rect 293126 3136 293132 3188
rect 293184 3176 293190 3188
rect 293862 3176 293868 3188
rect 293184 3148 293868 3176
rect 293184 3136 293190 3148
rect 293862 3136 293868 3148
rect 293920 3136 293926 3188
rect 309778 3136 309784 3188
rect 309836 3176 309842 3188
rect 323578 3176 323584 3188
rect 309836 3148 323584 3176
rect 309836 3136 309842 3148
rect 323578 3136 323584 3148
rect 323636 3136 323642 3188
rect 327626 3136 327632 3188
rect 327684 3176 327690 3188
rect 335173 3179 335231 3185
rect 335173 3176 335185 3179
rect 327684 3148 335185 3176
rect 327684 3136 327690 3148
rect 335173 3145 335185 3148
rect 335219 3145 335231 3179
rect 335173 3139 335231 3145
rect 343082 3136 343088 3188
rect 343140 3176 343146 3188
rect 369857 3179 369915 3185
rect 369857 3176 369869 3179
rect 343140 3148 369869 3176
rect 343140 3136 343146 3148
rect 369857 3145 369869 3148
rect 369903 3145 369915 3179
rect 369857 3139 369915 3145
rect 95694 3068 95700 3120
rect 95752 3108 95758 3120
rect 96522 3108 96528 3120
rect 95752 3080 96528 3108
rect 95752 3068 95758 3080
rect 96522 3068 96528 3080
rect 96580 3068 96586 3120
rect 97258 3108 97264 3120
rect 96632 3080 97264 3108
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 15838 3040 15844 3052
rect 10100 3012 15844 3040
rect 10100 3000 10106 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 68278 3000 68284 3052
rect 68336 3040 68342 3052
rect 71038 3040 71044 3052
rect 68336 3012 71044 3040
rect 68336 3000 68342 3012
rect 71038 3000 71044 3012
rect 71096 3000 71102 3052
rect 93302 3000 93308 3052
rect 93360 3040 93366 3052
rect 96632 3040 96660 3080
rect 97258 3068 97264 3080
rect 97316 3068 97322 3120
rect 98086 3068 98092 3120
rect 98144 3108 98150 3120
rect 99190 3108 99196 3120
rect 98144 3080 99196 3108
rect 98144 3068 98150 3080
rect 99190 3068 99196 3080
rect 99248 3068 99254 3120
rect 102778 3068 102784 3120
rect 102836 3108 102842 3120
rect 103422 3108 103428 3120
rect 102836 3080 103428 3108
rect 102836 3068 102842 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 103974 3068 103980 3120
rect 104032 3108 104038 3120
rect 104802 3108 104808 3120
rect 104032 3080 104808 3108
rect 104032 3068 104038 3080
rect 104802 3068 104808 3080
rect 104860 3068 104866 3120
rect 106366 3068 106372 3120
rect 106424 3108 106430 3120
rect 107562 3108 107568 3120
rect 106424 3080 107568 3108
rect 106424 3068 106430 3080
rect 107562 3068 107568 3080
rect 107620 3068 107626 3120
rect 111150 3068 111156 3120
rect 111208 3108 111214 3120
rect 111702 3108 111708 3120
rect 111208 3080 111708 3108
rect 111208 3068 111214 3080
rect 111702 3068 111708 3080
rect 111760 3068 111766 3120
rect 264238 3108 264244 3120
rect 111812 3080 264244 3108
rect 93360 3012 96660 3040
rect 93360 3000 93366 3012
rect 96890 3000 96896 3052
rect 96948 3040 96954 3052
rect 111812 3040 111840 3080
rect 264238 3068 264244 3080
rect 264296 3068 264302 3120
rect 313366 3068 313372 3120
rect 313424 3108 313430 3120
rect 325510 3108 325516 3120
rect 313424 3080 325516 3108
rect 313424 3068 313430 3080
rect 325510 3068 325516 3080
rect 325568 3068 325574 3120
rect 335906 3068 335912 3120
rect 335964 3108 335970 3120
rect 363233 3111 363291 3117
rect 363233 3108 363245 3111
rect 335964 3080 363245 3108
rect 335964 3068 335970 3080
rect 363233 3077 363245 3080
rect 363279 3077 363291 3111
rect 363233 3071 363291 3077
rect 363322 3068 363328 3120
rect 363380 3108 363386 3120
rect 370332 3108 370360 3284
rect 403437 3281 403449 3284
rect 403483 3281 403495 3315
rect 403728 3312 403756 3352
rect 409509 3349 409521 3352
rect 409555 3349 409567 3383
rect 413373 3383 413431 3389
rect 413373 3380 413385 3383
rect 409509 3343 409567 3349
rect 409616 3352 413385 3380
rect 403437 3275 403495 3281
rect 403544 3284 403756 3312
rect 403805 3315 403863 3321
rect 370406 3204 370412 3256
rect 370464 3244 370470 3256
rect 393869 3247 393927 3253
rect 393869 3244 393881 3247
rect 370464 3216 393881 3244
rect 370464 3204 370470 3216
rect 393869 3213 393881 3216
rect 393915 3213 393927 3247
rect 393869 3207 393927 3213
rect 402425 3247 402483 3253
rect 402425 3213 402437 3247
rect 402471 3244 402483 3247
rect 403345 3247 403403 3253
rect 403345 3244 403357 3247
rect 402471 3216 403357 3244
rect 402471 3213 402483 3216
rect 402425 3207 402483 3213
rect 403345 3213 403357 3216
rect 403391 3213 403403 3247
rect 403544 3244 403572 3284
rect 403805 3281 403817 3315
rect 403851 3312 403863 3315
rect 407114 3312 407120 3324
rect 403851 3284 407120 3312
rect 403851 3281 403863 3284
rect 403805 3275 403863 3281
rect 407114 3272 407120 3284
rect 407172 3272 407178 3324
rect 407298 3272 407304 3324
rect 407356 3312 407362 3324
rect 409616 3312 409644 3352
rect 413373 3349 413385 3352
rect 413419 3349 413431 3383
rect 413373 3343 413431 3349
rect 413557 3383 413615 3389
rect 413557 3349 413569 3383
rect 413603 3380 413615 3383
rect 417418 3380 417424 3392
rect 413603 3352 417424 3380
rect 413603 3349 413615 3352
rect 413557 3343 413615 3349
rect 417418 3340 417424 3352
rect 417476 3340 417482 3392
rect 417970 3340 417976 3392
rect 418028 3380 418034 3392
rect 418157 3383 418215 3389
rect 418157 3380 418169 3383
rect 418028 3352 418169 3380
rect 418028 3340 418034 3352
rect 418157 3349 418169 3352
rect 418203 3349 418215 3383
rect 418157 3343 418215 3349
rect 418249 3383 418307 3389
rect 418249 3349 418261 3383
rect 418295 3380 418307 3383
rect 435358 3380 435364 3392
rect 418295 3352 435364 3380
rect 418295 3349 418307 3352
rect 418249 3343 418307 3349
rect 435358 3340 435364 3352
rect 435416 3340 435422 3392
rect 443104 3380 443132 3420
rect 444190 3408 444196 3460
rect 444248 3448 444254 3460
rect 446398 3448 446404 3460
rect 444248 3420 446404 3448
rect 444248 3408 444254 3420
rect 446398 3408 446404 3420
rect 446456 3408 446462 3460
rect 446582 3408 446588 3460
rect 446640 3448 446646 3460
rect 451936 3448 451964 3488
rect 459738 3476 459744 3488
rect 459796 3476 459802 3528
rect 487062 3476 487068 3528
rect 487120 3516 487126 3528
rect 498930 3516 498936 3528
rect 487120 3488 498936 3516
rect 487120 3476 487126 3488
rect 498930 3476 498936 3488
rect 498988 3476 498994 3528
rect 500862 3476 500868 3528
rect 500920 3516 500926 3528
rect 526254 3516 526260 3528
rect 500920 3488 526260 3516
rect 500920 3476 500926 3488
rect 526254 3476 526260 3488
rect 526312 3476 526318 3528
rect 528462 3476 528468 3528
rect 528520 3516 528526 3528
rect 578602 3516 578608 3528
rect 528520 3488 578608 3516
rect 528520 3476 528526 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 446640 3420 451964 3448
rect 446640 3408 446646 3420
rect 452470 3408 452476 3460
rect 452528 3448 452534 3460
rect 457438 3448 457444 3460
rect 452528 3420 457444 3448
rect 452528 3408 452534 3420
rect 457438 3408 457444 3420
rect 457496 3408 457502 3460
rect 462038 3408 462044 3460
rect 462096 3448 462102 3460
rect 466454 3448 466460 3460
rect 462096 3420 466460 3448
rect 462096 3408 462102 3420
rect 466454 3408 466460 3420
rect 466512 3408 466518 3460
rect 488442 3408 488448 3460
rect 488500 3448 488506 3460
rect 501230 3448 501236 3460
rect 488500 3420 501236 3448
rect 488500 3408 488506 3420
rect 501230 3408 501236 3420
rect 501288 3408 501294 3460
rect 502242 3408 502248 3460
rect 502300 3448 502306 3460
rect 528646 3448 528652 3460
rect 502300 3420 528652 3448
rect 502300 3408 502306 3420
rect 528646 3408 528652 3420
rect 528704 3408 528710 3460
rect 529750 3408 529756 3460
rect 529808 3448 529814 3460
rect 580994 3448 581000 3460
rect 529808 3420 581000 3448
rect 529808 3408 529814 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 444558 3380 444564 3392
rect 443104 3352 444564 3380
rect 444558 3340 444564 3352
rect 444616 3340 444622 3392
rect 459646 3340 459652 3392
rect 459704 3380 459710 3392
rect 464338 3380 464344 3392
rect 459704 3352 464344 3380
rect 459704 3340 459710 3352
rect 464338 3340 464344 3352
rect 464396 3340 464402 3392
rect 482830 3340 482836 3392
rect 482888 3380 482894 3392
rect 489362 3380 489368 3392
rect 482888 3352 489368 3380
rect 482888 3340 482894 3352
rect 489362 3340 489368 3352
rect 489420 3340 489426 3392
rect 492582 3340 492588 3392
rect 492640 3380 492646 3392
rect 508406 3380 508412 3392
rect 492640 3352 508412 3380
rect 492640 3340 492646 3352
rect 508406 3340 508412 3352
rect 508464 3340 508470 3392
rect 509697 3383 509755 3389
rect 509697 3349 509709 3383
rect 509743 3380 509755 3383
rect 516778 3380 516784 3392
rect 509743 3352 516784 3380
rect 509743 3349 509755 3352
rect 509697 3343 509755 3349
rect 516778 3340 516784 3352
rect 516836 3340 516842 3392
rect 517422 3340 517428 3392
rect 517480 3380 517486 3392
rect 557166 3380 557172 3392
rect 517480 3352 557172 3380
rect 517480 3340 517486 3352
rect 557166 3340 557172 3352
rect 557224 3340 557230 3392
rect 558178 3340 558184 3392
rect 558236 3380 558242 3392
rect 558236 3352 569172 3380
rect 558236 3340 558242 3352
rect 407356 3284 409644 3312
rect 407356 3272 407362 3284
rect 409690 3272 409696 3324
rect 409748 3312 409754 3324
rect 431218 3312 431224 3324
rect 409748 3284 431224 3312
rect 409748 3272 409754 3284
rect 431218 3272 431224 3284
rect 431276 3272 431282 3324
rect 441798 3272 441804 3324
rect 441856 3312 441862 3324
rect 449158 3312 449164 3324
rect 441856 3284 449164 3312
rect 441856 3272 441862 3284
rect 449158 3272 449164 3284
rect 449216 3272 449222 3324
rect 464430 3272 464436 3324
rect 464488 3312 464494 3324
rect 464982 3312 464988 3324
rect 464488 3284 464988 3312
rect 464488 3272 464494 3284
rect 464982 3272 464988 3284
rect 465040 3272 465046 3324
rect 481542 3272 481548 3324
rect 481600 3312 481606 3324
rect 486970 3312 486976 3324
rect 481600 3284 486976 3312
rect 481600 3272 481606 3284
rect 486970 3272 486976 3284
rect 487028 3272 487034 3324
rect 488350 3272 488356 3324
rect 488408 3312 488414 3324
rect 502426 3312 502432 3324
rect 488408 3284 502432 3312
rect 488408 3272 488414 3284
rect 502426 3272 502432 3284
rect 502484 3272 502490 3324
rect 514662 3272 514668 3324
rect 514720 3312 514726 3324
rect 552382 3312 552388 3324
rect 514720 3284 552388 3312
rect 514720 3272 514726 3284
rect 552382 3272 552388 3284
rect 552440 3272 552446 3324
rect 556798 3272 556804 3324
rect 556856 3312 556862 3324
rect 565538 3312 565544 3324
rect 556856 3284 565544 3312
rect 556856 3272 556862 3284
rect 565538 3272 565544 3284
rect 565596 3272 565602 3324
rect 403345 3207 403403 3213
rect 403452 3216 403572 3244
rect 403621 3247 403679 3253
rect 381170 3136 381176 3188
rect 381228 3176 381234 3188
rect 403253 3179 403311 3185
rect 403253 3176 403265 3179
rect 381228 3148 403265 3176
rect 381228 3136 381234 3148
rect 403253 3145 403265 3148
rect 403299 3145 403311 3179
rect 403253 3139 403311 3145
rect 374638 3108 374644 3120
rect 363380 3080 370360 3108
rect 372264 3080 374644 3108
rect 363380 3068 363386 3080
rect 264330 3040 264336 3052
rect 96948 3012 98776 3040
rect 96948 3000 96954 3012
rect 79042 2932 79048 2984
rect 79100 2972 79106 2984
rect 82909 2975 82967 2981
rect 82909 2972 82921 2975
rect 79100 2944 82921 2972
rect 79100 2932 79106 2944
rect 82909 2941 82921 2944
rect 82955 2941 82967 2975
rect 82909 2935 82967 2941
rect 86126 2932 86132 2984
rect 86184 2972 86190 2984
rect 98641 2975 98699 2981
rect 98641 2972 98653 2975
rect 86184 2944 98653 2972
rect 86184 2932 86190 2944
rect 98641 2941 98653 2944
rect 98687 2941 98699 2975
rect 98748 2972 98776 3012
rect 99392 3012 111840 3040
rect 111904 3012 264336 3040
rect 99392 2972 99420 3012
rect 106918 2972 106924 2984
rect 98748 2944 99420 2972
rect 100404 2944 106924 2972
rect 98641 2935 98699 2941
rect 75454 2864 75460 2916
rect 75512 2904 75518 2916
rect 100404 2904 100432 2944
rect 106918 2932 106924 2944
rect 106976 2932 106982 2984
rect 75512 2876 100432 2904
rect 75512 2864 75518 2876
rect 100478 2864 100484 2916
rect 100536 2904 100542 2916
rect 111904 2904 111932 3012
rect 264330 3000 264336 3012
rect 264388 3000 264394 3052
rect 320450 3000 320456 3052
rect 320508 3040 320514 3052
rect 328546 3040 328552 3052
rect 320508 3012 328552 3040
rect 320508 3000 320514 3012
rect 328546 3000 328552 3012
rect 328604 3000 328610 3052
rect 338298 3000 338304 3052
rect 338356 3040 338362 3052
rect 339402 3040 339408 3052
rect 338356 3012 339408 3040
rect 338356 3000 338362 3012
rect 339402 3000 339408 3012
rect 339460 3000 339466 3052
rect 350258 3000 350264 3052
rect 350316 3040 350322 3052
rect 372264 3040 372292 3080
rect 374638 3068 374644 3080
rect 374696 3068 374702 3120
rect 375190 3068 375196 3120
rect 375248 3108 375254 3120
rect 403452 3108 403480 3216
rect 403621 3213 403633 3247
rect 403667 3244 403679 3247
rect 413370 3244 413376 3256
rect 403667 3216 413376 3244
rect 403667 3213 403679 3216
rect 403621 3207 403679 3213
rect 413370 3204 413376 3216
rect 413428 3204 413434 3256
rect 414385 3247 414443 3253
rect 414385 3213 414397 3247
rect 414431 3244 414443 3247
rect 416777 3247 416835 3253
rect 416777 3244 416789 3247
rect 414431 3216 416789 3244
rect 414431 3213 414443 3216
rect 414385 3207 414443 3213
rect 416777 3213 416789 3216
rect 416823 3213 416835 3247
rect 416777 3207 416835 3213
rect 416866 3204 416872 3256
rect 416924 3244 416930 3256
rect 438118 3244 438124 3256
rect 416924 3216 438124 3244
rect 416924 3204 416930 3216
rect 438118 3204 438124 3216
rect 438176 3204 438182 3256
rect 485038 3204 485044 3256
rect 485096 3244 485102 3256
rect 488166 3244 488172 3256
rect 485096 3216 488172 3244
rect 485096 3204 485102 3216
rect 488166 3204 488172 3216
rect 488224 3204 488230 3256
rect 489822 3204 489828 3256
rect 489880 3244 489886 3256
rect 504818 3244 504824 3256
rect 489880 3216 504824 3244
rect 489880 3204 489886 3216
rect 504818 3204 504824 3216
rect 504876 3204 504882 3256
rect 511810 3204 511816 3256
rect 511868 3244 511874 3256
rect 540149 3247 540207 3253
rect 540149 3244 540161 3247
rect 511868 3216 540161 3244
rect 511868 3204 511874 3216
rect 540149 3213 540161 3216
rect 540195 3213 540207 3247
rect 540149 3207 540207 3213
rect 540238 3204 540244 3256
rect 540296 3244 540302 3256
rect 541710 3244 541716 3256
rect 540296 3216 541716 3244
rect 540296 3204 540302 3216
rect 541710 3204 541716 3216
rect 541768 3204 541774 3256
rect 547138 3204 547144 3256
rect 547196 3244 547202 3256
rect 550082 3244 550088 3256
rect 547196 3216 550088 3244
rect 547196 3204 547202 3216
rect 550082 3204 550088 3216
rect 550140 3204 550146 3256
rect 558362 3244 558368 3256
rect 554884 3216 558368 3244
rect 403529 3179 403587 3185
rect 403529 3145 403541 3179
rect 403575 3176 403587 3179
rect 422849 3179 422907 3185
rect 403575 3148 418568 3176
rect 403575 3145 403587 3148
rect 403529 3139 403587 3145
rect 375248 3080 403480 3108
rect 375248 3068 375254 3080
rect 403618 3068 403624 3120
rect 403676 3108 403682 3120
rect 409509 3111 409567 3117
rect 403676 3080 409460 3108
rect 403676 3068 403682 3080
rect 350316 3012 372292 3040
rect 350316 3000 350322 3012
rect 373994 3000 374000 3052
rect 374052 3040 374058 3052
rect 375282 3040 375288 3052
rect 374052 3012 375288 3040
rect 374052 3000 374058 3012
rect 375282 3000 375288 3012
rect 375340 3000 375346 3052
rect 378870 3000 378876 3052
rect 378928 3040 378934 3052
rect 409432 3040 409460 3080
rect 409509 3077 409521 3111
rect 409555 3108 409567 3111
rect 414658 3108 414664 3120
rect 409555 3080 414664 3108
rect 409555 3077 409567 3080
rect 409509 3071 409567 3077
rect 414658 3068 414664 3080
rect 414716 3068 414722 3120
rect 415670 3068 415676 3120
rect 415728 3108 415734 3120
rect 416682 3108 416688 3120
rect 415728 3080 416688 3108
rect 415728 3068 415734 3080
rect 416682 3068 416688 3080
rect 416740 3068 416746 3120
rect 416777 3111 416835 3117
rect 416777 3077 416789 3111
rect 416823 3108 416835 3111
rect 418249 3111 418307 3117
rect 418249 3108 418261 3111
rect 416823 3080 418261 3108
rect 416823 3077 416835 3080
rect 416777 3071 416835 3077
rect 418249 3077 418261 3080
rect 418295 3077 418307 3111
rect 418540 3108 418568 3148
rect 422849 3145 422861 3179
rect 422895 3176 422907 3179
rect 430574 3176 430580 3188
rect 422895 3148 430580 3176
rect 422895 3145 422907 3148
rect 422849 3139 422907 3145
rect 430574 3136 430580 3148
rect 430632 3136 430638 3188
rect 493318 3136 493324 3188
rect 493376 3176 493382 3188
rect 496538 3176 496544 3188
rect 493376 3148 496544 3176
rect 493376 3136 493382 3148
rect 496538 3136 496544 3148
rect 496596 3136 496602 3188
rect 510522 3136 510528 3188
rect 510580 3176 510586 3188
rect 510580 3148 540284 3176
rect 510580 3136 510586 3148
rect 424318 3108 424324 3120
rect 418540 3080 424324 3108
rect 418249 3071 418307 3077
rect 424318 3068 424324 3080
rect 424376 3068 424382 3120
rect 470318 3068 470324 3120
rect 470376 3108 470382 3120
rect 470686 3108 470692 3120
rect 470376 3080 470692 3108
rect 470376 3068 470382 3080
rect 470686 3068 470692 3080
rect 470744 3068 470750 3120
rect 501598 3068 501604 3120
rect 501656 3108 501662 3120
rect 506014 3108 506020 3120
rect 501656 3080 506020 3108
rect 501656 3068 501662 3080
rect 506014 3068 506020 3080
rect 506072 3068 506078 3120
rect 511902 3068 511908 3120
rect 511960 3108 511966 3120
rect 540256 3108 540284 3148
rect 540330 3136 540336 3188
rect 540388 3176 540394 3188
rect 544102 3176 544108 3188
rect 540388 3148 544108 3176
rect 540388 3136 540394 3148
rect 544102 3136 544108 3148
rect 544160 3136 544166 3188
rect 545298 3108 545304 3120
rect 511960 3080 539088 3108
rect 540256 3080 545304 3108
rect 511960 3068 511966 3080
rect 412634 3040 412640 3052
rect 378928 3012 409368 3040
rect 409432 3012 412640 3040
rect 378928 3000 378934 3012
rect 112346 2932 112352 2984
rect 112404 2972 112410 2984
rect 113082 2972 113088 2984
rect 112404 2944 113088 2972
rect 112404 2932 112410 2944
rect 113082 2932 113088 2944
rect 113140 2932 113146 2984
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 115934 2932 115940 2984
rect 115992 2972 115998 2984
rect 116946 2972 116952 2984
rect 115992 2944 116952 2972
rect 115992 2932 115998 2944
rect 116946 2932 116952 2944
rect 117004 2932 117010 2984
rect 119430 2932 119436 2984
rect 119488 2972 119494 2984
rect 119982 2972 119988 2984
rect 119488 2944 119988 2972
rect 119488 2932 119494 2944
rect 119982 2932 119988 2944
rect 120040 2932 120046 2984
rect 120626 2932 120632 2984
rect 120684 2972 120690 2984
rect 121362 2972 121368 2984
rect 120684 2944 121368 2972
rect 120684 2932 120690 2944
rect 121362 2932 121368 2944
rect 121420 2932 121426 2984
rect 266906 2972 266912 2984
rect 121564 2944 266912 2972
rect 100536 2876 111932 2904
rect 100536 2864 100542 2876
rect 114738 2864 114744 2916
rect 114796 2904 114802 2916
rect 121457 2907 121515 2913
rect 121457 2904 121469 2907
rect 114796 2876 121469 2904
rect 114796 2864 114802 2876
rect 121457 2873 121469 2876
rect 121503 2873 121515 2907
rect 121457 2867 121515 2873
rect 98641 2839 98699 2845
rect 98641 2805 98653 2839
rect 98687 2836 98699 2839
rect 105538 2836 105544 2848
rect 98687 2808 105544 2836
rect 98687 2805 98699 2808
rect 98641 2799 98699 2805
rect 105538 2796 105544 2808
rect 105596 2796 105602 2848
rect 107562 2796 107568 2848
rect 107620 2836 107626 2848
rect 121564 2836 121592 2944
rect 266906 2932 266912 2944
rect 266964 2932 266970 2984
rect 341886 2932 341892 2984
rect 341944 2972 341950 2984
rect 351822 2972 351828 2984
rect 341944 2944 351828 2972
rect 341944 2932 341950 2944
rect 351822 2932 351828 2944
rect 351880 2932 351886 2984
rect 360930 2932 360936 2984
rect 360988 2972 360994 2984
rect 374733 2975 374791 2981
rect 374733 2972 374745 2975
rect 360988 2944 374745 2972
rect 360988 2932 360994 2944
rect 374733 2941 374745 2944
rect 374779 2941 374791 2975
rect 374733 2935 374791 2941
rect 377582 2932 377588 2984
rect 377640 2972 377646 2984
rect 403621 2975 403679 2981
rect 403621 2972 403633 2975
rect 377640 2944 403633 2972
rect 377640 2932 377646 2944
rect 403621 2941 403633 2944
rect 403667 2941 403679 2975
rect 403621 2935 403679 2941
rect 406102 2932 406108 2984
rect 406160 2972 406166 2984
rect 409138 2972 409144 2984
rect 406160 2944 409144 2972
rect 406160 2932 406166 2944
rect 409138 2932 409144 2944
rect 409196 2932 409202 2984
rect 121641 2907 121699 2913
rect 121641 2873 121653 2907
rect 121687 2904 121699 2907
rect 268378 2904 268384 2916
rect 121687 2876 268384 2904
rect 121687 2873 121699 2876
rect 121641 2867 121699 2873
rect 268378 2864 268384 2876
rect 268436 2864 268442 2916
rect 369857 2907 369915 2913
rect 369857 2873 369869 2907
rect 369903 2904 369915 2907
rect 376018 2904 376024 2916
rect 369903 2876 376024 2904
rect 369903 2873 369915 2876
rect 369857 2867 369915 2873
rect 376018 2864 376024 2876
rect 376076 2864 376082 2916
rect 384666 2864 384672 2916
rect 384724 2904 384730 2916
rect 409233 2907 409291 2913
rect 409233 2904 409245 2907
rect 384724 2876 409245 2904
rect 384724 2864 384730 2876
rect 409233 2873 409245 2876
rect 409279 2873 409291 2907
rect 409340 2904 409368 3012
rect 412634 3000 412640 3012
rect 412692 3000 412698 3052
rect 427078 3040 427084 3052
rect 418816 3012 427084 3040
rect 409414 2932 409420 2984
rect 409472 2972 409478 2984
rect 418816 2972 418844 3012
rect 427078 3000 427084 3012
rect 427136 3000 427142 3052
rect 445386 3000 445392 3052
rect 445444 3040 445450 3052
rect 451918 3040 451924 3052
rect 445444 3012 451924 3040
rect 445444 3000 445450 3012
rect 451918 3000 451924 3012
rect 451976 3000 451982 3052
rect 477402 3000 477408 3052
rect 477460 3040 477466 3052
rect 479886 3040 479892 3052
rect 477460 3012 479892 3040
rect 477460 3000 477466 3012
rect 479886 3000 479892 3012
rect 479944 3000 479950 3052
rect 507762 3000 507768 3052
rect 507820 3040 507826 3052
rect 538122 3040 538128 3052
rect 507820 3012 538128 3040
rect 507820 3000 507826 3012
rect 538122 3000 538128 3012
rect 538180 3000 538186 3052
rect 539060 3040 539088 3080
rect 545298 3068 545304 3080
rect 545356 3068 545362 3120
rect 545758 3068 545764 3120
rect 545816 3108 545822 3120
rect 554774 3108 554780 3120
rect 545816 3080 554780 3108
rect 545816 3068 545822 3080
rect 554774 3068 554780 3080
rect 554832 3068 554838 3120
rect 546494 3040 546500 3052
rect 539060 3012 546500 3040
rect 546494 3000 546500 3012
rect 546552 3000 546558 3052
rect 547230 3000 547236 3052
rect 547288 3040 547294 3052
rect 548886 3040 548892 3052
rect 547288 3012 548892 3040
rect 547288 3000 547294 3012
rect 548886 3000 548892 3012
rect 548944 3000 548950 3052
rect 549898 3000 549904 3052
rect 549956 3040 549962 3052
rect 554884 3040 554912 3216
rect 558362 3204 558368 3216
rect 558420 3204 558426 3256
rect 569144 3244 569172 3352
rect 569218 3340 569224 3392
rect 569276 3380 569282 3392
rect 570230 3380 570236 3392
rect 569276 3352 570236 3380
rect 569276 3340 569282 3352
rect 570230 3340 570236 3352
rect 570288 3340 570294 3392
rect 576210 3244 576216 3256
rect 569144 3216 576216 3244
rect 576210 3204 576216 3216
rect 576268 3204 576274 3256
rect 549956 3012 554912 3040
rect 549956 3000 549962 3012
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 577406 3040 577412 3052
rect 572036 3012 577412 3040
rect 572036 3000 572042 3012
rect 577406 3000 577412 3012
rect 577464 3000 577470 3052
rect 409472 2944 418844 2972
rect 418893 2975 418951 2981
rect 409472 2932 409478 2944
rect 418893 2941 418905 2975
rect 418939 2972 418951 2975
rect 426618 2972 426624 2984
rect 418939 2944 426624 2972
rect 418939 2941 418951 2944
rect 418893 2935 418951 2941
rect 426618 2932 426624 2944
rect 426676 2932 426682 2984
rect 506382 2932 506388 2984
rect 506440 2972 506446 2984
rect 535730 2972 535736 2984
rect 506440 2944 535736 2972
rect 506440 2932 506446 2944
rect 535730 2932 535736 2944
rect 535788 2932 535794 2984
rect 540149 2975 540207 2981
rect 540149 2941 540161 2975
rect 540195 2972 540207 2975
rect 547690 2972 547696 2984
rect 540195 2944 547696 2972
rect 540195 2941 540207 2944
rect 540149 2935 540207 2941
rect 547690 2932 547696 2944
rect 547748 2932 547754 2984
rect 551186 2972 551192 2984
rect 547800 2944 551192 2972
rect 416038 2904 416044 2916
rect 409340 2876 416044 2904
rect 409233 2867 409291 2873
rect 416038 2864 416044 2876
rect 416096 2864 416102 2916
rect 421558 2864 421564 2916
rect 421616 2904 421622 2916
rect 422202 2904 422208 2916
rect 421616 2876 422208 2904
rect 421616 2864 421622 2876
rect 422202 2864 422208 2876
rect 422260 2864 422266 2916
rect 465626 2864 465632 2916
rect 465684 2904 465690 2916
rect 466362 2904 466368 2916
rect 465684 2876 466368 2904
rect 465684 2864 465690 2876
rect 466362 2864 466368 2876
rect 466420 2864 466426 2916
rect 505002 2864 505008 2916
rect 505060 2904 505066 2916
rect 533430 2904 533436 2916
rect 505060 2876 533436 2904
rect 505060 2864 505066 2876
rect 533430 2864 533436 2876
rect 533488 2864 533494 2916
rect 107620 2808 121592 2836
rect 107620 2796 107626 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 269758 2836 269764 2848
rect 121880 2808 269764 2836
rect 121880 2796 121886 2808
rect 269758 2796 269764 2808
rect 269816 2796 269822 2848
rect 310974 2796 310980 2848
rect 311032 2836 311038 2848
rect 385678 2836 385684 2848
rect 311032 2808 385684 2836
rect 311032 2796 311038 2808
rect 385678 2796 385684 2808
rect 385736 2796 385742 2848
rect 395430 2796 395436 2848
rect 395488 2836 395494 2848
rect 416133 2839 416191 2845
rect 416133 2836 416145 2839
rect 395488 2808 416145 2836
rect 395488 2796 395494 2808
rect 416133 2805 416145 2808
rect 416179 2805 416191 2839
rect 416133 2799 416191 2805
rect 418157 2839 418215 2845
rect 418157 2805 418169 2839
rect 418203 2836 418215 2839
rect 427725 2839 427783 2845
rect 427725 2836 427737 2839
rect 418203 2808 427737 2836
rect 418203 2805 418215 2808
rect 418157 2799 418215 2805
rect 427725 2805 427737 2808
rect 427771 2805 427783 2839
rect 460198 2836 460204 2848
rect 427725 2799 427783 2805
rect 456076 2808 460204 2836
rect 456076 2780 456104 2808
rect 460198 2796 460204 2808
rect 460256 2796 460262 2848
rect 463234 2796 463240 2848
rect 463292 2836 463298 2848
rect 463602 2836 463608 2848
rect 463292 2808 463608 2836
rect 463292 2796 463298 2808
rect 463602 2796 463608 2808
rect 463660 2796 463666 2848
rect 471514 2796 471520 2848
rect 471572 2836 471578 2848
rect 471882 2836 471888 2848
rect 471572 2808 471888 2836
rect 471572 2796 471578 2808
rect 471882 2796 471888 2808
rect 471940 2796 471946 2848
rect 503714 2796 503720 2848
rect 503772 2836 503778 2848
rect 531038 2836 531044 2848
rect 503772 2808 531044 2836
rect 503772 2796 503778 2808
rect 531038 2796 531044 2808
rect 531096 2796 531102 2848
rect 542998 2796 543004 2848
rect 543056 2836 543062 2848
rect 547800 2836 547828 2944
rect 551186 2932 551192 2944
rect 551244 2932 551250 2984
rect 543056 2808 547828 2836
rect 543056 2796 543062 2808
rect 456058 2728 456064 2780
rect 456116 2728 456122 2780
rect 345474 688 345480 740
rect 345532 728 345538 740
rect 346302 728 346308 740
rect 345532 700 346308 728
rect 345532 688 345538 700
rect 346302 688 346308 700
rect 346360 688 346366 740
rect 139670 552 139676 604
rect 139728 592 139734 604
rect 140682 592 140688 604
rect 139728 564 140688 592
rect 139728 552 139734 564
rect 140682 552 140688 564
rect 140740 552 140746 604
rect 172974 552 172980 604
rect 173032 592 173038 604
rect 173802 592 173808 604
rect 173032 564 173808 592
rect 173032 552 173038 564
rect 173802 552 173808 564
rect 173860 552 173866 604
rect 180150 552 180156 604
rect 180208 592 180214 604
rect 180702 592 180708 604
rect 180208 564 180708 592
rect 180208 552 180214 564
rect 180702 552 180708 564
rect 180760 552 180766 604
rect 205082 552 205088 604
rect 205140 592 205146 604
rect 205542 592 205548 604
rect 205140 564 205548 592
rect 205140 552 205146 564
rect 205542 552 205548 564
rect 205600 552 205606 604
rect 206278 552 206284 604
rect 206336 592 206342 604
rect 206922 592 206928 604
rect 206336 564 206928 592
rect 206336 552 206342 564
rect 206922 552 206928 564
rect 206980 552 206986 604
rect 220538 552 220544 604
rect 220596 592 220602 604
rect 220722 592 220728 604
rect 220596 564 220728 592
rect 220596 552 220602 564
rect 220722 552 220728 564
rect 220780 552 220786 604
rect 393038 592 393044 604
rect 392999 564 393044 592
rect 393038 552 393044 564
rect 393096 552 393102 604
rect 413278 552 413284 604
rect 413336 592 413342 604
rect 414385 595 414443 601
rect 414385 592 414397 595
rect 413336 564 414397 592
rect 413336 552 413342 564
rect 414385 561 414397 564
rect 414431 561 414443 595
rect 414385 555 414443 561
rect 435818 552 435824 604
rect 435876 592 435882 604
rect 436002 592 436008 604
rect 435876 564 436008 592
rect 435876 552 435882 564
rect 436002 552 436008 564
rect 436060 552 436066 604
rect 453666 552 453672 604
rect 453724 592 453730 604
rect 453942 592 453948 604
rect 453724 564 453948 592
rect 453724 552 453730 564
rect 453942 552 453948 564
rect 454000 552 454006 604
rect 477770 552 477776 604
rect 477828 592 477834 604
rect 478690 592 478696 604
rect 477828 564 478696 592
rect 477828 552 477834 564
rect 478690 552 478696 564
rect 478748 552 478754 604
rect 480346 552 480352 604
rect 480404 592 480410 604
rect 481082 592 481088 604
rect 480404 564 481088 592
rect 480404 552 480410 564
rect 481082 552 481088 564
rect 481140 552 481146 604
rect 499758 552 499764 604
rect 499816 592 499822 604
rect 500126 592 500132 604
rect 499816 564 500132 592
rect 499816 552 499822 564
rect 500126 552 500132 564
rect 500184 552 500190 604
rect 506658 552 506664 604
rect 506716 592 506722 604
rect 507210 592 507216 604
rect 506716 564 507216 592
rect 506716 552 506722 564
rect 507210 552 507216 564
rect 507268 552 507274 604
rect 513558 552 513564 604
rect 513616 592 513622 604
rect 514386 592 514392 604
rect 513616 564 514392 592
rect 513616 552 513622 564
rect 514386 552 514392 564
rect 514444 552 514450 604
rect 520366 552 520372 604
rect 520424 592 520430 604
rect 521470 592 521476 604
rect 520424 564 521476 592
rect 520424 552 520430 564
rect 521470 552 521476 564
rect 521528 552 521534 604
<< via1 >>
rect 218980 700952 219032 701004
rect 393320 700952 393372 701004
rect 355968 700884 356020 700936
rect 543464 700884 543516 700936
rect 202788 700816 202840 700868
rect 390560 700816 390612 700868
rect 170312 700748 170364 700800
rect 396080 700748 396132 700800
rect 154120 700680 154172 700732
rect 401600 700680 401652 700732
rect 137836 700612 137888 700664
rect 398840 700612 398892 700664
rect 105452 700544 105504 700596
rect 404360 700544 404412 700596
rect 89168 700476 89220 700528
rect 409880 700476 409932 700528
rect 72976 700408 73028 700460
rect 407120 700408 407172 700460
rect 40500 700340 40552 700392
rect 411260 700340 411312 700392
rect 24308 700272 24360 700324
rect 416780 700272 416832 700324
rect 353208 700204 353260 700256
rect 527180 700204 527232 700256
rect 267648 700136 267700 700188
rect 383660 700136 383712 700188
rect 362868 700068 362920 700120
rect 478512 700068 478564 700120
rect 360108 700000 360160 700052
rect 462320 700000 462372 700052
rect 283840 699932 283892 699984
rect 385040 699932 385092 699984
rect 332508 699864 332560 699916
rect 375380 699864 375432 699916
rect 371148 699796 371200 699848
rect 413652 699796 413704 699848
rect 348792 699728 348844 699780
rect 378140 699728 378192 699780
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 364984 699660 365036 699712
rect 365628 699660 365680 699712
rect 368388 699660 368440 699712
rect 397460 699660 397512 699712
rect 344928 696940 344980 696992
rect 580172 696940 580224 696992
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 347688 685856 347740 685908
rect 580172 685856 580224 685908
rect 429292 684428 429344 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 419540 681708 419592 681760
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 342168 673480 342220 673532
rect 580172 673480 580224 673532
rect 269028 670692 269080 670744
rect 577504 670692 577556 670744
rect 3424 667904 3476 667956
rect 425060 667904 425112 667956
rect 429476 666587 429528 666596
rect 429476 666553 429485 666587
rect 429485 666553 429519 666587
rect 429519 666553 429528 666587
rect 429476 666544 429528 666553
rect 494152 666544 494204 666596
rect 559380 666544 559432 666596
rect 429292 656820 429344 656872
rect 559196 656863 559248 656872
rect 559196 656829 559205 656863
rect 559205 656829 559239 656863
rect 559239 656829 559248 656863
rect 559196 656820 559248 656829
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 422300 652740 422352 652792
rect 336648 650020 336700 650072
rect 580172 650020 580224 650072
rect 429200 647275 429252 647284
rect 429200 647241 429209 647275
rect 429209 647241 429243 647275
rect 429243 647241 429252 647275
rect 429200 647232 429252 647241
rect 559288 647232 559340 647284
rect 411260 645124 411312 645176
rect 412548 645124 412600 645176
rect 365168 643968 365220 644020
rect 429200 643968 429252 644020
rect 300768 643900 300820 643952
rect 380992 643900 381044 643952
rect 357348 643832 357400 643884
rect 494060 643832 494112 643884
rect 235908 643764 235960 643816
rect 388904 643764 388956 643816
rect 349436 643696 349488 643748
rect 559288 643696 559340 643748
rect 365628 643084 365680 643136
rect 373080 643084 373132 643136
rect 283656 643016 283708 643068
rect 427820 643016 427872 643068
rect 429016 643016 429068 643068
rect 523132 643016 523184 643068
rect 307300 642948 307352 643000
rect 473360 642948 473412 643000
rect 331036 642880 331088 642932
rect 532332 642880 532384 642932
rect 265164 642812 265216 642864
rect 320824 642812 320876 642864
rect 323124 642812 323176 642864
rect 532240 642812 532292 642864
rect 320456 642744 320508 642796
rect 530400 642744 530452 642796
rect 288900 642676 288952 642728
rect 307668 642676 307720 642728
rect 315212 642676 315264 642728
rect 532148 642676 532200 642728
rect 267832 642608 267884 642660
rect 269028 642608 269080 642660
rect 304632 642608 304684 642660
rect 532056 642608 532108 642660
rect 236276 642540 236328 642592
rect 290004 642540 290056 642592
rect 294144 642540 294196 642592
rect 531044 642540 531096 642592
rect 270500 642472 270552 642524
rect 530676 642472 530728 642524
rect 252008 642404 252060 642456
rect 263600 642404 263652 642456
rect 278320 642404 278372 642456
rect 580908 642404 580960 642456
rect 257344 642336 257396 642388
rect 580632 642336 580684 642388
rect 86224 642268 86276 642320
rect 438860 642268 438912 642320
rect 438952 642268 439004 642320
rect 454684 642268 454736 642320
rect 5448 642200 5500 642252
rect 433616 642200 433668 642252
rect 5356 642132 5408 642184
rect 441528 642132 441580 642184
rect 7932 642064 7984 642116
rect 446772 642064 446824 642116
rect 446864 642064 446916 642116
rect 486240 642064 486292 642116
rect 5264 641996 5316 642048
rect 449440 641996 449492 642048
rect 7656 641928 7708 641980
rect 462596 641928 462648 641980
rect 462964 641928 463016 641980
rect 502064 641928 502116 641980
rect 5172 641860 5224 641912
rect 465172 641860 465224 641912
rect 5080 641792 5132 641844
rect 473084 641792 473136 641844
rect 485136 641792 485188 641844
rect 517796 641792 517848 641844
rect 4988 641724 5040 641776
rect 488908 641724 488960 641776
rect 427820 641656 427872 641708
rect 580356 641656 580408 641708
rect 333612 641588 333664 641640
rect 530216 641588 530268 641640
rect 317788 641520 317840 641572
rect 529848 641520 529900 641572
rect 312544 641452 312596 641504
rect 530492 641452 530544 641504
rect 309968 641384 310020 641436
rect 529756 641384 529808 641436
rect 299388 641316 299440 641368
rect 531964 641316 532016 641368
rect 286232 641248 286284 641300
rect 530952 641248 531004 641300
rect 275744 641180 275796 641232
rect 530768 641180 530820 641232
rect 262588 641112 262640 641164
rect 530584 641112 530636 641164
rect 246764 641044 246816 641096
rect 529572 641044 529624 641096
rect 3976 640976 4028 641028
rect 258724 640976 258776 641028
rect 291476 640976 291528 641028
rect 580080 640976 580132 641028
rect 238852 640908 238904 640960
rect 529480 640908 529532 640960
rect 8208 640840 8260 640892
rect 428372 640840 428424 640892
rect 473360 640840 473412 640892
rect 579896 640840 579948 640892
rect 8116 640772 8168 640824
rect 431040 640772 431092 640824
rect 8024 640704 8076 640756
rect 436284 640704 436336 640756
rect 6552 640636 6604 640688
rect 444196 640772 444248 640824
rect 6460 640568 6512 640620
rect 452016 640568 452068 640620
rect 7748 640500 7800 640552
rect 459928 640500 459980 640552
rect 6368 640432 6420 640484
rect 467840 640432 467892 640484
rect 7564 640364 7616 640416
rect 475752 640364 475804 640416
rect 4804 640296 4856 640348
rect 515220 640296 515272 640348
rect 320824 640228 320876 640280
rect 580724 640228 580776 640280
rect 307668 640160 307720 640212
rect 579988 640160 580040 640212
rect 296812 640092 296864 640144
rect 531136 640092 531188 640144
rect 339224 640024 339276 640076
rect 580172 640024 580224 640076
rect 229744 639956 229796 640008
rect 478052 639956 478104 640008
rect 220912 639888 220964 639940
rect 235264 639888 235316 639940
rect 263600 639888 263652 639940
rect 580540 639888 580592 639940
rect 281264 639820 281316 639872
rect 530860 639820 530912 639872
rect 273168 639752 273220 639804
rect 580816 639752 580868 639804
rect 3332 639684 3384 639736
rect 438952 639684 439004 639736
rect 457076 639684 457128 639736
rect 4068 639616 4120 639668
rect 446864 639616 446916 639668
rect 7840 639548 7892 639600
rect 5540 639480 5592 639532
rect 23296 639480 23348 639532
rect 6276 639412 6328 639464
rect 156328 639480 156380 639532
rect 162676 639480 162728 639532
rect 201500 639480 201552 639532
rect 211068 639480 211120 639532
rect 480628 639616 480680 639668
rect 60648 639208 60700 639260
rect 66168 639208 66220 639260
rect 579804 639140 579856 639192
rect 580356 639140 580408 639192
rect 530216 627852 530268 627904
rect 579804 627852 579856 627904
rect 3240 624860 3292 624912
rect 8208 624860 8260 624912
rect 2780 610580 2832 610632
rect 5448 610580 5500 610632
rect 530308 604392 530360 604444
rect 579804 604392 579856 604444
rect 3240 596028 3292 596080
rect 8116 596028 8168 596080
rect 532332 593308 532384 593360
rect 579804 593308 579856 593360
rect 3240 567740 3292 567792
rect 8024 567740 8076 567792
rect 530400 557472 530452 557524
rect 579804 557472 579856 557524
rect 2780 553052 2832 553104
rect 5356 553052 5408 553104
rect 532240 546388 532292 546440
rect 579804 546388 579856 546440
rect 3240 539520 3292 539572
rect 86224 539520 86276 539572
rect 529848 534012 529900 534064
rect 579804 534012 579856 534064
rect 530492 510552 530544 510604
rect 579804 510552 579856 510604
rect 3240 510348 3292 510400
rect 6552 510348 6604 510400
rect 532148 499468 532200 499520
rect 579804 499468 579856 499520
rect 2780 496680 2832 496732
rect 5264 496680 5316 496732
rect 529756 487092 529808 487144
rect 579804 487092 579856 487144
rect 3240 481108 3292 481160
rect 7932 481108 7984 481160
rect 532056 463632 532108 463684
rect 579804 463632 579856 463684
rect 3148 452412 3200 452464
rect 6460 452412 6512 452464
rect 531228 440172 531280 440224
rect 579896 440172 579948 440224
rect 3148 438744 3200 438796
rect 7840 438744 7892 438796
rect 531136 416712 531188 416764
rect 579896 416712 579948 416764
rect 531964 405628 532016 405680
rect 579896 405628 579948 405680
rect 3148 395428 3200 395480
rect 7748 395428 7800 395480
rect 531044 393252 531096 393304
rect 579896 393252 579948 393304
rect 2780 380604 2832 380656
rect 5172 380604 5224 380656
rect 3332 366460 3384 366512
rect 7656 366460 7708 366512
rect 530952 346332 531004 346384
rect 579804 346332 579856 346384
rect 71044 338036 71096 338088
rect 264888 338036 264940 338088
rect 295800 338036 295852 338088
rect 332508 338036 332560 338088
rect 400220 338036 400272 338088
rect 405004 338036 405056 338088
rect 411812 338036 411864 338088
rect 412088 338036 412140 338088
rect 419172 338036 419224 338088
rect 427452 338036 427504 338088
rect 445484 338036 445536 338088
rect 451740 338036 451792 338088
rect 490840 338036 490892 338088
rect 509148 338036 509200 338088
rect 542360 338036 542412 338088
rect 66904 337968 66956 338020
rect 261208 337968 261260 338020
rect 322756 337968 322808 338020
rect 395252 337968 395304 338020
rect 3240 337900 3292 337952
rect 6368 337900 6420 337952
rect 57244 337900 57296 337952
rect 257528 337900 257580 337952
rect 309784 337900 309836 337952
rect 50344 337832 50396 337884
rect 251364 337832 251416 337884
rect 268384 337832 268436 337884
rect 288716 337832 288768 337884
rect 311900 337832 311952 337884
rect 312268 337832 312320 337884
rect 313464 337832 313516 337884
rect 314108 337832 314160 337884
rect 314660 337832 314712 337884
rect 315396 337832 315448 337884
rect 316040 337900 316092 337952
rect 316684 337900 316736 337952
rect 317604 337900 317656 337952
rect 318340 337900 318392 337952
rect 320180 337900 320232 337952
rect 320916 337900 320968 337952
rect 385684 337900 385736 337952
rect 389732 337900 389784 337952
rect 402612 337968 402664 338020
rect 416688 337968 416740 338020
rect 443644 337968 443696 338020
rect 407764 337900 407816 337952
rect 415492 337900 415544 337952
rect 416044 337900 416096 337952
rect 443000 337900 443052 337952
rect 387984 337832 388036 337884
rect 391204 337832 391256 337884
rect 397092 337832 397144 337884
rect 441252 337832 441304 337884
rect 450360 337968 450412 338020
rect 451924 337968 451976 338020
rect 459008 337968 459060 338020
rect 477316 337968 477368 338020
rect 480260 337968 480312 338020
rect 498752 337968 498804 338020
rect 499488 337968 499540 338020
rect 512828 337968 512880 338020
rect 547144 337968 547196 338020
rect 490196 337900 490248 337952
rect 501604 337900 501656 337952
rect 503444 337900 503496 337952
rect 503628 337900 503680 337952
rect 512276 337900 512328 337952
rect 547236 337900 547288 337952
rect 451004 337832 451056 337884
rect 453304 337832 453356 337884
rect 462044 337832 462096 337884
rect 463608 337832 463660 337884
rect 468116 337832 468168 337884
rect 487160 337832 487212 337884
rect 499764 337832 499816 337884
rect 501236 337832 501288 337884
rect 46204 337764 46256 337816
rect 247684 337764 247736 337816
rect 269764 337764 269816 337816
rect 292396 337764 292448 337816
rect 294604 337764 294656 337816
rect 375104 337764 375156 337816
rect 375288 337764 375340 337816
rect 39304 337696 39356 337748
rect 240416 337696 240468 337748
rect 248420 337696 248472 337748
rect 249524 337696 249576 337748
rect 249984 337696 250036 337748
rect 250812 337696 250864 337748
rect 258724 337696 258776 337748
rect 266728 337696 266780 337748
rect 287704 337696 287756 337748
rect 373264 337696 373316 337748
rect 376024 337696 376076 337748
rect 406292 337764 406344 337816
rect 409788 337764 409840 337816
rect 439964 337764 440016 337816
rect 445024 337764 445076 337816
rect 456524 337764 456576 337816
rect 464988 337764 465040 337816
rect 468760 337764 468812 337816
rect 482836 337764 482888 337816
rect 497556 337764 497608 337816
rect 509884 337764 509936 337816
rect 409972 337696 410024 337748
rect 412548 337696 412600 337748
rect 441804 337696 441856 337748
rect 442356 337696 442408 337748
rect 454684 337696 454736 337748
rect 456064 337696 456116 337748
rect 463884 337696 463936 337748
rect 477960 337696 478012 337748
rect 478788 337696 478840 337748
rect 479156 337696 479208 337748
rect 32404 337628 32456 337680
rect 264336 337628 264388 337680
rect 281448 337628 281500 337680
rect 283564 337628 283616 337680
rect 365904 337628 365956 337680
rect 366916 337628 366968 337680
rect 418528 337628 418580 337680
rect 420828 337628 420880 337680
rect 446128 337628 446180 337680
rect 449256 337628 449308 337680
rect 457168 337628 457220 337680
rect 466368 337628 466420 337680
rect 469404 337628 469456 337680
rect 475476 337628 475528 337680
rect 477592 337628 477644 337680
rect 480352 337696 480404 337748
rect 481548 337696 481600 337748
rect 489000 337696 489052 337748
rect 28264 337560 28316 337612
rect 17224 337492 17276 337544
rect 228180 337492 228232 337544
rect 234896 337492 234948 337544
rect 248328 337560 248380 337612
rect 244648 337492 244700 337544
rect 246304 337492 246356 337544
rect 290004 337560 290056 337612
rect 293868 337560 293920 337612
rect 380624 337560 380676 337612
rect 391572 337560 391624 337612
rect 393136 337560 393188 337612
rect 432052 337560 432104 337612
rect 262864 337492 262916 337544
rect 285036 337492 285088 337544
rect 286968 337492 287020 337544
rect 376944 337492 376996 337544
rect 24124 337424 24176 337476
rect 15844 337356 15896 337408
rect 228180 337356 228232 337408
rect 235448 337356 235500 337408
rect 261484 337424 261536 337476
rect 239772 337356 239824 337408
rect 257344 337356 257396 337408
rect 263048 337356 263100 337408
rect 61384 337288 61436 337340
rect 252008 337288 252060 337340
rect 255964 337288 256016 337340
rect 259368 337288 259420 337340
rect 264244 337424 264296 337476
rect 279608 337424 279660 337476
rect 280068 337424 280120 337476
rect 369584 337424 369636 337476
rect 384028 337492 384080 337544
rect 275928 337356 275980 337408
rect 276664 337356 276716 337408
rect 371424 337356 371476 337408
rect 372528 337356 372580 337408
rect 389088 337492 389140 337544
rect 413468 337424 413520 337476
rect 420368 337424 420420 337476
rect 421012 337356 421064 337408
rect 429108 337492 429160 337544
rect 434628 337560 434680 337612
rect 452844 337560 452896 337612
rect 453948 337560 454000 337612
rect 463240 337560 463292 337612
rect 478512 337560 478564 337612
rect 483204 337560 483256 337612
rect 483480 337628 483532 337680
rect 484216 337628 484268 337680
rect 485872 337628 485924 337680
rect 489184 337628 489236 337680
rect 491392 337628 491444 337680
rect 492588 337628 492640 337680
rect 493232 337628 493284 337680
rect 493968 337628 494020 337680
rect 484584 337560 484636 337612
rect 492680 337560 492732 337612
rect 495716 337560 495768 337612
rect 496728 337560 496780 337612
rect 496912 337628 496964 337680
rect 498844 337628 498896 337680
rect 499948 337696 500000 337748
rect 500776 337696 500828 337748
rect 502616 337696 502668 337748
rect 504272 337696 504324 337748
rect 505008 337696 505060 337748
rect 505468 337696 505520 337748
rect 506388 337696 506440 337748
rect 506756 337696 506808 337748
rect 507768 337696 507820 337748
rect 507952 337696 508004 337748
rect 509148 337696 509200 337748
rect 510988 337696 511040 337748
rect 511908 337696 511960 337748
rect 502432 337628 502484 337680
rect 503536 337628 503588 337680
rect 514668 337832 514720 337884
rect 515864 337764 515916 337816
rect 520832 337832 520884 337884
rect 556804 337832 556856 337884
rect 516508 337696 516560 337748
rect 517428 337696 517480 337748
rect 553400 337764 553452 337816
rect 554872 337696 554924 337748
rect 516784 337628 516836 337680
rect 518348 337628 518400 337680
rect 560300 337628 560352 337680
rect 510804 337560 510856 337612
rect 517704 337560 517756 337612
rect 518808 337560 518860 337612
rect 518992 337560 519044 337612
rect 520096 337560 520148 337612
rect 522028 337560 522080 337612
rect 446680 337492 446732 337544
rect 451188 337492 451240 337544
rect 461400 337492 461452 337544
rect 479800 337492 479852 337544
rect 446404 337424 446456 337476
rect 458364 337424 458416 337476
rect 429568 337356 429620 337408
rect 430488 337356 430540 337408
rect 447324 337356 447376 337408
rect 448428 337356 448480 337408
rect 460204 337356 460256 337408
rect 460848 337356 460900 337408
rect 466920 337356 466972 337408
rect 270408 337288 270460 337340
rect 284944 337288 284996 337340
rect 338948 337288 339000 337340
rect 365720 337288 365772 337340
rect 378508 337288 378560 337340
rect 403900 337288 403952 337340
rect 409144 337288 409196 337340
rect 428372 337288 428424 337340
rect 428556 337288 428608 337340
rect 442264 337288 442316 337340
rect 449808 337288 449860 337340
rect 481640 337492 481692 337544
rect 482836 337492 482888 337544
rect 494520 337492 494572 337544
rect 513564 337492 513616 337544
rect 513840 337492 513892 337544
rect 563152 337560 563204 337612
rect 567200 337492 567252 337544
rect 480996 337424 481048 337476
rect 485044 337424 485096 337476
rect 485320 337424 485372 337476
rect 493324 337424 493376 337476
rect 496268 337424 496320 337476
rect 517612 337424 517664 337476
rect 519544 337424 519596 337476
rect 484676 337356 484728 337408
rect 485688 337356 485740 337408
rect 491484 337356 491536 337408
rect 498108 337356 498160 337408
rect 520372 337356 520424 337408
rect 523224 337356 523276 337408
rect 569224 337424 569276 337476
rect 526904 337356 526956 337408
rect 571984 337356 572036 337408
rect 485964 337288 486016 337340
rect 506664 337288 506716 337340
rect 517152 337288 517204 337340
rect 549904 337288 549956 337340
rect 84844 337220 84896 337272
rect 272248 337220 272300 337272
rect 283656 337220 283708 337272
rect 337108 337220 337160 337272
rect 339408 337220 339460 337272
rect 97264 337152 97316 337204
rect 277768 337152 277820 337204
rect 316684 337152 316736 337204
rect 346308 337220 346360 337272
rect 407488 337220 407540 337272
rect 104808 337084 104860 337136
rect 283196 337084 283248 337136
rect 353208 337152 353260 337204
rect 411168 337152 411220 337204
rect 413376 337220 413428 337272
rect 417332 337152 417384 337204
rect 417608 337152 417660 337204
rect 422208 337220 422260 337272
rect 424968 337220 425020 337272
rect 447968 337220 448020 337272
rect 508596 337220 508648 337272
rect 540244 337220 540296 337272
rect 424048 337152 424100 337204
rect 433248 337152 433300 337204
rect 449164 337152 449216 337204
rect 453396 337152 453448 337204
rect 460756 337152 460808 337204
rect 515312 337152 515364 337204
rect 526812 337152 526864 337204
rect 528744 337152 528796 337204
rect 529756 337152 529808 337204
rect 558184 337152 558236 337204
rect 357348 337084 357400 337136
rect 413652 337084 413704 337136
rect 414664 337084 414716 337136
rect 422852 337084 422904 337136
rect 423588 337084 423640 337136
rect 111708 337016 111760 337068
rect 286876 337016 286928 337068
rect 360108 337016 360160 337068
rect 414848 337016 414900 337068
rect 420276 337016 420328 337068
rect 431868 337016 431920 337068
rect 451648 337084 451700 337136
rect 507308 337084 507360 337136
rect 538220 337084 538272 337136
rect 436008 337016 436060 337068
rect 454040 337016 454092 337068
rect 487712 337016 487764 337068
rect 488448 337016 488500 337068
rect 495072 337016 495124 337068
rect 496084 337016 496136 337068
rect 509792 337016 509844 337068
rect 540336 337016 540388 337068
rect 118608 336948 118660 337000
rect 290556 336948 290608 337000
rect 366364 336948 366416 337000
rect 410524 336948 410576 337000
rect 416412 336948 416464 337000
rect 420184 336948 420236 337000
rect 125508 336880 125560 336932
rect 294236 336880 294288 336932
rect 363696 336880 363748 336932
rect 105544 336812 105596 336864
rect 274088 336812 274140 336864
rect 366456 336812 366508 336864
rect 395436 336880 395488 336932
rect 400772 336880 400824 336932
rect 421932 336880 421984 336932
rect 424416 336948 424468 337000
rect 398932 336812 398984 336864
rect 106924 336744 106976 336796
rect 268568 336744 268620 336796
rect 363604 336744 363656 336796
rect 374644 336744 374696 336796
rect 381544 336744 381596 336796
rect 382464 336744 382516 336796
rect 382924 336744 382976 336796
rect 386144 336744 386196 336796
rect 389916 336744 389968 336796
rect 393412 336744 393464 336796
rect 396724 336744 396776 336796
rect 404452 336812 404504 336864
rect 413284 336812 413336 336864
rect 401048 336744 401100 336796
rect 408132 336744 408184 336796
rect 410616 336744 410668 336796
rect 413008 336744 413060 336796
rect 416136 336744 416188 336796
rect 424692 336812 424744 336864
rect 427084 336880 427136 336932
rect 438768 336948 438820 337000
rect 503444 336948 503496 337000
rect 545764 336948 545816 337000
rect 431224 336812 431276 336864
rect 440608 336880 440660 336932
rect 435364 336812 435416 336864
rect 442448 336812 442500 336864
rect 424324 336744 424376 336796
rect 425888 336744 425940 336796
rect 432604 336744 432656 336796
rect 435732 336744 435784 336796
rect 436928 336744 436980 336796
rect 438124 336744 438176 336796
rect 444288 336744 444340 336796
rect 446496 336744 446548 336796
rect 453488 336880 453540 336932
rect 460204 336880 460256 336932
rect 464436 336880 464488 336932
rect 476120 336880 476172 336932
rect 477776 336880 477828 336932
rect 504916 336880 504968 336932
rect 534080 336880 534132 336932
rect 464344 336812 464396 336864
rect 466276 336812 466328 336864
rect 467748 336812 467800 336864
rect 469956 336812 470008 336864
rect 543004 336812 543056 336864
rect 447784 336744 447836 336796
rect 455328 336744 455380 336796
rect 457444 336744 457496 336796
rect 462596 336744 462648 336796
rect 464436 336744 464488 336796
rect 465724 336744 465776 336796
rect 469864 336744 469916 336796
rect 471244 336744 471296 336796
rect 474924 336744 474976 336796
rect 476028 336744 476080 336796
rect 356796 336676 356848 336728
rect 370504 336676 370556 336728
rect 375748 336676 375800 336728
rect 380992 336676 381044 336728
rect 381360 336676 381412 336728
rect 524512 336744 524564 336796
rect 525616 336744 525668 336796
rect 527548 336744 527600 336796
rect 528468 336744 528520 336796
rect 529388 336744 529440 336796
rect 529848 336744 529900 336796
rect 531320 336744 531372 336796
rect 252560 336268 252612 336320
rect 253848 336268 253900 336320
rect 229100 335588 229152 335640
rect 229836 335588 229888 335640
rect 230480 335588 230532 335640
rect 230940 335588 230992 335640
rect 241520 335588 241572 335640
rect 241980 335588 242032 335640
rect 259644 335588 259696 335640
rect 260288 335588 260340 335640
rect 296812 335588 296864 335640
rect 297548 335588 297600 335640
rect 299480 335588 299532 335640
rect 300124 335588 300176 335640
rect 302332 335588 302384 335640
rect 303068 335588 303120 335640
rect 303620 335588 303672 335640
rect 304356 335588 304408 335640
rect 306380 335588 306432 335640
rect 306748 335588 306800 335640
rect 307852 335588 307904 335640
rect 308036 335588 308088 335640
rect 310704 335588 310756 335640
rect 311164 335588 311216 335640
rect 323124 335588 323176 335640
rect 323860 335588 323912 335640
rect 328644 335588 328696 335640
rect 329380 335588 329432 335640
rect 335360 335588 335412 335640
rect 336188 335588 336240 335640
rect 339500 335588 339552 335640
rect 340420 335588 340472 335640
rect 345020 335588 345072 335640
rect 345940 335588 345992 335640
rect 350540 335588 350592 335640
rect 351460 335588 351512 335640
rect 354680 335588 354732 335640
rect 355140 335588 355192 335640
rect 357624 335588 357676 335640
rect 358268 335588 358320 335640
rect 360200 335588 360252 335640
rect 360660 335588 360712 335640
rect 361672 335588 361724 335640
rect 362500 335588 362552 335640
rect 367192 335588 367244 335640
rect 368020 335588 368072 335640
rect 378232 335588 378284 335640
rect 379060 335588 379112 335640
rect 405924 335588 405976 335640
rect 406660 335588 406712 335640
rect 422300 335588 422352 335640
rect 423220 335588 423272 335640
rect 430580 335588 430632 335640
rect 431132 335588 431184 335640
rect 470692 335588 470744 335640
rect 471428 335588 471480 335640
rect 245660 335520 245712 335572
rect 246488 335520 246540 335572
rect 334072 335384 334124 335436
rect 357624 335291 357676 335300
rect 357624 335257 357633 335291
rect 357633 335257 357667 335291
rect 357667 335257 357676 335291
rect 357624 335248 357676 335257
rect 334164 335180 334216 335232
rect 254124 335112 254176 335164
rect 255044 335112 255096 335164
rect 340880 334568 340932 334620
rect 341708 334568 341760 334620
rect 251824 334364 251876 334416
rect 253204 334364 253256 334416
rect 362960 334364 363012 334416
rect 363788 334364 363840 334416
rect 253204 334228 253256 334280
rect 255688 334228 255740 334280
rect 294052 333931 294104 333940
rect 294052 333897 294061 333931
rect 294061 333897 294095 333931
rect 294095 333897 294104 333931
rect 294052 333888 294104 333897
rect 237472 333616 237524 333668
rect 238300 333616 238352 333668
rect 324412 333276 324464 333328
rect 325056 333276 325108 333328
rect 433708 333276 433760 333328
rect 434168 333276 434220 333328
rect 466552 333276 466604 333328
rect 467104 333276 467156 333328
rect 325700 332732 325752 332784
rect 326436 332732 326488 332784
rect 359096 331848 359148 331900
rect 359280 331848 359332 331900
rect 349160 331780 349212 331832
rect 349620 331780 349672 331832
rect 333980 331576 334032 331628
rect 334256 331576 334308 331628
rect 343640 331508 343692 331560
rect 344100 331508 344152 331560
rect 364524 331372 364576 331424
rect 364984 331372 365036 331424
rect 231952 331236 232004 331288
rect 232780 331236 232832 331288
rect 309692 331236 309744 331288
rect 342628 331279 342680 331288
rect 342628 331245 342637 331279
rect 342637 331245 342671 331279
rect 342671 331245 342680 331279
rect 342628 331236 342680 331245
rect 393136 331279 393188 331288
rect 393136 331245 393145 331279
rect 393145 331245 393179 331279
rect 393179 331245 393188 331279
rect 393136 331236 393188 331245
rect 305184 331168 305236 331220
rect 416780 331168 416832 331220
rect 416964 331168 417016 331220
rect 422300 331168 422352 331220
rect 422484 331168 422536 331220
rect 305276 331100 305328 331152
rect 451556 330488 451608 330540
rect 292764 328992 292816 329044
rect 293224 328992 293276 329044
rect 241796 328448 241848 328500
rect 242440 328448 242492 328500
rect 265256 328448 265308 328500
rect 265532 328448 265584 328500
rect 267096 328448 267148 328500
rect 270776 328448 270828 328500
rect 271052 328448 271104 328500
rect 295616 328491 295668 328500
rect 295616 328457 295625 328491
rect 295625 328457 295659 328491
rect 295659 328457 295668 328491
rect 295616 328448 295668 328457
rect 309416 328491 309468 328500
rect 309416 328457 309425 328491
rect 309425 328457 309459 328491
rect 309459 328457 309468 328491
rect 309416 328448 309468 328457
rect 330024 328448 330076 328500
rect 330576 328448 330628 328500
rect 331496 328448 331548 328500
rect 331680 328448 331732 328500
rect 332692 328448 332744 328500
rect 332968 328448 333020 328500
rect 334440 328448 334492 328500
rect 334808 328448 334860 328500
rect 336924 328448 336976 328500
rect 337200 328448 337252 328500
rect 342628 328491 342680 328500
rect 342628 328457 342637 328491
rect 342637 328457 342671 328491
rect 342671 328457 342680 328491
rect 342628 328448 342680 328457
rect 397736 328448 397788 328500
rect 397920 328448 397972 328500
rect 252652 328423 252704 328432
rect 252652 328389 252661 328423
rect 252661 328389 252695 328423
rect 252695 328389 252704 328423
rect 252652 328380 252704 328389
rect 416964 328380 417016 328432
rect 422484 328380 422536 328432
rect 428004 328380 428056 328432
rect 433708 328423 433760 328432
rect 433708 328389 433717 328423
rect 433717 328389 433751 328423
rect 433751 328389 433760 328423
rect 433708 328380 433760 328389
rect 472164 328380 472216 328432
rect 236276 327088 236328 327140
rect 236920 327088 236972 327140
rect 370044 327131 370096 327140
rect 370044 327097 370053 327131
rect 370053 327097 370087 327131
rect 370087 327097 370096 327131
rect 370044 327088 370096 327097
rect 375564 327131 375616 327140
rect 375564 327097 375573 327131
rect 375573 327097 375607 327131
rect 375607 327097 375616 327131
rect 375564 327088 375616 327097
rect 393044 327088 393096 327140
rect 292764 327063 292816 327072
rect 292764 327029 292773 327063
rect 292773 327029 292807 327063
rect 292807 327029 292816 327063
rect 292764 327020 292816 327029
rect 318984 326179 319036 326188
rect 318984 326145 318993 326179
rect 318993 326145 319027 326179
rect 319027 326145 319036 326179
rect 318984 326136 319036 326145
rect 357624 325839 357676 325848
rect 357624 325805 357633 325839
rect 357633 325805 357667 325839
rect 357667 325805 357676 325839
rect 357624 325796 357676 325805
rect 356520 325703 356572 325712
rect 356520 325669 356529 325703
rect 356529 325669 356563 325703
rect 356563 325669 356572 325703
rect 356520 325660 356572 325669
rect 230664 325567 230716 325576
rect 230664 325533 230673 325567
rect 230673 325533 230707 325567
rect 230707 325533 230716 325567
rect 230664 325524 230716 325533
rect 393044 324164 393096 324216
rect 2780 323552 2832 323604
rect 5080 323552 5132 323604
rect 530860 322872 530912 322924
rect 580080 322872 580132 322924
rect 249984 321691 250036 321700
rect 249984 321657 249993 321691
rect 249993 321657 250027 321691
rect 250027 321657 250036 321691
rect 249984 321648 250036 321657
rect 261024 321648 261076 321700
rect 231952 321580 232004 321632
rect 259736 321580 259788 321632
rect 324504 321580 324556 321632
rect 359096 321580 359148 321632
rect 392216 321580 392268 321632
rect 408684 321580 408736 321632
rect 466552 321623 466604 321632
rect 466552 321589 466561 321623
rect 466561 321589 466595 321623
rect 466595 321589 466604 321623
rect 466552 321580 466604 321589
rect 261024 321512 261076 321564
rect 324412 321512 324464 321564
rect 400404 321512 400456 321564
rect 400588 321512 400640 321564
rect 232044 321444 232096 321496
rect 408776 321444 408828 321496
rect 252652 320127 252704 320136
rect 252652 320093 252661 320127
rect 252661 320093 252695 320127
rect 252695 320093 252704 320127
rect 252652 320084 252704 320093
rect 230848 318792 230900 318844
rect 259644 318835 259696 318844
rect 259644 318801 259653 318835
rect 259653 318801 259687 318835
rect 259687 318801 259696 318835
rect 259644 318792 259696 318801
rect 359004 318835 359056 318844
rect 359004 318801 359013 318835
rect 359013 318801 359047 318835
rect 359047 318801 359056 318835
rect 359004 318792 359056 318801
rect 392124 318835 392176 318844
rect 392124 318801 392133 318835
rect 392133 318801 392167 318835
rect 392167 318801 392176 318835
rect 392124 318792 392176 318801
rect 416872 318835 416924 318844
rect 416872 318801 416881 318835
rect 416881 318801 416915 318835
rect 416915 318801 416924 318835
rect 416872 318792 416924 318801
rect 422392 318835 422444 318844
rect 422392 318801 422401 318835
rect 422401 318801 422435 318835
rect 422435 318801 422444 318835
rect 422392 318792 422444 318801
rect 427912 318835 427964 318844
rect 427912 318801 427921 318835
rect 427921 318801 427955 318835
rect 427955 318801 427964 318835
rect 427912 318792 427964 318801
rect 433800 318792 433852 318844
rect 466552 318835 466604 318844
rect 466552 318801 466561 318835
rect 466561 318801 466595 318835
rect 466595 318801 466604 318835
rect 466552 318792 466604 318801
rect 472072 318835 472124 318844
rect 472072 318801 472081 318835
rect 472081 318801 472115 318835
rect 472115 318801 472124 318835
rect 472072 318792 472124 318801
rect 283012 318724 283064 318776
rect 283104 318724 283156 318776
rect 288624 318767 288676 318776
rect 288624 318733 288633 318767
rect 288633 318733 288667 318767
rect 288667 318733 288676 318767
rect 288624 318724 288676 318733
rect 327264 318767 327316 318776
rect 327264 318733 327273 318767
rect 327273 318733 327307 318767
rect 327307 318733 327316 318767
rect 327264 318724 327316 318733
rect 332784 318767 332836 318776
rect 332784 318733 332793 318767
rect 332793 318733 332827 318767
rect 332827 318733 332836 318767
rect 332784 318724 332836 318733
rect 347964 318724 348016 318776
rect 348056 318724 348108 318776
rect 352012 318724 352064 318776
rect 353484 318724 353536 318776
rect 353576 318724 353628 318776
rect 371424 318724 371476 318776
rect 375564 318724 375616 318776
rect 375748 318724 375800 318776
rect 376944 318724 376996 318776
rect 381084 318724 381136 318776
rect 381268 318724 381320 318776
rect 382280 318724 382332 318776
rect 382464 318724 382516 318776
rect 387892 318724 387944 318776
rect 387984 318724 388036 318776
rect 397736 318767 397788 318776
rect 397736 318733 397745 318767
rect 397745 318733 397779 318767
rect 397779 318733 397788 318767
rect 397736 318724 397788 318733
rect 352104 318656 352156 318708
rect 249984 317475 250036 317484
rect 249984 317441 249993 317475
rect 249993 317441 250027 317475
rect 250027 317441 250036 317475
rect 249984 317432 250036 317441
rect 292764 317475 292816 317484
rect 292764 317441 292773 317475
rect 292773 317441 292807 317475
rect 292807 317441 292816 317475
rect 292764 317432 292816 317441
rect 319168 317432 319220 317484
rect 255412 317364 255464 317416
rect 255596 317364 255648 317416
rect 283012 317364 283064 317416
rect 283288 317364 283340 317416
rect 375748 317407 375800 317416
rect 375748 317373 375757 317407
rect 375757 317373 375791 317407
rect 375791 317373 375800 317407
rect 375748 317364 375800 317373
rect 381268 317407 381320 317416
rect 381268 317373 381277 317407
rect 381277 317373 381311 317407
rect 381311 317373 381320 317407
rect 381268 317364 381320 317373
rect 382280 317407 382332 317416
rect 382280 317373 382289 317407
rect 382289 317373 382323 317407
rect 382323 317373 382332 317407
rect 382280 317364 382332 317373
rect 387892 317407 387944 317416
rect 387892 317373 387901 317407
rect 387901 317373 387935 317407
rect 387935 317373 387944 317407
rect 387892 317364 387944 317373
rect 451556 316072 451608 316124
rect 451740 316072 451792 316124
rect 277676 316004 277728 316056
rect 277860 316004 277912 316056
rect 294144 316004 294196 316056
rect 357532 316004 357584 316056
rect 357808 316004 357860 316056
rect 232044 315936 232096 315988
rect 356520 315979 356572 315988
rect 356520 315945 356529 315979
rect 356529 315945 356563 315979
rect 356563 315945 356572 315979
rect 356520 315936 356572 315945
rect 451556 315979 451608 315988
rect 451556 315945 451565 315979
rect 451565 315945 451599 315979
rect 451599 315945 451608 315979
rect 451556 315936 451608 315945
rect 397736 312171 397788 312180
rect 397736 312137 397745 312171
rect 397745 312137 397779 312171
rect 397779 312137 397788 312171
rect 397736 312128 397788 312137
rect 294144 311924 294196 311976
rect 230664 311856 230716 311908
rect 230848 311856 230900 311908
rect 249984 311856 250036 311908
rect 277584 311899 277636 311908
rect 277584 311865 277593 311899
rect 277593 311865 277627 311899
rect 277627 311865 277636 311899
rect 277584 311856 277636 311865
rect 433432 311856 433484 311908
rect 433800 311856 433852 311908
rect 249892 311788 249944 311840
rect 294144 311788 294196 311840
rect 346584 311831 346636 311840
rect 346584 311797 346593 311831
rect 346593 311797 346627 311831
rect 346627 311797 346636 311831
rect 346584 311788 346636 311797
rect 416780 311788 416832 311840
rect 416964 311788 417016 311840
rect 422300 311788 422352 311840
rect 422484 311788 422536 311840
rect 427820 311788 427872 311840
rect 428004 311788 428056 311840
rect 466460 311788 466512 311840
rect 466644 311788 466696 311840
rect 471980 311788 472032 311840
rect 472164 311788 472216 311840
rect 371332 309315 371384 309324
rect 371332 309281 371341 309315
rect 371341 309281 371375 309315
rect 371375 309281 371384 309315
rect 371332 309272 371384 309281
rect 376852 309315 376904 309324
rect 376852 309281 376861 309315
rect 376861 309281 376895 309315
rect 376895 309281 376904 309315
rect 376852 309272 376904 309281
rect 252560 309136 252612 309188
rect 252744 309136 252796 309188
rect 267096 309179 267148 309188
rect 267096 309145 267105 309179
rect 267105 309145 267139 309179
rect 267139 309145 267148 309179
rect 267096 309136 267148 309145
rect 287152 309136 287204 309188
rect 287244 309136 287296 309188
rect 288624 309179 288676 309188
rect 288624 309145 288633 309179
rect 288633 309145 288667 309179
rect 288667 309145 288676 309179
rect 288624 309136 288676 309145
rect 305184 309136 305236 309188
rect 305276 309136 305328 309188
rect 319168 309204 319220 309256
rect 342628 309204 342680 309256
rect 324228 309136 324280 309188
rect 324504 309136 324556 309188
rect 327264 309179 327316 309188
rect 327264 309145 327273 309179
rect 327273 309145 327307 309179
rect 327307 309145 327316 309179
rect 327264 309136 327316 309145
rect 332784 309179 332836 309188
rect 332784 309145 332793 309179
rect 332793 309145 332827 309179
rect 332827 309145 332836 309179
rect 332784 309136 332836 309145
rect 334440 309179 334492 309188
rect 334440 309145 334449 309179
rect 334449 309145 334483 309179
rect 334483 309145 334492 309179
rect 334440 309136 334492 309145
rect 336832 309136 336884 309188
rect 336924 309136 336976 309188
rect 342444 309136 342496 309188
rect 346584 309179 346636 309188
rect 346584 309145 346593 309179
rect 346593 309145 346627 309179
rect 346627 309145 346636 309179
rect 346584 309136 346636 309145
rect 393228 309179 393280 309188
rect 393228 309145 393237 309179
rect 393237 309145 393271 309179
rect 393271 309145 393280 309179
rect 393228 309136 393280 309145
rect 400312 309136 400364 309188
rect 400404 309136 400456 309188
rect 236276 309068 236328 309120
rect 236368 309068 236420 309120
rect 270684 309111 270736 309120
rect 270684 309077 270693 309111
rect 270693 309077 270727 309111
rect 270727 309077 270736 309111
rect 270684 309068 270736 309077
rect 309324 309111 309376 309120
rect 309324 309077 309333 309111
rect 309333 309077 309367 309111
rect 309367 309077 309376 309111
rect 309324 309068 309376 309077
rect 318984 309068 319036 309120
rect 375748 309111 375800 309120
rect 375748 309077 375757 309111
rect 375757 309077 375791 309111
rect 375791 309077 375800 309111
rect 375748 309068 375800 309077
rect 376852 309111 376904 309120
rect 376852 309077 376861 309111
rect 376861 309077 376895 309111
rect 376895 309077 376904 309111
rect 376852 309068 376904 309077
rect 416964 309068 417016 309120
rect 422484 309111 422536 309120
rect 422484 309077 422493 309111
rect 422493 309077 422527 309111
rect 422527 309077 422536 309111
rect 422484 309068 422536 309077
rect 428004 309111 428056 309120
rect 428004 309077 428013 309111
rect 428013 309077 428047 309111
rect 428047 309077 428056 309111
rect 428004 309068 428056 309077
rect 433432 309111 433484 309120
rect 433432 309077 433441 309111
rect 433441 309077 433475 309111
rect 433475 309077 433484 309111
rect 433432 309068 433484 309077
rect 466644 309068 466696 309120
rect 472164 309068 472216 309120
rect 342444 309043 342496 309052
rect 342444 309009 342453 309043
rect 342453 309009 342487 309043
rect 342487 309009 342496 309043
rect 342444 309000 342496 309009
rect 261024 307776 261076 307828
rect 261116 307776 261168 307828
rect 267096 307819 267148 307828
rect 267096 307785 267105 307819
rect 267105 307785 267139 307819
rect 267139 307785 267148 307819
rect 267096 307776 267148 307785
rect 334440 307819 334492 307828
rect 334440 307785 334449 307819
rect 334449 307785 334483 307819
rect 334483 307785 334492 307819
rect 334440 307776 334492 307785
rect 381268 307819 381320 307828
rect 381268 307785 381277 307819
rect 381277 307785 381311 307819
rect 381311 307785 381320 307819
rect 381268 307776 381320 307785
rect 387892 307819 387944 307828
rect 387892 307785 387901 307819
rect 387901 307785 387935 307819
rect 387935 307785 387944 307819
rect 387892 307776 387944 307785
rect 243084 307708 243136 307760
rect 292764 307751 292816 307760
rect 292764 307717 292773 307751
rect 292773 307717 292807 307751
rect 292807 307717 292816 307751
rect 292764 307708 292816 307717
rect 277584 306391 277636 306400
rect 277584 306357 277593 306391
rect 277593 306357 277627 306391
rect 277627 306357 277636 306391
rect 277584 306348 277636 306357
rect 357532 306348 357584 306400
rect 357624 306348 357676 306400
rect 365812 306348 365864 306400
rect 365996 306348 366048 306400
rect 387892 304895 387944 304904
rect 387892 304861 387901 304895
rect 387901 304861 387935 304895
rect 387935 304861 387944 304895
rect 387892 304852 387944 304861
rect 230664 304283 230716 304292
rect 230664 304249 230673 304283
rect 230673 304249 230707 304283
rect 230707 304249 230716 304283
rect 230664 304240 230716 304249
rect 298284 302268 298336 302320
rect 347964 302268 348016 302320
rect 400404 302268 400456 302320
rect 347964 302132 348016 302184
rect 298376 302064 298428 302116
rect 382464 302064 382516 302116
rect 408776 302243 408828 302252
rect 408776 302209 408785 302243
rect 408785 302209 408819 302243
rect 408819 302209 408828 302243
rect 408776 302200 408828 302209
rect 400496 302064 400548 302116
rect 451556 302107 451608 302116
rect 451556 302073 451565 302107
rect 451565 302073 451599 302107
rect 451599 302073 451608 302107
rect 451556 302064 451608 302073
rect 422484 299931 422536 299940
rect 422484 299897 422493 299931
rect 422493 299897 422527 299931
rect 422527 299897 422536 299931
rect 422484 299888 422536 299897
rect 277584 299548 277636 299600
rect 342536 299548 342588 299600
rect 230848 299480 230900 299532
rect 265164 299480 265216 299532
rect 265256 299480 265308 299532
rect 270776 299480 270828 299532
rect 309416 299480 309468 299532
rect 370136 299480 370188 299532
rect 370228 299480 370280 299532
rect 375656 299480 375708 299532
rect 375748 299480 375800 299532
rect 376944 299480 376996 299532
rect 416872 299523 416924 299532
rect 416872 299489 416881 299523
rect 416881 299489 416915 299523
rect 416915 299489 416924 299523
rect 416872 299480 416924 299489
rect 428004 299523 428056 299532
rect 428004 299489 428013 299523
rect 428013 299489 428047 299523
rect 428047 299489 428056 299523
rect 428004 299480 428056 299489
rect 433708 299480 433760 299532
rect 466552 299523 466604 299532
rect 466552 299489 466561 299523
rect 466561 299489 466595 299523
rect 466595 299489 466604 299523
rect 466552 299480 466604 299489
rect 472072 299523 472124 299532
rect 472072 299489 472081 299523
rect 472081 299489 472115 299523
rect 472115 299489 472124 299523
rect 472072 299480 472124 299489
rect 241796 299455 241848 299464
rect 241796 299421 241805 299455
rect 241805 299421 241839 299455
rect 241839 299421 241848 299455
rect 241796 299412 241848 299421
rect 277584 299412 277636 299464
rect 281816 299412 281868 299464
rect 305184 299455 305236 299464
rect 305184 299421 305193 299455
rect 305193 299421 305227 299455
rect 305227 299421 305236 299455
rect 305184 299412 305236 299421
rect 310704 299455 310756 299464
rect 310704 299421 310713 299455
rect 310713 299421 310747 299455
rect 310747 299421 310756 299455
rect 310704 299412 310756 299421
rect 331404 299412 331456 299464
rect 331496 299412 331548 299464
rect 334256 299412 334308 299464
rect 334440 299412 334492 299464
rect 346584 299455 346636 299464
rect 346584 299421 346593 299455
rect 346593 299421 346627 299455
rect 346627 299421 346636 299455
rect 346584 299412 346636 299421
rect 382464 299455 382516 299464
rect 382464 299421 382473 299455
rect 382473 299421 382507 299455
rect 382507 299421 382516 299455
rect 382464 299412 382516 299421
rect 324504 299387 324556 299396
rect 324504 299353 324513 299387
rect 324513 299353 324547 299387
rect 324547 299353 324556 299387
rect 324504 299344 324556 299353
rect 292764 298231 292816 298240
rect 292764 298197 292773 298231
rect 292773 298197 292807 298231
rect 292807 298197 292816 298231
rect 292764 298188 292816 298197
rect 232044 298120 232096 298172
rect 242992 298163 243044 298172
rect 242992 298129 243001 298163
rect 243001 298129 243035 298163
rect 243035 298129 243044 298163
rect 242992 298120 243044 298129
rect 261024 298120 261076 298172
rect 261208 298120 261260 298172
rect 356612 298120 356664 298172
rect 371240 298120 371292 298172
rect 371608 298120 371660 298172
rect 387984 298120 388036 298172
rect 408776 298163 408828 298172
rect 408776 298129 408785 298163
rect 408785 298129 408819 298163
rect 408819 298129 408828 298163
rect 408776 298120 408828 298129
rect 236276 298095 236328 298104
rect 236276 298061 236285 298095
rect 236285 298061 236319 298095
rect 236319 298061 236328 298095
rect 236276 298052 236328 298061
rect 249892 298095 249944 298104
rect 249892 298061 249901 298095
rect 249901 298061 249935 298095
rect 249935 298061 249944 298095
rect 249892 298052 249944 298061
rect 254216 298052 254268 298104
rect 254492 298052 254544 298104
rect 255504 298095 255556 298104
rect 255504 298061 255513 298095
rect 255513 298061 255547 298095
rect 255547 298061 255556 298095
rect 255504 298052 255556 298061
rect 265256 298095 265308 298104
rect 265256 298061 265265 298095
rect 265265 298061 265299 298095
rect 265299 298061 265308 298095
rect 265256 298052 265308 298061
rect 267096 298052 267148 298104
rect 270776 298052 270828 298104
rect 270868 298052 270920 298104
rect 277584 298095 277636 298104
rect 277584 298061 277593 298095
rect 277593 298061 277627 298095
rect 277627 298061 277636 298095
rect 277584 298052 277636 298061
rect 292764 298052 292816 298104
rect 295708 298095 295760 298104
rect 295708 298061 295717 298095
rect 295717 298061 295751 298095
rect 295751 298061 295760 298095
rect 295708 298052 295760 298061
rect 331404 298095 331456 298104
rect 331404 298061 331413 298095
rect 331413 298061 331447 298095
rect 331447 298061 331456 298095
rect 331404 298052 331456 298061
rect 334256 298095 334308 298104
rect 334256 298061 334265 298095
rect 334265 298061 334299 298095
rect 334299 298061 334308 298095
rect 334256 298052 334308 298061
rect 352104 298052 352156 298104
rect 353484 298095 353536 298104
rect 353484 298061 353493 298095
rect 353493 298061 353527 298095
rect 353527 298061 353536 298095
rect 353484 298052 353536 298061
rect 365904 298052 365956 298104
rect 370136 298095 370188 298104
rect 370136 298061 370145 298095
rect 370145 298061 370179 298095
rect 370179 298061 370188 298095
rect 370136 298052 370188 298061
rect 400496 298052 400548 298104
rect 400588 298052 400640 298104
rect 261024 297984 261076 298036
rect 261116 297984 261168 298036
rect 352196 297984 352248 298036
rect 365904 297916 365956 297968
rect 298376 296667 298428 296676
rect 298376 296633 298385 296667
rect 298385 296633 298419 296667
rect 298419 296633 298428 296667
rect 298376 296624 298428 296633
rect 3332 294380 3384 294432
rect 7564 294380 7616 294432
rect 295708 293267 295760 293276
rect 295708 293233 295717 293267
rect 295717 293233 295751 293267
rect 295751 293233 295760 293267
rect 295708 293224 295760 293233
rect 408776 293063 408828 293072
rect 408776 293029 408785 293063
rect 408785 293029 408819 293063
rect 408819 293029 408828 293063
rect 408776 293020 408828 293029
rect 327264 292612 327316 292664
rect 330024 292612 330076 292664
rect 332784 292612 332836 292664
rect 387984 292612 388036 292664
rect 230664 292544 230716 292596
rect 230848 292544 230900 292596
rect 451556 292612 451608 292664
rect 288624 292476 288676 292528
rect 327264 292476 327316 292528
rect 330024 292476 330076 292528
rect 332784 292476 332836 292528
rect 387984 292476 388036 292528
rect 451464 292476 451516 292528
rect 466460 292476 466512 292528
rect 466644 292476 466696 292528
rect 471980 292476 472032 292528
rect 472164 292476 472216 292528
rect 288624 292340 288676 292392
rect 357624 291864 357676 291916
rect 357808 291864 357860 291916
rect 376852 289892 376904 289944
rect 241796 289867 241848 289876
rect 241796 289833 241805 289867
rect 241805 289833 241839 289867
rect 241839 289833 241848 289867
rect 241796 289824 241848 289833
rect 281632 289867 281684 289876
rect 281632 289833 281641 289867
rect 281641 289833 281675 289867
rect 281675 289833 281684 289867
rect 281632 289824 281684 289833
rect 305184 289867 305236 289876
rect 305184 289833 305193 289867
rect 305193 289833 305227 289867
rect 305227 289833 305236 289867
rect 305184 289824 305236 289833
rect 309324 289824 309376 289876
rect 309600 289824 309652 289876
rect 310704 289867 310756 289876
rect 310704 289833 310713 289867
rect 310713 289833 310747 289867
rect 310747 289833 310756 289867
rect 310704 289824 310756 289833
rect 324504 289867 324556 289876
rect 324504 289833 324513 289867
rect 324513 289833 324547 289867
rect 324547 289833 324556 289867
rect 324504 289824 324556 289833
rect 346584 289867 346636 289876
rect 346584 289833 346593 289867
rect 346593 289833 346627 289867
rect 346627 289833 346636 289867
rect 346584 289824 346636 289833
rect 376944 289824 376996 289876
rect 381084 289824 381136 289876
rect 381360 289824 381412 289876
rect 382464 289867 382516 289876
rect 382464 289833 382473 289867
rect 382473 289833 382507 289867
rect 382507 289833 382516 289867
rect 382464 289824 382516 289833
rect 259644 289799 259696 289808
rect 259644 289765 259653 289799
rect 259653 289765 259687 289799
rect 259687 289765 259696 289799
rect 259644 289756 259696 289765
rect 287244 289799 287296 289808
rect 287244 289765 287253 289799
rect 287253 289765 287287 289799
rect 287287 289765 287296 289799
rect 287244 289756 287296 289765
rect 347964 289756 348016 289808
rect 356428 289756 356480 289808
rect 375564 289756 375616 289808
rect 375748 289756 375800 289808
rect 392124 289756 392176 289808
rect 392216 289756 392268 289808
rect 236460 289688 236512 289740
rect 309324 289731 309376 289740
rect 309324 289697 309333 289731
rect 309333 289697 309367 289731
rect 309367 289697 309376 289731
rect 309324 289688 309376 289697
rect 348056 289688 348108 289740
rect 356520 289688 356572 289740
rect 370228 289688 370280 289740
rect 249892 288439 249944 288448
rect 249892 288405 249901 288439
rect 249901 288405 249935 288439
rect 249935 288405 249944 288439
rect 249892 288396 249944 288405
rect 255504 288439 255556 288448
rect 255504 288405 255513 288439
rect 255513 288405 255547 288439
rect 255547 288405 255556 288439
rect 255504 288396 255556 288405
rect 265256 288439 265308 288448
rect 265256 288405 265265 288439
rect 265265 288405 265299 288439
rect 265299 288405 265308 288439
rect 265256 288396 265308 288405
rect 292672 288439 292724 288448
rect 292672 288405 292681 288439
rect 292681 288405 292715 288439
rect 292715 288405 292724 288439
rect 292672 288396 292724 288405
rect 331404 288439 331456 288448
rect 331404 288405 331413 288439
rect 331413 288405 331447 288439
rect 331447 288405 331456 288439
rect 331404 288396 331456 288405
rect 353576 288396 353628 288448
rect 298468 287036 298520 287088
rect 352012 287036 352064 287088
rect 352104 287036 352156 287088
rect 231952 285880 232004 285932
rect 232320 285880 232372 285932
rect 249892 285855 249944 285864
rect 249892 285821 249901 285855
rect 249901 285821 249935 285855
rect 249935 285821 249944 285855
rect 249892 285812 249944 285821
rect 230664 282956 230716 283008
rect 331404 282888 331456 282940
rect 342536 282931 342588 282940
rect 342536 282897 342545 282931
rect 342545 282897 342579 282931
rect 342579 282897 342588 282931
rect 342536 282888 342588 282897
rect 364524 282888 364576 282940
rect 381084 282888 381136 282940
rect 422300 282888 422352 282940
rect 422484 282888 422536 282940
rect 427820 282888 427872 282940
rect 428004 282888 428056 282940
rect 230664 282820 230716 282872
rect 242992 282820 243044 282872
rect 243176 282820 243228 282872
rect 259736 282752 259788 282804
rect 331496 282752 331548 282804
rect 334440 282752 334492 282804
rect 364616 282752 364668 282804
rect 381176 282752 381228 282804
rect 408776 282795 408828 282804
rect 408776 282761 408785 282795
rect 408785 282761 408819 282795
rect 408819 282761 408828 282795
rect 408776 282752 408828 282761
rect 342536 280279 342588 280288
rect 342536 280245 342545 280279
rect 342545 280245 342579 280279
rect 342579 280245 342588 280279
rect 342536 280236 342588 280245
rect 267004 280211 267056 280220
rect 267004 280177 267013 280211
rect 267013 280177 267047 280211
rect 267047 280177 267056 280211
rect 267004 280168 267056 280177
rect 277676 280168 277728 280220
rect 281724 280168 281776 280220
rect 281908 280168 281960 280220
rect 287244 280211 287296 280220
rect 287244 280177 287253 280211
rect 287253 280177 287287 280211
rect 287287 280177 287296 280211
rect 287244 280168 287296 280177
rect 292672 280168 292724 280220
rect 292764 280168 292816 280220
rect 309416 280168 309468 280220
rect 324412 280168 324464 280220
rect 324688 280168 324740 280220
rect 352012 280168 352064 280220
rect 3148 280100 3200 280152
rect 6276 280100 6328 280152
rect 230664 280100 230716 280152
rect 233332 280100 233384 280152
rect 233516 280100 233568 280152
rect 241796 280143 241848 280152
rect 241796 280109 241805 280143
rect 241805 280109 241839 280143
rect 241839 280109 241848 280143
rect 241796 280100 241848 280109
rect 242808 280100 242860 280152
rect 243176 280100 243228 280152
rect 244464 280100 244516 280152
rect 244556 280100 244608 280152
rect 265164 280100 265216 280152
rect 265256 280100 265308 280152
rect 270592 280100 270644 280152
rect 270868 280100 270920 280152
rect 283104 280143 283156 280152
rect 283104 280109 283113 280143
rect 283113 280109 283147 280143
rect 283147 280109 283156 280143
rect 283104 280100 283156 280109
rect 295432 280100 295484 280152
rect 295708 280100 295760 280152
rect 298468 280100 298520 280152
rect 305184 280143 305236 280152
rect 305184 280109 305193 280143
rect 305193 280109 305227 280143
rect 305227 280109 305236 280143
rect 305184 280100 305236 280109
rect 310704 280143 310756 280152
rect 310704 280109 310713 280143
rect 310713 280109 310747 280143
rect 310747 280109 310756 280143
rect 310704 280100 310756 280109
rect 318984 280100 319036 280152
rect 319076 280100 319128 280152
rect 327264 280143 327316 280152
rect 327264 280109 327273 280143
rect 327273 280109 327307 280143
rect 327307 280109 327316 280143
rect 327264 280100 327316 280109
rect 331128 280100 331180 280152
rect 331496 280100 331548 280152
rect 334440 280100 334492 280152
rect 346584 280143 346636 280152
rect 346584 280109 346593 280143
rect 346593 280109 346627 280143
rect 346627 280109 346636 280143
rect 346584 280100 346636 280109
rect 352104 280100 352156 280152
rect 353576 280100 353628 280152
rect 353668 280100 353720 280152
rect 356428 280100 356480 280152
rect 356520 280100 356572 280152
rect 359004 280100 359056 280152
rect 359096 280100 359148 280152
rect 364616 280100 364668 280152
rect 369952 280100 370004 280152
rect 370228 280100 370280 280152
rect 371424 280143 371476 280152
rect 371424 280109 371433 280143
rect 371433 280109 371467 280143
rect 371467 280109 371476 280143
rect 371424 280100 371476 280109
rect 375472 280100 375524 280152
rect 375748 280100 375800 280152
rect 376944 280143 376996 280152
rect 376944 280109 376953 280143
rect 376953 280109 376987 280143
rect 376987 280109 376996 280143
rect 376944 280100 376996 280109
rect 386696 280100 386748 280152
rect 386788 280100 386840 280152
rect 387984 280100 388036 280152
rect 388076 280100 388128 280152
rect 393228 280143 393280 280152
rect 393228 280109 393237 280143
rect 393237 280109 393271 280143
rect 393271 280109 393280 280143
rect 393228 280100 393280 280109
rect 400496 280143 400548 280152
rect 400496 280109 400505 280143
rect 400505 280109 400539 280143
rect 400539 280109 400548 280143
rect 400496 280100 400548 280109
rect 416872 280143 416924 280152
rect 416872 280109 416881 280143
rect 416881 280109 416915 280143
rect 416915 280109 416924 280143
rect 416872 280100 416924 280109
rect 433616 280143 433668 280152
rect 433616 280109 433625 280143
rect 433625 280109 433659 280143
rect 433659 280109 433668 280143
rect 433616 280100 433668 280109
rect 466552 280143 466604 280152
rect 466552 280109 466561 280143
rect 466561 280109 466595 280143
rect 466595 280109 466604 280143
rect 466552 280100 466604 280109
rect 472072 280143 472124 280152
rect 472072 280109 472081 280143
rect 472081 280109 472115 280143
rect 472115 280109 472124 280143
rect 472072 280100 472124 280109
rect 298284 280032 298336 280084
rect 348056 278808 348108 278860
rect 236368 278740 236420 278792
rect 236644 278740 236696 278792
rect 250076 278740 250128 278792
rect 254216 278740 254268 278792
rect 254492 278740 254544 278792
rect 347964 278740 348016 278792
rect 392124 278740 392176 278792
rect 392216 278740 392268 278792
rect 451280 278740 451332 278792
rect 451556 278740 451608 278792
rect 270592 278715 270644 278724
rect 270592 278681 270601 278715
rect 270601 278681 270635 278715
rect 270635 278681 270644 278715
rect 270592 278672 270644 278681
rect 295432 278715 295484 278724
rect 295432 278681 295441 278715
rect 295441 278681 295475 278715
rect 295475 278681 295484 278715
rect 295432 278672 295484 278681
rect 375472 278715 375524 278724
rect 375472 278681 375481 278715
rect 375481 278681 375515 278715
rect 375515 278681 375524 278715
rect 375472 278672 375524 278681
rect 408776 278715 408828 278724
rect 408776 278681 408785 278715
rect 408785 278681 408819 278715
rect 408819 278681 408828 278715
rect 408776 278672 408828 278681
rect 277676 275111 277728 275120
rect 277676 275077 277685 275111
rect 277685 275077 277719 275111
rect 277719 275077 277728 275111
rect 277676 275068 277728 275077
rect 451556 273751 451608 273760
rect 451556 273717 451565 273751
rect 451565 273717 451599 273751
rect 451599 273717 451608 273751
rect 451556 273708 451608 273717
rect 230848 273275 230900 273284
rect 230848 273241 230857 273275
rect 230857 273241 230891 273275
rect 230891 273241 230900 273275
rect 230848 273232 230900 273241
rect 254216 273300 254268 273352
rect 330024 273300 330076 273352
rect 332784 273300 332836 273352
rect 356428 273300 356480 273352
rect 357624 273300 357676 273352
rect 254124 273164 254176 273216
rect 272064 273164 272116 273216
rect 288624 273164 288676 273216
rect 294144 273164 294196 273216
rect 330024 273164 330076 273216
rect 332784 273164 332836 273216
rect 356428 273164 356480 273216
rect 357624 273164 357676 273216
rect 364524 273207 364576 273216
rect 364524 273173 364533 273207
rect 364533 273173 364567 273207
rect 364567 273173 364576 273207
rect 364524 273164 364576 273173
rect 382464 273164 382516 273216
rect 272064 273028 272116 273080
rect 288624 273028 288676 273080
rect 294144 273028 294196 273080
rect 382464 273028 382516 273080
rect 327264 272187 327316 272196
rect 327264 272153 327273 272187
rect 327273 272153 327307 272187
rect 327307 272153 327316 272187
rect 327264 272144 327316 272153
rect 334348 270623 334400 270632
rect 334348 270589 334357 270623
rect 334357 270589 334391 270623
rect 334391 270589 334400 270623
rect 334348 270580 334400 270589
rect 232044 270512 232096 270564
rect 232320 270512 232372 270564
rect 236368 270512 236420 270564
rect 241796 270555 241848 270564
rect 241796 270521 241805 270555
rect 241805 270521 241839 270555
rect 241839 270521 241848 270555
rect 241796 270512 241848 270521
rect 267004 270512 267056 270564
rect 267096 270512 267148 270564
rect 283104 270555 283156 270564
rect 283104 270521 283113 270555
rect 283113 270521 283147 270555
rect 283147 270521 283156 270555
rect 283104 270512 283156 270521
rect 305184 270555 305236 270564
rect 305184 270521 305193 270555
rect 305193 270521 305227 270555
rect 305227 270521 305236 270555
rect 305184 270512 305236 270521
rect 309324 270512 309376 270564
rect 309600 270512 309652 270564
rect 310704 270555 310756 270564
rect 310704 270521 310713 270555
rect 310713 270521 310747 270555
rect 310747 270521 310756 270555
rect 310704 270512 310756 270521
rect 346584 270555 346636 270564
rect 346584 270521 346593 270555
rect 346593 270521 346627 270555
rect 346627 270521 346636 270555
rect 346584 270512 346636 270521
rect 371424 270555 371476 270564
rect 371424 270521 371433 270555
rect 371433 270521 371467 270555
rect 371467 270521 371476 270555
rect 371424 270512 371476 270521
rect 376944 270555 376996 270564
rect 376944 270521 376953 270555
rect 376953 270521 376987 270555
rect 376987 270521 376996 270555
rect 376944 270512 376996 270521
rect 380992 270512 381044 270564
rect 381084 270512 381136 270564
rect 393228 270555 393280 270564
rect 393228 270521 393237 270555
rect 393237 270521 393271 270555
rect 393271 270521 393280 270555
rect 393228 270512 393280 270521
rect 400588 270512 400640 270564
rect 416964 270512 417016 270564
rect 433708 270512 433760 270564
rect 466644 270512 466696 270564
rect 472164 270512 472216 270564
rect 236276 270444 236328 270496
rect 252744 270487 252796 270496
rect 252744 270453 252753 270487
rect 252753 270453 252787 270487
rect 252787 270453 252796 270487
rect 252744 270444 252796 270453
rect 287244 270487 287296 270496
rect 287244 270453 287253 270487
rect 287253 270453 287287 270487
rect 287287 270453 287296 270487
rect 287244 270444 287296 270453
rect 392124 270487 392176 270496
rect 392124 270453 392133 270487
rect 392133 270453 392167 270487
rect 392167 270453 392176 270487
rect 392124 270444 392176 270453
rect 309324 270419 309376 270428
rect 309324 270385 309333 270419
rect 309333 270385 309367 270419
rect 309367 270385 309376 270419
rect 309324 270376 309376 270385
rect 381084 270419 381136 270428
rect 381084 270385 381093 270419
rect 381093 270385 381127 270419
rect 381127 270385 381136 270419
rect 381084 270376 381136 270385
rect 270776 269084 270828 269136
rect 277768 269084 277820 269136
rect 295616 269084 295668 269136
rect 259368 267724 259420 267776
rect 259552 267724 259604 267776
rect 3332 266296 3384 266348
rect 229744 266296 229796 266348
rect 530768 264868 530820 264920
rect 580172 264868 580224 264920
rect 392216 264256 392268 264308
rect 230848 263576 230900 263628
rect 231952 263576 232004 263628
rect 236276 263576 236328 263628
rect 243176 263576 243228 263628
rect 267004 263619 267056 263628
rect 267004 263585 267013 263619
rect 267013 263585 267047 263619
rect 267047 263585 267056 263619
rect 267004 263576 267056 263585
rect 324412 263619 324464 263628
rect 324412 263585 324421 263619
rect 324421 263585 324455 263619
rect 324455 263585 324464 263619
rect 324412 263576 324464 263585
rect 334348 263576 334400 263628
rect 342536 263619 342588 263628
rect 342536 263585 342545 263619
rect 342545 263585 342579 263619
rect 342579 263585 342588 263619
rect 342536 263576 342588 263585
rect 364524 263576 364576 263628
rect 422300 263576 422352 263628
rect 422484 263576 422536 263628
rect 427820 263576 427872 263628
rect 428004 263576 428056 263628
rect 236368 263508 236420 263560
rect 331312 263508 331364 263560
rect 230940 263440 230992 263492
rect 243176 263440 243228 263492
rect 331496 263440 331548 263492
rect 358912 263508 358964 263560
rect 334440 263440 334492 263492
rect 352012 263440 352064 263492
rect 352288 263440 352340 263492
rect 359096 263440 359148 263492
rect 364616 263440 364668 263492
rect 375656 263440 375708 263492
rect 397368 263440 397420 263492
rect 397736 263440 397788 263492
rect 408776 263483 408828 263492
rect 408776 263449 408785 263483
rect 408785 263449 408819 263483
rect 408819 263449 408828 263483
rect 408776 263440 408828 263449
rect 451556 263483 451608 263492
rect 451556 263449 451565 263483
rect 451565 263449 451599 263483
rect 451599 263449 451608 263483
rect 451556 263440 451608 263449
rect 252744 260899 252796 260908
rect 252744 260865 252753 260899
rect 252753 260865 252787 260899
rect 252787 260865 252796 260899
rect 252744 260856 252796 260865
rect 287244 260899 287296 260908
rect 287244 260865 287253 260899
rect 287253 260865 287287 260899
rect 287287 260865 287296 260899
rect 287244 260856 287296 260865
rect 292764 260856 292816 260908
rect 309416 260856 309468 260908
rect 324412 260899 324464 260908
rect 324412 260865 324421 260899
rect 324421 260865 324455 260899
rect 324455 260865 324464 260899
rect 324412 260856 324464 260865
rect 342536 260899 342588 260908
rect 342536 260865 342545 260899
rect 342545 260865 342579 260899
rect 342579 260865 342588 260899
rect 342536 260856 342588 260865
rect 348056 260856 348108 260908
rect 241796 260831 241848 260840
rect 241796 260797 241805 260831
rect 241805 260797 241839 260831
rect 241839 260797 241848 260831
rect 241796 260788 241848 260797
rect 242808 260788 242860 260840
rect 243176 260788 243228 260840
rect 244464 260788 244516 260840
rect 249984 260788 250036 260840
rect 254032 260788 254084 260840
rect 254216 260788 254268 260840
rect 255504 260788 255556 260840
rect 277584 260788 277636 260840
rect 277676 260788 277728 260840
rect 283104 260831 283156 260840
rect 283104 260797 283113 260831
rect 283113 260797 283147 260831
rect 283147 260797 283156 260831
rect 283104 260788 283156 260797
rect 244556 260720 244608 260772
rect 250076 260720 250128 260772
rect 295432 260788 295484 260840
rect 295616 260788 295668 260840
rect 305184 260831 305236 260840
rect 305184 260797 305193 260831
rect 305193 260797 305227 260831
rect 305227 260797 305236 260831
rect 305184 260788 305236 260797
rect 310704 260831 310756 260840
rect 310704 260797 310713 260831
rect 310713 260797 310747 260831
rect 310747 260797 310756 260831
rect 310704 260788 310756 260797
rect 318984 260788 319036 260840
rect 319076 260788 319128 260840
rect 327264 260831 327316 260840
rect 327264 260797 327273 260831
rect 327273 260797 327307 260831
rect 327307 260797 327316 260831
rect 327264 260788 327316 260797
rect 331128 260788 331180 260840
rect 331496 260788 331548 260840
rect 334440 260788 334492 260840
rect 346584 260831 346636 260840
rect 346584 260797 346593 260831
rect 346593 260797 346627 260831
rect 346627 260797 346636 260831
rect 346584 260788 346636 260797
rect 348148 260788 348200 260840
rect 356520 260856 356572 260908
rect 381176 260856 381228 260908
rect 359096 260788 359148 260840
rect 364248 260788 364300 260840
rect 364616 260788 364668 260840
rect 371424 260831 371476 260840
rect 371424 260797 371433 260831
rect 371433 260797 371467 260831
rect 371467 260797 371476 260831
rect 371424 260788 371476 260797
rect 375656 260788 375708 260840
rect 376944 260831 376996 260840
rect 376944 260797 376953 260831
rect 376953 260797 376987 260831
rect 376987 260797 376996 260831
rect 376944 260788 376996 260797
rect 400496 260831 400548 260840
rect 400496 260797 400505 260831
rect 400505 260797 400539 260831
rect 400539 260797 400548 260831
rect 400496 260788 400548 260797
rect 416872 260831 416924 260840
rect 416872 260797 416881 260831
rect 416881 260797 416915 260831
rect 416915 260797 416924 260831
rect 416872 260788 416924 260797
rect 433616 260831 433668 260840
rect 433616 260797 433625 260831
rect 433625 260797 433659 260831
rect 433659 260797 433668 260831
rect 433616 260788 433668 260797
rect 466552 260831 466604 260840
rect 466552 260797 466561 260831
rect 466561 260797 466595 260831
rect 466595 260797 466604 260831
rect 466552 260788 466604 260797
rect 472072 260831 472124 260840
rect 472072 260797 472081 260831
rect 472081 260797 472115 260831
rect 472115 260797 472124 260831
rect 472072 260788 472124 260797
rect 255596 260720 255648 260772
rect 292764 260720 292816 260772
rect 309416 260720 309468 260772
rect 342536 260720 342588 260772
rect 356428 260720 356480 260772
rect 397368 260720 397420 260772
rect 397736 260720 397788 260772
rect 231860 259471 231912 259480
rect 231860 259437 231869 259471
rect 231869 259437 231903 259471
rect 231903 259437 231912 259471
rect 231860 259428 231912 259437
rect 267004 259471 267056 259480
rect 267004 259437 267013 259471
rect 267013 259437 267047 259471
rect 267047 259437 267056 259471
rect 267004 259428 267056 259437
rect 282000 259360 282052 259412
rect 295432 259403 295484 259412
rect 295432 259369 295441 259403
rect 295441 259369 295475 259403
rect 295475 259369 295484 259403
rect 295432 259360 295484 259369
rect 451556 259403 451608 259412
rect 451556 259369 451565 259403
rect 451565 259369 451599 259403
rect 451599 259369 451608 259403
rect 451556 259360 451608 259369
rect 292856 258000 292908 258052
rect 231860 254600 231912 254652
rect 232044 254600 232096 254652
rect 348148 254600 348200 254652
rect 353668 254600 353720 254652
rect 230940 254439 230992 254448
rect 230940 254405 230949 254439
rect 230949 254405 230983 254439
rect 230983 254405 230992 254439
rect 230940 254396 230992 254405
rect 330024 253988 330076 254040
rect 356428 254031 356480 254040
rect 356428 253997 356437 254031
rect 356437 253997 356471 254031
rect 356471 253997 356480 254031
rect 356428 253988 356480 253997
rect 357624 253988 357676 254040
rect 236368 253852 236420 253904
rect 272064 253852 272116 253904
rect 288624 253852 288676 253904
rect 294144 253852 294196 253904
rect 330024 253852 330076 253904
rect 357624 253852 357676 253904
rect 382464 253852 382516 253904
rect 236276 253716 236328 253768
rect 272064 253716 272116 253768
rect 288624 253716 288676 253768
rect 294144 253716 294196 253768
rect 382464 253716 382516 253768
rect 530676 252492 530728 252544
rect 579620 252492 579672 252544
rect 334348 251311 334400 251320
rect 334348 251277 334357 251311
rect 334357 251277 334391 251311
rect 334391 251277 334400 251311
rect 334348 251268 334400 251277
rect 359004 251311 359056 251320
rect 359004 251277 359013 251311
rect 359013 251277 359047 251311
rect 359047 251277 359056 251311
rect 359004 251268 359056 251277
rect 241796 251243 241848 251252
rect 241796 251209 241805 251243
rect 241805 251209 241839 251243
rect 241839 251209 241848 251243
rect 241796 251200 241848 251209
rect 283104 251243 283156 251252
rect 283104 251209 283113 251243
rect 283113 251209 283147 251243
rect 283147 251209 283156 251243
rect 283104 251200 283156 251209
rect 305184 251243 305236 251252
rect 305184 251209 305193 251243
rect 305193 251209 305227 251243
rect 305227 251209 305236 251243
rect 305184 251200 305236 251209
rect 309324 251243 309376 251252
rect 309324 251209 309333 251243
rect 309333 251209 309367 251243
rect 309367 251209 309376 251243
rect 309324 251200 309376 251209
rect 310704 251243 310756 251252
rect 310704 251209 310713 251243
rect 310713 251209 310747 251243
rect 310747 251209 310756 251243
rect 310704 251200 310756 251209
rect 327264 251243 327316 251252
rect 327264 251209 327273 251243
rect 327273 251209 327307 251243
rect 327307 251209 327316 251243
rect 327264 251200 327316 251209
rect 342444 251243 342496 251252
rect 342444 251209 342453 251243
rect 342453 251209 342487 251243
rect 342487 251209 342496 251243
rect 342444 251200 342496 251209
rect 346584 251243 346636 251252
rect 346584 251209 346593 251243
rect 346593 251209 346627 251243
rect 346627 251209 346636 251243
rect 346584 251200 346636 251209
rect 371424 251243 371476 251252
rect 371424 251209 371433 251243
rect 371433 251209 371467 251243
rect 371467 251209 371476 251243
rect 371424 251200 371476 251209
rect 375564 251243 375616 251252
rect 375564 251209 375573 251243
rect 375573 251209 375607 251243
rect 375607 251209 375616 251243
rect 375564 251200 375616 251209
rect 376944 251243 376996 251252
rect 376944 251209 376953 251243
rect 376953 251209 376987 251243
rect 376987 251209 376996 251243
rect 376944 251200 376996 251209
rect 381084 251200 381136 251252
rect 381360 251200 381412 251252
rect 400588 251200 400640 251252
rect 416964 251200 417016 251252
rect 433708 251200 433760 251252
rect 466644 251200 466696 251252
rect 472164 251200 472216 251252
rect 252744 251175 252796 251184
rect 252744 251141 252753 251175
rect 252753 251141 252787 251175
rect 252787 251141 252796 251175
rect 252744 251132 252796 251141
rect 270592 251132 270644 251184
rect 270960 251132 271012 251184
rect 287244 251175 287296 251184
rect 287244 251141 287253 251175
rect 287253 251141 287287 251175
rect 287287 251141 287296 251175
rect 287244 251132 287296 251141
rect 298284 251132 298336 251184
rect 334348 251175 334400 251184
rect 334348 251141 334357 251175
rect 334357 251141 334391 251175
rect 334391 251141 334400 251175
rect 334348 251132 334400 251141
rect 359004 251175 359056 251184
rect 359004 251141 359013 251175
rect 359013 251141 359047 251175
rect 359047 251141 359056 251175
rect 359004 251132 359056 251141
rect 370044 251132 370096 251184
rect 254032 251064 254084 251116
rect 254216 251064 254268 251116
rect 356428 251107 356480 251116
rect 356428 251073 356437 251107
rect 356437 251073 356471 251107
rect 356471 251073 356480 251107
rect 356428 251064 356480 251073
rect 381084 251107 381136 251116
rect 381084 251073 381093 251107
rect 381093 251073 381127 251107
rect 381127 251073 381136 251107
rect 381084 251064 381136 251073
rect 386604 249840 386656 249892
rect 386696 249840 386748 249892
rect 392124 249840 392176 249892
rect 392216 249840 392268 249892
rect 259552 249772 259604 249824
rect 259736 249772 259788 249824
rect 292856 249704 292908 249756
rect 324228 245420 324280 245472
rect 324412 245420 324464 245472
rect 232044 244332 232096 244384
rect 233332 244264 233384 244316
rect 233516 244264 233568 244316
rect 236276 244307 236328 244316
rect 236276 244273 236285 244307
rect 236285 244273 236319 244307
rect 236319 244273 236328 244307
rect 236276 244264 236328 244273
rect 356428 244264 356480 244316
rect 231952 244196 232004 244248
rect 230940 244171 230992 244180
rect 230940 244137 230949 244171
rect 230949 244137 230983 244171
rect 230983 244137 230992 244171
rect 230940 244128 230992 244137
rect 334348 244171 334400 244180
rect 334348 244137 334357 244171
rect 334357 244137 334391 244171
rect 334391 244137 334400 244171
rect 334348 244128 334400 244137
rect 386696 244264 386748 244316
rect 422300 244264 422352 244316
rect 422484 244264 422536 244316
rect 427820 244264 427872 244316
rect 428004 244264 428056 244316
rect 386604 244196 386656 244248
rect 356520 244128 356572 244180
rect 359004 244171 359056 244180
rect 359004 244137 359013 244171
rect 359013 244137 359047 244171
rect 359047 244137 359056 244171
rect 359004 244128 359056 244137
rect 408776 244128 408828 244180
rect 408960 244128 409012 244180
rect 451556 244171 451608 244180
rect 451556 244137 451565 244171
rect 451565 244137 451599 244171
rect 451599 244137 451608 244171
rect 451556 244128 451608 244137
rect 298192 242675 298244 242684
rect 298192 242641 298201 242675
rect 298201 242641 298235 242675
rect 298235 242641 298244 242675
rect 298192 242632 298244 242641
rect 364248 242156 364300 242208
rect 364616 242156 364668 242208
rect 281908 241587 281960 241596
rect 281908 241553 281917 241587
rect 281917 241553 281951 241587
rect 281951 241553 281960 241587
rect 281908 241544 281960 241553
rect 242992 241476 243044 241528
rect 243176 241476 243228 241528
rect 252744 241519 252796 241528
rect 252744 241485 252753 241519
rect 252753 241485 252787 241519
rect 252787 241485 252796 241519
rect 252744 241476 252796 241485
rect 254032 241476 254084 241528
rect 254216 241476 254268 241528
rect 259552 241476 259604 241528
rect 259736 241476 259788 241528
rect 287244 241519 287296 241528
rect 287244 241485 287253 241519
rect 287253 241485 287287 241519
rect 287287 241485 287296 241519
rect 287244 241476 287296 241485
rect 309508 241476 309560 241528
rect 309600 241476 309652 241528
rect 331128 241476 331180 241528
rect 331496 241476 331548 241528
rect 348056 241519 348108 241528
rect 348056 241485 348065 241519
rect 348065 241485 348099 241519
rect 348099 241485 348108 241519
rect 348056 241476 348108 241485
rect 353576 241519 353628 241528
rect 353576 241485 353585 241519
rect 353585 241485 353619 241519
rect 353619 241485 353628 241519
rect 353576 241476 353628 241485
rect 369952 241519 370004 241528
rect 369952 241485 369961 241519
rect 369961 241485 369995 241519
rect 369995 241485 370004 241519
rect 369952 241476 370004 241485
rect 375748 241476 375800 241528
rect 375840 241476 375892 241528
rect 381176 241476 381228 241528
rect 281908 241451 281960 241460
rect 281908 241417 281917 241451
rect 281917 241417 281951 241451
rect 281951 241417 281960 241451
rect 281908 241408 281960 241417
rect 466552 241408 466604 241460
rect 466644 241408 466696 241460
rect 236276 240227 236328 240236
rect 236276 240193 236285 240227
rect 236285 240193 236319 240227
rect 236319 240193 236328 240227
rect 236276 240184 236328 240193
rect 292764 240116 292816 240168
rect 292856 240116 292908 240168
rect 392216 240116 392268 240168
rect 392400 240116 392452 240168
rect 231952 240048 232004 240100
rect 232228 240048 232280 240100
rect 236276 240091 236328 240100
rect 236276 240057 236285 240091
rect 236285 240057 236319 240091
rect 236319 240057 236328 240091
rect 236276 240048 236328 240057
rect 295524 240048 295576 240100
rect 298192 240048 298244 240100
rect 298284 240048 298336 240100
rect 298284 238688 298336 238740
rect 298560 238688 298612 238740
rect 348056 238731 348108 238740
rect 348056 238697 348065 238731
rect 348065 238697 348099 238731
rect 348099 238697 348108 238731
rect 348056 238688 348108 238697
rect 295524 237371 295576 237380
rect 295524 237337 295533 237371
rect 295533 237337 295567 237371
rect 295567 237337 295576 237371
rect 295524 237328 295576 237337
rect 2780 237260 2832 237312
rect 4988 237260 5040 237312
rect 392216 236716 392268 236768
rect 324228 236648 324280 236700
rect 324412 236648 324464 236700
rect 364616 235900 364668 235952
rect 230940 234676 230992 234728
rect 353576 234676 353628 234728
rect 356520 234676 356572 234728
rect 381084 234719 381136 234728
rect 381084 234685 381093 234719
rect 381093 234685 381127 234719
rect 381127 234685 381136 234719
rect 381084 234676 381136 234685
rect 261116 234608 261168 234660
rect 327356 234608 327408 234660
rect 330116 234608 330168 234660
rect 352012 234651 352064 234660
rect 352012 234617 352021 234651
rect 352021 234617 352055 234651
rect 352055 234617 352064 234651
rect 352012 234608 352064 234617
rect 357716 234608 357768 234660
rect 408776 234676 408828 234728
rect 451556 234676 451608 234728
rect 230848 234540 230900 234592
rect 261024 234540 261076 234592
rect 272064 234540 272116 234592
rect 281908 234583 281960 234592
rect 281908 234549 281917 234583
rect 281917 234549 281951 234583
rect 281951 234549 281960 234583
rect 281908 234540 281960 234549
rect 288624 234540 288676 234592
rect 294144 234540 294196 234592
rect 327264 234540 327316 234592
rect 330024 234540 330076 234592
rect 353576 234540 353628 234592
rect 357624 234540 357676 234592
rect 371424 234540 371476 234592
rect 382464 234540 382516 234592
rect 408684 234540 408736 234592
rect 451464 234540 451516 234592
rect 272064 234404 272116 234456
rect 288624 234404 288676 234456
rect 294144 234404 294196 234456
rect 371424 234404 371476 234456
rect 382464 234404 382516 234456
rect 334348 231956 334400 232008
rect 359004 231956 359056 232008
rect 242992 231820 243044 231872
rect 243084 231820 243136 231872
rect 277584 231820 277636 231872
rect 277676 231820 277728 231872
rect 282920 231820 282972 231872
rect 283104 231820 283156 231872
rect 305184 231820 305236 231872
rect 305368 231820 305420 231872
rect 310704 231820 310756 231872
rect 310888 231820 310940 231872
rect 318984 231820 319036 231872
rect 319076 231820 319128 231872
rect 331496 231820 331548 231872
rect 334440 231820 334492 231872
rect 346584 231820 346636 231872
rect 346768 231820 346820 231872
rect 359096 231820 359148 231872
rect 369952 231820 370004 231872
rect 370044 231820 370096 231872
rect 375564 231820 375616 231872
rect 375840 231820 375892 231872
rect 376760 231820 376812 231872
rect 376944 231820 376996 231872
rect 381176 231820 381228 231872
rect 393136 231820 393188 231872
rect 393228 231820 393280 231872
rect 397736 231820 397788 231872
rect 397920 231820 397972 231872
rect 400312 231820 400364 231872
rect 400588 231820 400640 231872
rect 416964 231820 417016 231872
rect 417148 231820 417200 231872
rect 433432 231820 433484 231872
rect 433708 231820 433760 231872
rect 472164 231820 472216 231872
rect 472348 231820 472400 231872
rect 259644 231795 259696 231804
rect 259644 231761 259653 231795
rect 259653 231761 259687 231795
rect 259687 231761 259696 231795
rect 259644 231752 259696 231761
rect 408684 231795 408736 231804
rect 408684 231761 408693 231795
rect 408693 231761 408727 231795
rect 408727 231761 408736 231795
rect 408684 231752 408736 231761
rect 243176 231727 243228 231736
rect 243176 231693 243185 231727
rect 243185 231693 243219 231727
rect 243219 231693 243228 231727
rect 243176 231684 243228 231693
rect 331496 231684 331548 231736
rect 236276 230571 236328 230580
rect 236276 230537 236285 230571
rect 236285 230537 236319 230571
rect 236319 230537 236328 230571
rect 236276 230528 236328 230537
rect 265164 230528 265216 230580
rect 265256 230528 265308 230580
rect 292764 230528 292816 230580
rect 292856 230528 292908 230580
rect 348056 230367 348108 230376
rect 348056 230333 348065 230367
rect 348065 230333 348099 230367
rect 348099 230333 348108 230367
rect 348056 230324 348108 230333
rect 352196 230324 352248 230376
rect 356428 229211 356480 229220
rect 356428 229177 356437 229211
rect 356437 229177 356471 229211
rect 356471 229177 356480 229211
rect 356428 229168 356480 229177
rect 356428 229075 356480 229084
rect 356428 229041 356437 229075
rect 356437 229041 356471 229075
rect 356471 229041 356480 229075
rect 356428 229032 356480 229041
rect 295524 227783 295576 227792
rect 295524 227749 295533 227783
rect 295533 227749 295567 227783
rect 295567 227749 295576 227783
rect 295524 227740 295576 227749
rect 233332 224952 233384 225004
rect 233516 224952 233568 225004
rect 254124 224952 254176 225004
rect 267096 224995 267148 225004
rect 267096 224961 267105 224995
rect 267105 224961 267139 224995
rect 267139 224961 267148 224995
rect 267096 224952 267148 224961
rect 295524 224952 295576 225004
rect 309324 224952 309376 225004
rect 324412 224995 324464 225004
rect 324412 224961 324421 224995
rect 324421 224961 324455 224995
rect 324455 224961 324464 224995
rect 324412 224952 324464 224961
rect 381176 224995 381228 225004
rect 381176 224961 381185 224995
rect 381185 224961 381219 224995
rect 381219 224961 381228 224995
rect 381176 224952 381228 224961
rect 386604 224952 386656 225004
rect 397736 224952 397788 225004
rect 422300 224952 422352 225004
rect 422484 224952 422536 225004
rect 427820 224952 427872 225004
rect 428004 224952 428056 225004
rect 254216 224816 254268 224868
rect 265164 224816 265216 224868
rect 265348 224816 265400 224868
rect 295616 224816 295668 224868
rect 356428 224927 356480 224936
rect 356428 224893 356437 224927
rect 356437 224893 356471 224927
rect 356471 224893 356480 224927
rect 356428 224884 356480 224893
rect 309416 224816 309468 224868
rect 386696 224816 386748 224868
rect 397736 224816 397788 224868
rect 243360 224204 243412 224256
rect 231952 222232 232004 222284
rect 232228 222232 232280 222284
rect 324412 222275 324464 222284
rect 324412 222241 324421 222275
rect 324421 222241 324455 222275
rect 324455 222241 324464 222275
rect 324412 222232 324464 222241
rect 230664 222164 230716 222216
rect 230940 222164 230992 222216
rect 252744 222164 252796 222216
rect 252928 222164 252980 222216
rect 259736 222164 259788 222216
rect 281908 222207 281960 222216
rect 281908 222173 281917 222207
rect 281917 222173 281951 222207
rect 281951 222173 281960 222207
rect 281908 222164 281960 222173
rect 287244 222164 287296 222216
rect 287428 222164 287480 222216
rect 381176 222207 381228 222216
rect 381176 222173 381185 222207
rect 381185 222173 381219 222207
rect 381219 222173 381228 222207
rect 381176 222164 381228 222173
rect 392216 222164 392268 222216
rect 393228 222164 393280 222216
rect 393412 222164 393464 222216
rect 408776 222164 408828 222216
rect 451280 222164 451332 222216
rect 451556 222164 451608 222216
rect 324412 222139 324464 222148
rect 324412 222105 324421 222139
rect 324421 222105 324455 222139
rect 324455 222105 324464 222139
rect 324412 222096 324464 222105
rect 466552 222096 466604 222148
rect 466644 222096 466696 222148
rect 236276 220804 236328 220856
rect 236460 220804 236512 220856
rect 267096 220847 267148 220856
rect 267096 220813 267105 220847
rect 267105 220813 267139 220847
rect 267139 220813 267148 220847
rect 267096 220804 267148 220813
rect 281908 220847 281960 220856
rect 281908 220813 281917 220847
rect 281917 220813 281951 220847
rect 281951 220813 281960 220847
rect 281908 220804 281960 220813
rect 298376 220804 298428 220856
rect 298560 220804 298612 220856
rect 331312 220804 331364 220856
rect 331588 220804 331640 220856
rect 352012 220804 352064 220856
rect 352196 220804 352248 220856
rect 324412 219555 324464 219564
rect 324412 219521 324421 219555
rect 324421 219521 324455 219555
rect 324455 219521 324464 219555
rect 324412 219512 324464 219521
rect 243084 219376 243136 219428
rect 243360 219376 243412 219428
rect 267096 219376 267148 219428
rect 331128 219376 331180 219428
rect 331312 219376 331364 219428
rect 364432 218059 364484 218068
rect 364432 218025 364441 218059
rect 364441 218025 364475 218059
rect 364475 218025 364484 218059
rect 364432 218016 364484 218025
rect 243084 217991 243136 218000
rect 243084 217957 243093 217991
rect 243093 217957 243127 217991
rect 243127 217957 243136 217991
rect 243084 217948 243136 217957
rect 577504 217948 577556 218000
rect 579620 217948 579672 218000
rect 254216 217404 254268 217456
rect 259736 217404 259788 217456
rect 254124 217336 254176 217388
rect 259644 217336 259696 217388
rect 236368 215976 236420 216028
rect 236552 215976 236604 216028
rect 298376 215432 298428 215484
rect 230940 215364 230992 215416
rect 281908 215364 281960 215416
rect 295616 215364 295668 215416
rect 370044 215364 370096 215416
rect 381084 215407 381136 215416
rect 381084 215373 381093 215407
rect 381093 215373 381127 215407
rect 381127 215373 381136 215407
rect 381084 215364 381136 215373
rect 309324 215339 309376 215348
rect 309324 215305 309333 215339
rect 309333 215305 309367 215339
rect 309367 215305 309376 215339
rect 309324 215296 309376 215305
rect 327356 215296 327408 215348
rect 330116 215296 330168 215348
rect 357716 215296 357768 215348
rect 397644 215339 397696 215348
rect 397644 215305 397653 215339
rect 397653 215305 397687 215339
rect 397687 215305 397696 215339
rect 397644 215296 397696 215305
rect 408776 215364 408828 215416
rect 451556 215364 451608 215416
rect 230848 215228 230900 215280
rect 231768 215228 231820 215280
rect 231952 215228 232004 215280
rect 233332 215228 233384 215280
rect 233516 215228 233568 215280
rect 272064 215228 272116 215280
rect 281908 215228 281960 215280
rect 327264 215228 327316 215280
rect 330024 215228 330076 215280
rect 357624 215228 357676 215280
rect 370044 215228 370096 215280
rect 371424 215228 371476 215280
rect 382464 215228 382516 215280
rect 408684 215228 408736 215280
rect 451464 215228 451516 215280
rect 272064 215092 272116 215144
rect 371424 215092 371476 215144
rect 382464 215092 382516 215144
rect 334348 212644 334400 212696
rect 356520 212576 356572 212628
rect 359004 212576 359056 212628
rect 252744 212508 252796 212560
rect 252836 212508 252888 212560
rect 270776 212508 270828 212560
rect 270960 212508 271012 212560
rect 277584 212508 277636 212560
rect 277676 212508 277728 212560
rect 305184 212508 305236 212560
rect 305368 212508 305420 212560
rect 309416 212508 309468 212560
rect 310704 212508 310756 212560
rect 310888 212508 310940 212560
rect 318984 212508 319036 212560
rect 319076 212508 319128 212560
rect 334440 212508 334492 212560
rect 346584 212508 346636 212560
rect 346768 212508 346820 212560
rect 347964 212508 348016 212560
rect 348148 212508 348200 212560
rect 352012 212508 352064 212560
rect 352104 212508 352156 212560
rect 353484 212508 353536 212560
rect 353668 212508 353720 212560
rect 356428 212508 356480 212560
rect 375564 212508 375616 212560
rect 375840 212508 375892 212560
rect 376760 212508 376812 212560
rect 376944 212508 376996 212560
rect 381176 212508 381228 212560
rect 393136 212508 393188 212560
rect 393228 212508 393280 212560
rect 397552 212508 397604 212560
rect 400312 212508 400364 212560
rect 400588 212508 400640 212560
rect 416964 212508 417016 212560
rect 417148 212508 417200 212560
rect 433432 212508 433484 212560
rect 433708 212508 433760 212560
rect 472164 212508 472216 212560
rect 472348 212508 472400 212560
rect 408684 212483 408736 212492
rect 408684 212449 408693 212483
rect 408693 212449 408727 212483
rect 408727 212449 408736 212483
rect 408684 212440 408736 212449
rect 298284 211259 298336 211268
rect 298284 211225 298293 211259
rect 298293 211225 298327 211259
rect 298327 211225 298336 211259
rect 298284 211216 298336 211225
rect 281724 211123 281776 211132
rect 281724 211089 281733 211123
rect 281733 211089 281767 211123
rect 281767 211089 281776 211123
rect 281724 211080 281776 211089
rect 295432 211123 295484 211132
rect 295432 211089 295441 211123
rect 295441 211089 295475 211123
rect 295475 211089 295484 211123
rect 295432 211080 295484 211089
rect 298284 211123 298336 211132
rect 298284 211089 298293 211123
rect 298293 211089 298327 211123
rect 298327 211089 298336 211123
rect 298284 211080 298336 211089
rect 356428 211123 356480 211132
rect 356428 211089 356437 211123
rect 356437 211089 356471 211123
rect 356471 211089 356480 211123
rect 356428 211080 356480 211089
rect 370044 211080 370096 211132
rect 370228 211080 370280 211132
rect 267004 209831 267056 209840
rect 267004 209797 267013 209831
rect 267013 209797 267047 209831
rect 267047 209797 267056 209831
rect 267004 209788 267056 209797
rect 265164 209763 265216 209772
rect 265164 209729 265173 209763
rect 265173 209729 265207 209763
rect 265207 209729 265216 209763
rect 265164 209720 265216 209729
rect 358912 208403 358964 208412
rect 358912 208369 358921 208403
rect 358921 208369 358955 208403
rect 358955 208369 358964 208403
rect 358912 208360 358964 208369
rect 295432 206252 295484 206304
rect 295708 206252 295760 206304
rect 259644 205640 259696 205692
rect 309416 205683 309468 205692
rect 309416 205649 309425 205683
rect 309425 205649 309459 205683
rect 309459 205649 309468 205683
rect 309416 205640 309468 205649
rect 324412 205683 324464 205692
rect 324412 205649 324421 205683
rect 324421 205649 324455 205683
rect 324455 205649 324464 205683
rect 324412 205640 324464 205649
rect 347964 205640 348016 205692
rect 353484 205640 353536 205692
rect 381176 205640 381228 205692
rect 422300 205640 422352 205692
rect 422484 205640 422536 205692
rect 427820 205640 427872 205692
rect 428004 205640 428056 205692
rect 236276 205615 236328 205624
rect 236276 205581 236285 205615
rect 236285 205581 236319 205615
rect 236319 205581 236328 205615
rect 236276 205572 236328 205581
rect 298284 205615 298336 205624
rect 298284 205581 298293 205615
rect 298293 205581 298327 205615
rect 298327 205581 298336 205615
rect 298284 205572 298336 205581
rect 259736 205504 259788 205556
rect 353576 205572 353628 205624
rect 530584 205572 530636 205624
rect 580172 205572 580224 205624
rect 348056 205504 348108 205556
rect 381176 205504 381228 205556
rect 233516 205164 233568 205216
rect 233516 205028 233568 205080
rect 331496 202920 331548 202972
rect 230664 202852 230716 202904
rect 230940 202852 230992 202904
rect 231952 202852 232004 202904
rect 232044 202852 232096 202904
rect 236276 202895 236328 202904
rect 236276 202861 236285 202895
rect 236285 202861 236319 202895
rect 236319 202861 236328 202895
rect 236276 202852 236328 202861
rect 252468 202852 252520 202904
rect 252560 202852 252612 202904
rect 309416 202895 309468 202904
rect 309416 202861 309425 202895
rect 309425 202861 309459 202895
rect 309459 202861 309468 202895
rect 309416 202852 309468 202861
rect 324412 202895 324464 202904
rect 324412 202861 324421 202895
rect 324421 202861 324455 202895
rect 324455 202861 324464 202895
rect 324412 202852 324464 202861
rect 342628 202852 342680 202904
rect 342720 202852 342772 202904
rect 352012 202852 352064 202904
rect 352104 202852 352156 202904
rect 393228 202852 393280 202904
rect 393412 202852 393464 202904
rect 397368 202852 397420 202904
rect 397736 202852 397788 202904
rect 408776 202852 408828 202904
rect 451280 202852 451332 202904
rect 451556 202852 451608 202904
rect 265256 202784 265308 202836
rect 281816 202784 281868 202836
rect 356428 202827 356480 202836
rect 356428 202793 356437 202827
rect 356437 202793 356471 202827
rect 356471 202793 356480 202827
rect 356428 202784 356480 202793
rect 466552 202784 466604 202836
rect 466644 202784 466696 202836
rect 331404 201535 331456 201544
rect 331404 201501 331413 201535
rect 331413 201501 331447 201535
rect 331447 201501 331456 201535
rect 331404 201492 331456 201501
rect 243084 201467 243136 201476
rect 243084 201433 243093 201467
rect 243093 201433 243127 201467
rect 243127 201433 243136 201467
rect 243084 201424 243136 201433
rect 375564 201424 375616 201476
rect 375840 201424 375892 201476
rect 381084 201424 381136 201476
rect 381360 201424 381412 201476
rect 292764 200064 292816 200116
rect 292856 200064 292908 200116
rect 295432 200064 295484 200116
rect 295708 200064 295760 200116
rect 236276 198679 236328 198688
rect 236276 198645 236285 198679
rect 236285 198645 236319 198679
rect 236319 198645 236328 198679
rect 236276 198636 236328 198645
rect 292856 198636 292908 198688
rect 331036 196596 331088 196648
rect 331404 196596 331456 196648
rect 342720 196596 342772 196648
rect 342904 196596 342956 196648
rect 230940 196052 230992 196104
rect 243176 196052 243228 196104
rect 270776 196095 270828 196104
rect 270776 196061 270785 196095
rect 270785 196061 270819 196095
rect 270819 196061 270828 196095
rect 270776 196052 270828 196061
rect 261116 195984 261168 196036
rect 281908 196052 281960 196104
rect 324412 196095 324464 196104
rect 324412 196061 324421 196095
rect 324421 196061 324455 196095
rect 324455 196061 324464 196095
rect 324412 196052 324464 196061
rect 364616 196052 364668 196104
rect 370044 196052 370096 196104
rect 309324 196027 309376 196036
rect 309324 195993 309333 196027
rect 309333 195993 309367 196027
rect 309367 195993 309376 196027
rect 309324 195984 309376 195993
rect 330116 195984 330168 196036
rect 358912 195984 358964 196036
rect 359096 195984 359148 196036
rect 397644 196027 397696 196036
rect 397644 195993 397653 196027
rect 397653 195993 397687 196027
rect 397687 195993 397696 196027
rect 397644 195984 397696 195993
rect 408776 196052 408828 196104
rect 451556 196052 451608 196104
rect 230848 195916 230900 195968
rect 243176 195916 243228 195968
rect 261024 195916 261076 195968
rect 277492 195916 277544 195968
rect 277676 195916 277728 195968
rect 281816 195916 281868 195968
rect 318892 195916 318944 195968
rect 319076 195916 319128 195968
rect 330024 195916 330076 195968
rect 364616 195916 364668 195968
rect 370044 195916 370096 195968
rect 371424 195916 371476 195968
rect 382464 195916 382516 195968
rect 408684 195916 408736 195968
rect 451464 195916 451516 195968
rect 371424 195780 371476 195832
rect 382464 195780 382516 195832
rect 392032 195236 392084 195288
rect 392308 195236 392360 195288
rect 3148 194284 3200 194336
rect 6184 194284 6236 194336
rect 334348 193332 334400 193384
rect 265164 193264 265216 193316
rect 265348 193264 265400 193316
rect 327356 193264 327408 193316
rect 331220 193264 331272 193316
rect 252560 193196 252612 193248
rect 252744 193196 252796 193248
rect 254124 193196 254176 193248
rect 254308 193196 254360 193248
rect 259736 193196 259788 193248
rect 266360 193196 266412 193248
rect 266544 193196 266596 193248
rect 267004 193196 267056 193248
rect 267096 193196 267148 193248
rect 294144 193196 294196 193248
rect 298376 193196 298428 193248
rect 305184 193196 305236 193248
rect 305368 193196 305420 193248
rect 309416 193196 309468 193248
rect 310704 193196 310756 193248
rect 310888 193196 310940 193248
rect 259644 193128 259696 193180
rect 270776 193171 270828 193180
rect 270776 193137 270785 193171
rect 270785 193137 270819 193171
rect 270819 193137 270828 193171
rect 270776 193128 270828 193137
rect 356520 193264 356572 193316
rect 386604 193264 386656 193316
rect 386788 193264 386840 193316
rect 334440 193196 334492 193248
rect 346584 193196 346636 193248
rect 346768 193196 346820 193248
rect 347964 193196 348016 193248
rect 348148 193196 348200 193248
rect 353484 193196 353536 193248
rect 353668 193196 353720 193248
rect 356428 193196 356480 193248
rect 376760 193196 376812 193248
rect 376944 193196 376996 193248
rect 393136 193196 393188 193248
rect 393228 193196 393280 193248
rect 397552 193196 397604 193248
rect 400312 193196 400364 193248
rect 400588 193196 400640 193248
rect 416964 193196 417016 193248
rect 417148 193196 417200 193248
rect 433432 193196 433484 193248
rect 433708 193196 433760 193248
rect 472164 193196 472216 193248
rect 472348 193196 472400 193248
rect 294236 193128 294288 193180
rect 327356 193128 327408 193180
rect 331220 193128 331272 193180
rect 298284 191879 298336 191888
rect 298284 191845 298293 191879
rect 298293 191845 298327 191879
rect 298327 191845 298336 191879
rect 298284 191836 298336 191845
rect 324412 191879 324464 191888
rect 324412 191845 324421 191879
rect 324421 191845 324455 191879
rect 324455 191845 324464 191879
rect 324412 191836 324464 191845
rect 266544 191768 266596 191820
rect 270408 191768 270460 191820
rect 270776 191768 270828 191820
rect 369768 191768 369820 191820
rect 370044 191768 370096 191820
rect 375472 191768 375524 191820
rect 375564 191768 375616 191820
rect 324228 191700 324280 191752
rect 324412 191700 324464 191752
rect 236368 189048 236420 189100
rect 295616 188479 295668 188488
rect 295616 188445 295625 188479
rect 295625 188445 295659 188479
rect 295659 188445 295668 188479
rect 295616 188436 295668 188445
rect 327172 188096 327224 188148
rect 327356 188096 327408 188148
rect 244464 186940 244516 186992
rect 244648 186940 244700 186992
rect 298284 186464 298336 186516
rect 233332 186328 233384 186380
rect 233516 186328 233568 186380
rect 267096 186396 267148 186448
rect 334440 186439 334492 186448
rect 334440 186405 334449 186439
rect 334449 186405 334483 186439
rect 334483 186405 334492 186439
rect 334440 186396 334492 186405
rect 321744 186328 321796 186380
rect 352104 186396 352156 186448
rect 357624 186396 357676 186448
rect 397736 186328 397788 186380
rect 422300 186328 422352 186380
rect 422484 186328 422536 186380
rect 267004 186260 267056 186312
rect 321652 186260 321704 186312
rect 352012 186260 352064 186312
rect 451464 186260 451516 186312
rect 451648 186260 451700 186312
rect 397736 186192 397788 186244
rect 230664 183540 230716 183592
rect 230940 183540 230992 183592
rect 252744 183540 252796 183592
rect 254308 183540 254360 183592
rect 277584 183540 277636 183592
rect 277676 183540 277728 183592
rect 287244 183540 287296 183592
rect 287428 183540 287480 183592
rect 294052 183540 294104 183592
rect 294236 183540 294288 183592
rect 295616 183583 295668 183592
rect 295616 183549 295625 183583
rect 295625 183549 295659 183583
rect 295659 183549 295668 183583
rect 295616 183540 295668 183549
rect 298376 183583 298428 183592
rect 298376 183549 298385 183583
rect 298385 183549 298419 183583
rect 298419 183549 298428 183583
rect 298376 183540 298428 183549
rect 318984 183540 319036 183592
rect 319076 183540 319128 183592
rect 331128 183540 331180 183592
rect 331496 183540 331548 183592
rect 334440 183583 334492 183592
rect 334440 183549 334449 183583
rect 334449 183549 334483 183583
rect 334483 183549 334492 183583
rect 334440 183540 334492 183549
rect 357532 183583 357584 183592
rect 357532 183549 357541 183583
rect 357541 183549 357575 183583
rect 357575 183549 357584 183583
rect 357532 183540 357584 183549
rect 381176 183540 381228 183592
rect 381360 183540 381412 183592
rect 393228 183540 393280 183592
rect 393412 183540 393464 183592
rect 408776 183540 408828 183592
rect 408960 183540 409012 183592
rect 254216 183472 254268 183524
rect 451648 183515 451700 183524
rect 451648 183481 451657 183515
rect 451657 183481 451691 183515
rect 451691 183481 451700 183515
rect 451648 183472 451700 183481
rect 466552 183472 466604 183524
rect 466644 183472 466696 183524
rect 252836 183404 252888 183456
rect 266452 183379 266504 183388
rect 266452 183345 266461 183379
rect 266461 183345 266495 183379
rect 266495 183345 266504 183379
rect 266452 183336 266504 183345
rect 386696 182180 386748 182232
rect 386788 182180 386840 182232
rect 252836 182155 252888 182164
rect 252836 182121 252845 182155
rect 252845 182121 252879 182155
rect 252879 182121 252888 182155
rect 252836 182112 252888 182121
rect 259736 182112 259788 182164
rect 259920 182112 259972 182164
rect 270592 182112 270644 182164
rect 270868 182112 270920 182164
rect 318984 182112 319036 182164
rect 319076 182112 319128 182164
rect 369952 182112 370004 182164
rect 370412 182112 370464 182164
rect 397368 182112 397420 182164
rect 397736 182112 397788 182164
rect 292764 180863 292816 180872
rect 292764 180829 292773 180863
rect 292773 180829 292807 180863
rect 292807 180829 292816 180863
rect 292764 180820 292816 180829
rect 232136 180795 232188 180804
rect 232136 180761 232145 180795
rect 232145 180761 232179 180795
rect 232179 180761 232188 180795
rect 232136 180752 232188 180761
rect 243176 180752 243228 180804
rect 243360 180752 243412 180804
rect 386696 180752 386748 180804
rect 392216 180752 392268 180804
rect 2780 179460 2832 179512
rect 4896 179460 4948 179512
rect 236368 179367 236420 179376
rect 236368 179333 236377 179367
rect 236377 179333 236411 179367
rect 236411 179333 236420 179367
rect 236368 179324 236420 179333
rect 359096 178780 359148 178832
rect 359004 178712 359056 178764
rect 254216 177284 254268 177336
rect 294052 176672 294104 176724
rect 277584 176604 277636 176656
rect 288624 176604 288676 176656
rect 298376 176740 298428 176792
rect 309416 176740 309468 176792
rect 408776 176740 408828 176792
rect 321652 176672 321704 176724
rect 327172 176672 327224 176724
rect 298284 176604 298336 176656
rect 309324 176604 309376 176656
rect 294144 176536 294196 176588
rect 321744 176536 321796 176588
rect 371424 176604 371476 176656
rect 382464 176604 382516 176656
rect 400404 176604 400456 176656
rect 400588 176604 400640 176656
rect 327264 176536 327316 176588
rect 427912 176715 427964 176724
rect 427912 176681 427921 176715
rect 427921 176681 427955 176715
rect 427955 176681 427964 176715
rect 427912 176672 427964 176681
rect 433616 176647 433668 176656
rect 433616 176613 433625 176647
rect 433625 176613 433659 176647
rect 433659 176613 433668 176647
rect 433616 176604 433668 176613
rect 408776 176536 408828 176588
rect 277584 176468 277636 176520
rect 288624 176468 288676 176520
rect 371424 176468 371476 176520
rect 382464 176468 382516 176520
rect 334348 175899 334400 175908
rect 334348 175865 334357 175899
rect 334357 175865 334391 175899
rect 334391 175865 334400 175899
rect 334348 175856 334400 175865
rect 324228 175380 324280 175432
rect 324504 175380 324556 175432
rect 230756 174360 230808 174412
rect 230940 174360 230992 174412
rect 265256 174020 265308 174072
rect 241796 173884 241848 173936
rect 241980 173884 242032 173936
rect 250076 173952 250128 174004
rect 265256 173884 265308 173936
rect 282920 173884 282972 173936
rect 283104 173884 283156 173936
rect 305184 173884 305236 173936
rect 305368 173884 305420 173936
rect 308128 173884 308180 173936
rect 308312 173884 308364 173936
rect 346584 173884 346636 173936
rect 346768 173884 346820 173936
rect 347964 173884 348016 173936
rect 348148 173884 348200 173936
rect 352012 173884 352064 173936
rect 352104 173884 352156 173936
rect 353484 173884 353536 173936
rect 353668 173884 353720 173936
rect 356428 173884 356480 173936
rect 356612 173884 356664 173936
rect 376760 173884 376812 173936
rect 376944 173884 376996 173936
rect 380808 173884 380860 173936
rect 380992 173884 381044 173936
rect 416964 173884 417016 173936
rect 417148 173884 417200 173936
rect 422484 173884 422536 173936
rect 422668 173884 422720 173936
rect 427912 173927 427964 173936
rect 427912 173893 427921 173927
rect 427921 173893 427955 173927
rect 427955 173893 427964 173927
rect 427912 173884 427964 173893
rect 433616 173927 433668 173936
rect 433616 173893 433625 173927
rect 433625 173893 433659 173927
rect 433659 173893 433668 173927
rect 433616 173884 433668 173893
rect 451740 173884 451792 173936
rect 472164 173884 472216 173936
rect 472348 173884 472400 173936
rect 249984 173816 250036 173868
rect 252836 172567 252888 172576
rect 252836 172533 252845 172567
rect 252845 172533 252879 172567
rect 252879 172533 252888 172567
rect 252836 172524 252888 172533
rect 254124 172567 254176 172576
rect 254124 172533 254133 172567
rect 254133 172533 254167 172567
rect 254167 172533 254176 172567
rect 254124 172524 254176 172533
rect 298284 172499 298336 172508
rect 298284 172465 298293 172499
rect 298293 172465 298327 172499
rect 298327 172465 298336 172499
rect 298284 172456 298336 172465
rect 309324 172499 309376 172508
rect 309324 172465 309333 172499
rect 309333 172465 309367 172499
rect 309367 172465 309376 172499
rect 309324 172456 309376 172465
rect 292764 171232 292816 171284
rect 292764 171096 292816 171148
rect 386604 171139 386656 171148
rect 386604 171105 386613 171139
rect 386613 171105 386647 171139
rect 386647 171105 386656 171139
rect 386604 171096 386656 171105
rect 392124 171139 392176 171148
rect 392124 171105 392133 171139
rect 392133 171105 392167 171139
rect 392167 171105 392176 171139
rect 392124 171096 392176 171105
rect 243084 171071 243136 171080
rect 243084 171037 243093 171071
rect 243093 171037 243127 171071
rect 243127 171037 243136 171071
rect 243084 171028 243136 171037
rect 295524 171071 295576 171080
rect 295524 171037 295533 171071
rect 295533 171037 295567 171071
rect 295567 171037 295576 171071
rect 295524 171028 295576 171037
rect 324504 171071 324556 171080
rect 324504 171037 324513 171071
rect 324513 171037 324547 171071
rect 324547 171037 324556 171071
rect 324504 171028 324556 171037
rect 238760 170280 238812 170332
rect 248328 170280 248380 170332
rect 280068 170144 280120 170196
rect 280068 169940 280120 169992
rect 289636 169940 289688 169992
rect 292948 169940 293000 169992
rect 267740 169872 267792 169924
rect 278688 169872 278740 169924
rect 475936 169872 475988 169924
rect 478144 169872 478196 169924
rect 326068 169804 326120 169856
rect 331312 169804 331364 169856
rect 425060 169804 425112 169856
rect 434536 169804 434588 169856
rect 334532 169736 334584 169788
rect 364524 167671 364576 167680
rect 364524 167637 364533 167671
rect 364533 167637 364567 167671
rect 364567 167637 364576 167671
rect 364524 167628 364576 167637
rect 270684 167016 270736 167068
rect 359004 167016 359056 167068
rect 422300 167016 422352 167068
rect 422484 167016 422536 167068
rect 230756 166948 230808 167000
rect 230940 166948 230992 167000
rect 281724 166948 281776 167000
rect 281908 166948 281960 167000
rect 298284 166991 298336 167000
rect 298284 166957 298293 166991
rect 298293 166957 298327 166991
rect 298327 166957 298336 166991
rect 298284 166948 298336 166957
rect 270776 166880 270828 166932
rect 359096 166880 359148 166932
rect 400312 164228 400364 164280
rect 400404 164228 400456 164280
rect 230664 164160 230716 164212
rect 230940 164160 230992 164212
rect 240140 164160 240192 164212
rect 240324 164160 240376 164212
rect 252560 164160 252612 164212
rect 252836 164160 252888 164212
rect 254124 164160 254176 164212
rect 254308 164160 254360 164212
rect 255504 164160 255556 164212
rect 255596 164160 255648 164212
rect 259644 164203 259696 164212
rect 259644 164169 259653 164203
rect 259653 164169 259687 164203
rect 259687 164169 259696 164203
rect 259644 164160 259696 164169
rect 272064 164160 272116 164212
rect 272248 164160 272300 164212
rect 283104 164203 283156 164212
rect 283104 164169 283113 164203
rect 283113 164169 283147 164203
rect 283147 164169 283156 164203
rect 283104 164160 283156 164169
rect 288624 164203 288676 164212
rect 288624 164169 288633 164203
rect 288633 164169 288667 164203
rect 288667 164169 288676 164203
rect 288624 164160 288676 164169
rect 305184 164160 305236 164212
rect 305276 164160 305328 164212
rect 308128 164160 308180 164212
rect 308312 164160 308364 164212
rect 309324 164203 309376 164212
rect 309324 164169 309333 164203
rect 309333 164169 309367 164203
rect 309367 164169 309376 164203
rect 309324 164160 309376 164169
rect 310704 164160 310756 164212
rect 310888 164160 310940 164212
rect 346584 164160 346636 164212
rect 346768 164160 346820 164212
rect 347964 164203 348016 164212
rect 347964 164169 347973 164203
rect 347973 164169 348007 164203
rect 348007 164169 348016 164203
rect 347964 164160 348016 164169
rect 353484 164160 353536 164212
rect 353576 164160 353628 164212
rect 356428 164160 356480 164212
rect 356520 164160 356572 164212
rect 357624 164203 357676 164212
rect 357624 164169 357633 164203
rect 357633 164169 357667 164203
rect 357667 164169 357676 164203
rect 357624 164160 357676 164169
rect 375196 164160 375248 164212
rect 375564 164160 375616 164212
rect 376760 164160 376812 164212
rect 376944 164160 376996 164212
rect 416872 164160 416924 164212
rect 417148 164160 417200 164212
rect 422392 164203 422444 164212
rect 422392 164169 422401 164203
rect 422401 164169 422435 164203
rect 422435 164169 422444 164203
rect 422392 164160 422444 164169
rect 427912 164203 427964 164212
rect 427912 164169 427921 164203
rect 427921 164169 427955 164203
rect 427955 164169 427964 164203
rect 427912 164160 427964 164169
rect 433248 164160 433300 164212
rect 433432 164160 433484 164212
rect 472072 164160 472124 164212
rect 472348 164160 472400 164212
rect 380992 164092 381044 164144
rect 381084 164092 381136 164144
rect 232136 162911 232188 162920
rect 232136 162877 232145 162911
rect 232145 162877 232179 162911
rect 232179 162877 232188 162911
rect 232136 162868 232188 162877
rect 352012 162843 352064 162852
rect 352012 162809 352021 162843
rect 352021 162809 352055 162843
rect 352055 162809 352064 162843
rect 352012 162800 352064 162809
rect 353484 162843 353536 162852
rect 353484 162809 353493 162843
rect 353493 162809 353527 162843
rect 353527 162809 353536 162843
rect 353484 162800 353536 162809
rect 356428 162843 356480 162852
rect 356428 162809 356437 162843
rect 356437 162809 356471 162843
rect 356471 162809 356480 162843
rect 356428 162800 356480 162809
rect 380992 162843 381044 162852
rect 380992 162809 381001 162843
rect 381001 162809 381035 162843
rect 381035 162809 381044 162843
rect 380992 162800 381044 162809
rect 386604 162800 386656 162852
rect 386788 162800 386840 162852
rect 387984 162843 388036 162852
rect 387984 162809 387993 162843
rect 387993 162809 388027 162843
rect 388027 162809 388036 162843
rect 387984 162800 388036 162809
rect 392124 162800 392176 162852
rect 392308 162800 392360 162852
rect 236368 161483 236420 161492
rect 236368 161449 236377 161483
rect 236377 161449 236411 161483
rect 236411 161449 236420 161483
rect 236368 161440 236420 161449
rect 243176 161440 243228 161492
rect 295524 161483 295576 161492
rect 295524 161449 295533 161483
rect 295533 161449 295567 161483
rect 295567 161449 295576 161483
rect 295524 161440 295576 161449
rect 324504 161483 324556 161492
rect 324504 161449 324513 161483
rect 324513 161449 324547 161483
rect 324547 161449 324556 161483
rect 324504 161440 324556 161449
rect 334348 161440 334400 161492
rect 334532 161440 334584 161492
rect 232136 161415 232188 161424
rect 232136 161381 232145 161415
rect 232145 161381 232179 161415
rect 232179 161381 232188 161415
rect 232136 161372 232188 161381
rect 265256 161415 265308 161424
rect 265256 161381 265265 161415
rect 265265 161381 265299 161415
rect 265299 161381 265308 161415
rect 265256 161372 265308 161381
rect 331404 161415 331456 161424
rect 331404 161381 331413 161415
rect 331413 161381 331447 161415
rect 331447 161381 331456 161415
rect 331404 161372 331456 161381
rect 287244 159332 287296 159384
rect 287428 159332 287480 159384
rect 294144 159332 294196 159384
rect 294328 159332 294380 159384
rect 294328 158652 294380 158704
rect 529664 158652 529716 158704
rect 579712 158652 579764 158704
rect 387984 158015 388036 158024
rect 387984 157981 387993 158015
rect 387993 157981 388027 158015
rect 388027 157981 388036 158015
rect 387984 157972 388036 157981
rect 243176 157428 243228 157480
rect 267004 157471 267056 157480
rect 267004 157437 267013 157471
rect 267013 157437 267047 157471
rect 267047 157437 267056 157471
rect 267004 157428 267056 157437
rect 281908 157360 281960 157412
rect 408592 157360 408644 157412
rect 243176 157292 243228 157344
rect 281816 157292 281868 157344
rect 318892 157292 318944 157344
rect 319076 157292 319128 157344
rect 336832 157292 336884 157344
rect 359096 157292 359148 157344
rect 371424 157292 371476 157344
rect 382464 157292 382516 157344
rect 336924 157224 336976 157276
rect 422392 157335 422444 157344
rect 422392 157301 422401 157335
rect 422401 157301 422435 157335
rect 422435 157301 422444 157335
rect 422392 157292 422444 157301
rect 427912 157335 427964 157344
rect 427912 157301 427921 157335
rect 427921 157301 427955 157335
rect 427955 157301 427964 157335
rect 427912 157292 427964 157301
rect 451648 157292 451700 157344
rect 408684 157224 408736 157276
rect 371424 157156 371476 157208
rect 382464 157156 382516 157208
rect 451648 157156 451700 157208
rect 347964 155771 348016 155780
rect 347964 155737 347973 155771
rect 347973 155737 348007 155771
rect 348007 155737 348016 155771
rect 347964 155728 348016 155737
rect 283104 154955 283156 154964
rect 283104 154921 283113 154955
rect 283113 154921 283147 154955
rect 283147 154921 283156 154955
rect 283104 154912 283156 154921
rect 288624 154955 288676 154964
rect 288624 154921 288633 154955
rect 288633 154921 288667 154955
rect 288667 154921 288676 154955
rect 288624 154912 288676 154921
rect 259644 154615 259696 154624
rect 259644 154581 259653 154615
rect 259653 154581 259687 154615
rect 259687 154581 259696 154615
rect 259644 154572 259696 154581
rect 357624 154615 357676 154624
rect 357624 154581 357633 154615
rect 357633 154581 357667 154615
rect 357667 154581 357676 154615
rect 357624 154572 357676 154581
rect 359004 154615 359056 154624
rect 359004 154581 359013 154615
rect 359013 154581 359047 154615
rect 359047 154581 359056 154615
rect 359004 154572 359056 154581
rect 364616 154572 364668 154624
rect 466552 154572 466604 154624
rect 466644 154572 466696 154624
rect 230848 154504 230900 154556
rect 231032 154504 231084 154556
rect 270684 154547 270736 154556
rect 270684 154513 270693 154547
rect 270693 154513 270727 154547
rect 270727 154513 270736 154547
rect 270684 154504 270736 154513
rect 271788 154504 271840 154556
rect 272064 154504 272116 154556
rect 342352 154504 342404 154556
rect 342536 154504 342588 154556
rect 352012 154547 352064 154556
rect 352012 154513 352021 154547
rect 352021 154513 352055 154547
rect 352055 154513 352064 154547
rect 352012 154504 352064 154513
rect 370044 154547 370096 154556
rect 370044 154513 370053 154547
rect 370053 154513 370087 154547
rect 370087 154513 370096 154547
rect 370044 154504 370096 154513
rect 375564 154504 375616 154556
rect 375748 154504 375800 154556
rect 393228 154504 393280 154556
rect 393412 154504 393464 154556
rect 408684 154547 408736 154556
rect 408684 154513 408693 154547
rect 408693 154513 408727 154547
rect 408727 154513 408736 154547
rect 408684 154504 408736 154513
rect 451648 154547 451700 154556
rect 451648 154513 451657 154547
rect 451657 154513 451691 154547
rect 451691 154513 451700 154547
rect 451648 154504 451700 154513
rect 466552 154479 466604 154488
rect 466552 154445 466561 154479
rect 466561 154445 466595 154479
rect 466595 154445 466604 154479
rect 466552 154436 466604 154445
rect 353484 153255 353536 153264
rect 353484 153221 353493 153255
rect 353493 153221 353527 153255
rect 353527 153221 353536 153255
rect 353484 153212 353536 153221
rect 356428 153255 356480 153264
rect 356428 153221 356437 153255
rect 356437 153221 356471 153255
rect 356471 153221 356480 153255
rect 356428 153212 356480 153221
rect 236276 153144 236328 153196
rect 236368 153144 236420 153196
rect 240140 153144 240192 153196
rect 240232 153144 240284 153196
rect 267004 153187 267056 153196
rect 267004 153153 267013 153187
rect 267013 153153 267047 153187
rect 267047 153153 267056 153187
rect 267004 153144 267056 153153
rect 309324 153144 309376 153196
rect 309508 153144 309560 153196
rect 318984 153144 319036 153196
rect 319076 153144 319128 153196
rect 321744 153187 321796 153196
rect 321744 153153 321753 153187
rect 321753 153153 321787 153187
rect 321787 153153 321796 153187
rect 321744 153144 321796 153153
rect 347964 153187 348016 153196
rect 347964 153153 347973 153187
rect 347973 153153 348007 153187
rect 348007 153153 348016 153187
rect 347964 153144 348016 153153
rect 400496 153187 400548 153196
rect 400496 153153 400505 153187
rect 400505 153153 400539 153187
rect 400539 153153 400548 153187
rect 400496 153144 400548 153153
rect 353484 153119 353536 153128
rect 353484 153085 353493 153119
rect 353493 153085 353527 153119
rect 353527 153085 353536 153119
rect 353484 153076 353536 153085
rect 232228 151784 232280 151836
rect 265256 151827 265308 151836
rect 265256 151793 265265 151827
rect 265265 151793 265299 151827
rect 265299 151793 265308 151827
rect 265256 151784 265308 151793
rect 295616 151784 295668 151836
rect 331404 151827 331456 151836
rect 292764 151759 292816 151768
rect 292764 151725 292773 151759
rect 292773 151725 292807 151759
rect 292807 151725 292816 151759
rect 292764 151716 292816 151725
rect 331404 151793 331413 151827
rect 331413 151793 331447 151827
rect 331447 151793 331456 151827
rect 331404 151784 331456 151793
rect 324596 151759 324648 151768
rect 324596 151725 324605 151759
rect 324605 151725 324639 151759
rect 324639 151725 324648 151759
rect 324596 151716 324648 151725
rect 295708 151648 295760 151700
rect 295708 150356 295760 150408
rect 351828 149676 351880 149728
rect 352012 149676 352064 149728
rect 294052 149107 294104 149116
rect 294052 149073 294061 149107
rect 294061 149073 294095 149107
rect 294095 149073 294104 149107
rect 294052 149064 294104 149073
rect 392308 148316 392360 148368
rect 331404 147704 331456 147756
rect 334348 147704 334400 147756
rect 359004 147704 359056 147756
rect 259644 147636 259696 147688
rect 327264 147636 327316 147688
rect 356428 147636 356480 147688
rect 259736 147568 259788 147620
rect 270684 147611 270736 147620
rect 270684 147577 270693 147611
rect 270693 147577 270727 147611
rect 270727 147577 270736 147611
rect 270684 147568 270736 147577
rect 327172 147568 327224 147620
rect 331404 147568 331456 147620
rect 334348 147568 334400 147620
rect 422300 147636 422352 147688
rect 422484 147636 422536 147688
rect 427820 147636 427872 147688
rect 428004 147636 428056 147688
rect 359004 147568 359056 147620
rect 370044 147611 370096 147620
rect 370044 147577 370053 147611
rect 370053 147577 370087 147611
rect 370087 147577 370096 147611
rect 370044 147568 370096 147577
rect 381084 147568 381136 147620
rect 400496 147611 400548 147620
rect 400496 147577 400505 147611
rect 400505 147577 400539 147611
rect 400539 147577 400548 147611
rect 400496 147568 400548 147577
rect 408684 147611 408736 147620
rect 408684 147577 408693 147611
rect 408693 147577 408727 147611
rect 408727 147577 408736 147611
rect 408684 147568 408736 147577
rect 451648 147611 451700 147620
rect 451648 147577 451657 147611
rect 451657 147577 451691 147611
rect 451691 147577 451700 147611
rect 451648 147568 451700 147577
rect 466552 147611 466604 147620
rect 466552 147577 466561 147611
rect 466561 147577 466595 147611
rect 466595 147577 466604 147611
rect 466552 147568 466604 147577
rect 356520 147432 356572 147484
rect 252560 145528 252612 145580
rect 252744 145528 252796 145580
rect 357624 144916 357676 144968
rect 357716 144916 357768 144968
rect 254216 144848 254268 144900
rect 254308 144848 254360 144900
rect 259736 144848 259788 144900
rect 259828 144848 259880 144900
rect 271972 144848 272024 144900
rect 272064 144848 272116 144900
rect 308128 144848 308180 144900
rect 308312 144848 308364 144900
rect 310704 144848 310756 144900
rect 310888 144848 310940 144900
rect 334440 144848 334492 144900
rect 346584 144848 346636 144900
rect 346768 144848 346820 144900
rect 352012 144848 352064 144900
rect 352196 144848 352248 144900
rect 356520 144848 356572 144900
rect 356612 144848 356664 144900
rect 364616 144848 364668 144900
rect 364708 144848 364760 144900
rect 376760 144848 376812 144900
rect 376944 144848 376996 144900
rect 393228 144891 393280 144900
rect 393228 144857 393237 144891
rect 393237 144857 393271 144891
rect 393271 144857 393280 144891
rect 393228 144848 393280 144857
rect 422392 144891 422444 144900
rect 422392 144857 422401 144891
rect 422401 144857 422435 144891
rect 422435 144857 422444 144891
rect 422392 144848 422444 144857
rect 433616 144848 433668 144900
rect 433800 144848 433852 144900
rect 347964 144823 348016 144832
rect 347964 144789 347973 144823
rect 347973 144789 348007 144823
rect 348007 144789 348016 144823
rect 347964 144780 348016 144789
rect 353484 144823 353536 144832
rect 353484 144789 353493 144823
rect 353493 144789 353527 144823
rect 353527 144789 353536 144823
rect 353484 144780 353536 144789
rect 267004 143556 267056 143608
rect 267096 143556 267148 143608
rect 321744 143599 321796 143608
rect 321744 143565 321753 143599
rect 321753 143565 321787 143599
rect 321787 143565 321796 143599
rect 321744 143556 321796 143565
rect 231952 143488 232004 143540
rect 232044 143488 232096 143540
rect 236276 143488 236328 143540
rect 236460 143488 236512 143540
rect 357532 143488 357584 143540
rect 357624 143488 357676 143540
rect 397736 143531 397788 143540
rect 397736 143497 397745 143531
rect 397745 143497 397779 143531
rect 397779 143497 397788 143531
rect 397736 143488 397788 143497
rect 400404 143488 400456 143540
rect 400496 143488 400548 143540
rect 472072 143531 472124 143540
rect 472072 143497 472081 143531
rect 472081 143497 472115 143531
rect 472115 143497 472124 143531
rect 472072 143488 472124 143497
rect 292764 142171 292816 142180
rect 292764 142137 292773 142171
rect 292773 142137 292807 142171
rect 292807 142137 292816 142171
rect 292764 142128 292816 142137
rect 324596 142171 324648 142180
rect 324596 142137 324605 142171
rect 324605 142137 324639 142171
rect 324639 142137 324648 142171
rect 324596 142128 324648 142137
rect 232044 142060 232096 142112
rect 236460 142103 236512 142112
rect 236460 142069 236469 142103
rect 236469 142069 236503 142103
rect 236503 142069 236512 142103
rect 236460 142060 236512 142069
rect 240140 142103 240192 142112
rect 240140 142069 240149 142103
rect 240149 142069 240183 142103
rect 240183 142069 240192 142103
rect 240140 142060 240192 142069
rect 266452 142103 266504 142112
rect 266452 142069 266461 142103
rect 266461 142069 266495 142103
rect 266495 142069 266504 142103
rect 266452 142060 266504 142069
rect 295616 140811 295668 140820
rect 295616 140777 295625 140811
rect 295625 140777 295659 140811
rect 295659 140777 295668 140811
rect 295616 140768 295668 140777
rect 294052 139383 294104 139392
rect 294052 139349 294061 139383
rect 294061 139349 294095 139383
rect 294095 139349 294104 139383
rect 294052 139340 294104 139349
rect 277584 138048 277636 138100
rect 342536 138048 342588 138100
rect 230756 137980 230808 138032
rect 244464 137980 244516 138032
rect 249984 137980 250036 138032
rect 230848 137912 230900 137964
rect 318984 137980 319036 138032
rect 277584 137912 277636 137964
rect 408776 138048 408828 138100
rect 428004 138048 428056 138100
rect 416872 137980 416924 138032
rect 466460 137980 466512 138032
rect 466644 137980 466696 138032
rect 319076 137912 319128 137964
rect 342536 137912 342588 137964
rect 397736 137955 397788 137964
rect 397736 137921 397745 137955
rect 397745 137921 397779 137955
rect 397779 137921 397788 137955
rect 397736 137912 397788 137921
rect 408684 137912 408736 137964
rect 416780 137912 416832 137964
rect 422392 137955 422444 137964
rect 422392 137921 422401 137955
rect 422401 137921 422435 137955
rect 422435 137921 422444 137955
rect 422392 137912 422444 137921
rect 244464 137844 244516 137896
rect 249984 137844 250036 137896
rect 359004 135328 359056 135380
rect 309324 135260 309376 135312
rect 309600 135260 309652 135312
rect 327172 135303 327224 135312
rect 327172 135269 327181 135303
rect 327181 135269 327215 135303
rect 327215 135269 327224 135303
rect 327172 135260 327224 135269
rect 381084 135260 381136 135312
rect 381268 135260 381320 135312
rect 392124 135303 392176 135312
rect 392124 135269 392133 135303
rect 392133 135269 392167 135303
rect 392167 135269 392176 135303
rect 392124 135260 392176 135269
rect 393228 135303 393280 135312
rect 393228 135269 393237 135303
rect 393237 135269 393271 135303
rect 393271 135269 393280 135303
rect 393228 135260 393280 135269
rect 427912 135303 427964 135312
rect 427912 135269 427921 135303
rect 427921 135269 427955 135303
rect 427955 135269 427964 135303
rect 427912 135260 427964 135269
rect 451648 135260 451700 135312
rect 451740 135260 451792 135312
rect 230848 135192 230900 135244
rect 231032 135192 231084 135244
rect 259644 135192 259696 135244
rect 259828 135192 259880 135244
rect 270684 135235 270736 135244
rect 270684 135201 270693 135235
rect 270693 135201 270727 135235
rect 270727 135201 270736 135235
rect 270684 135192 270736 135201
rect 281632 135235 281684 135244
rect 281632 135201 281641 135235
rect 281641 135201 281675 135235
rect 281675 135201 281684 135235
rect 281632 135192 281684 135201
rect 352104 135192 352156 135244
rect 352196 135192 352248 135244
rect 356428 135192 356480 135244
rect 359004 135192 359056 135244
rect 370044 135235 370096 135244
rect 370044 135201 370053 135235
rect 370053 135201 370087 135235
rect 370087 135201 370096 135235
rect 370044 135192 370096 135201
rect 375564 135192 375616 135244
rect 408684 135235 408736 135244
rect 408684 135201 408693 135235
rect 408693 135201 408727 135235
rect 408727 135201 408736 135235
rect 408684 135192 408736 135201
rect 334440 135124 334492 135176
rect 356520 135124 356572 135176
rect 375748 135124 375800 135176
rect 284300 134036 284352 134088
rect 293776 134036 293828 134088
rect 514576 134036 514628 134088
rect 514852 134036 514904 134088
rect 540980 133900 541032 133952
rect 545856 133900 545908 133952
rect 243084 133875 243136 133884
rect 243084 133841 243093 133875
rect 243093 133841 243127 133875
rect 243127 133841 243136 133875
rect 243084 133832 243136 133841
rect 325608 133832 325660 133884
rect 333888 133832 333940 133884
rect 298376 133807 298428 133816
rect 298376 133773 298385 133807
rect 298385 133773 298419 133807
rect 298419 133773 298428 133807
rect 298376 133764 298428 133773
rect 348424 133696 348476 133748
rect 354588 133696 354640 133748
rect 236460 132515 236512 132524
rect 236460 132481 236469 132515
rect 236469 132481 236503 132515
rect 236503 132481 236512 132515
rect 236460 132472 236512 132481
rect 240324 132472 240376 132524
rect 266544 132472 266596 132524
rect 327172 132515 327224 132524
rect 327172 132481 327181 132515
rect 327181 132481 327215 132515
rect 327215 132481 327224 132515
rect 327172 132472 327224 132481
rect 265348 132447 265400 132456
rect 265348 132413 265357 132447
rect 265357 132413 265391 132447
rect 265391 132413 265400 132447
rect 265348 132404 265400 132413
rect 309324 132447 309376 132456
rect 309324 132413 309333 132447
rect 309333 132413 309367 132447
rect 309367 132413 309376 132447
rect 309324 132404 309376 132413
rect 321744 132447 321796 132456
rect 321744 132413 321753 132447
rect 321753 132413 321787 132447
rect 321787 132413 321796 132447
rect 321744 132404 321796 132413
rect 324504 132404 324556 132456
rect 295524 131087 295576 131096
rect 295524 131053 295533 131087
rect 295533 131053 295567 131087
rect 295567 131053 295576 131087
rect 295524 131044 295576 131053
rect 271972 130364 272024 130416
rect 272156 130364 272208 130416
rect 281816 129004 281868 129056
rect 233332 128324 233384 128376
rect 233516 128324 233568 128376
rect 381084 128324 381136 128376
rect 400404 128324 400456 128376
rect 422300 128324 422352 128376
rect 422484 128324 422536 128376
rect 466460 128324 466512 128376
rect 270684 128299 270736 128308
rect 270684 128265 270693 128299
rect 270693 128265 270727 128299
rect 270727 128265 270736 128299
rect 270684 128256 270736 128265
rect 370044 128299 370096 128308
rect 370044 128265 370053 128299
rect 370053 128265 370087 128299
rect 370087 128265 370096 128299
rect 370044 128256 370096 128265
rect 381176 128256 381228 128308
rect 400496 128256 400548 128308
rect 408684 128299 408736 128308
rect 408684 128265 408693 128299
rect 408693 128265 408727 128299
rect 408727 128265 408736 128299
rect 408684 128256 408736 128265
rect 466552 128256 466604 128308
rect 472072 128299 472124 128308
rect 472072 128265 472081 128299
rect 472081 128265 472115 128299
rect 472115 128265 472124 128299
rect 472072 128256 472124 128265
rect 241796 125536 241848 125588
rect 241980 125536 242032 125588
rect 252744 125536 252796 125588
rect 252928 125536 252980 125588
rect 254216 125536 254268 125588
rect 254308 125536 254360 125588
rect 255504 125536 255556 125588
rect 255596 125536 255648 125588
rect 259736 125536 259788 125588
rect 259828 125536 259880 125588
rect 266544 125536 266596 125588
rect 266728 125536 266780 125588
rect 267004 125536 267056 125588
rect 267280 125536 267332 125588
rect 283104 125579 283156 125588
rect 283104 125545 283113 125579
rect 283113 125545 283147 125579
rect 283147 125545 283156 125579
rect 283104 125536 283156 125545
rect 308128 125536 308180 125588
rect 308312 125536 308364 125588
rect 310704 125579 310756 125588
rect 310704 125545 310713 125579
rect 310713 125545 310747 125579
rect 310747 125545 310756 125579
rect 310704 125536 310756 125545
rect 346584 125579 346636 125588
rect 346584 125545 346593 125579
rect 346593 125545 346627 125579
rect 346627 125545 346636 125579
rect 346584 125536 346636 125545
rect 352012 125536 352064 125588
rect 352196 125536 352248 125588
rect 357624 125536 357676 125588
rect 357716 125536 357768 125588
rect 364616 125536 364668 125588
rect 376944 125579 376996 125588
rect 376944 125545 376953 125579
rect 376953 125545 376987 125579
rect 376987 125545 376996 125579
rect 376944 125536 376996 125545
rect 386696 125536 386748 125588
rect 386788 125536 386840 125588
rect 387984 125536 388036 125588
rect 388076 125536 388128 125588
rect 392216 125536 392268 125588
rect 392308 125536 392360 125588
rect 393228 125579 393280 125588
rect 393228 125545 393237 125579
rect 393237 125545 393271 125579
rect 393271 125545 393280 125579
rect 393228 125536 393280 125545
rect 422392 125579 422444 125588
rect 422392 125545 422401 125579
rect 422401 125545 422435 125579
rect 422435 125545 422444 125579
rect 422392 125536 422444 125545
rect 427912 125579 427964 125588
rect 427912 125545 427921 125579
rect 427921 125545 427955 125579
rect 427955 125545 427964 125579
rect 427912 125536 427964 125545
rect 433616 125579 433668 125588
rect 433616 125545 433625 125579
rect 433625 125545 433659 125579
rect 433659 125545 433668 125579
rect 433616 125536 433668 125545
rect 466644 125536 466696 125588
rect 466736 125536 466788 125588
rect 265348 124627 265400 124636
rect 265348 124593 265357 124627
rect 265357 124593 265391 124627
rect 265391 124593 265400 124627
rect 265348 124584 265400 124593
rect 236368 124244 236420 124296
rect 236460 124244 236512 124296
rect 231952 124219 232004 124228
rect 231952 124185 231961 124219
rect 231961 124185 231995 124219
rect 231995 124185 232004 124219
rect 231952 124176 232004 124185
rect 243268 124176 243320 124228
rect 298376 124219 298428 124228
rect 298376 124185 298385 124219
rect 298385 124185 298419 124219
rect 298419 124185 298428 124219
rect 298376 124176 298428 124185
rect 356428 124176 356480 124228
rect 356520 124176 356572 124228
rect 400496 124108 400548 124160
rect 451464 124151 451516 124160
rect 451464 124117 451473 124151
rect 451473 124117 451507 124151
rect 451507 124117 451516 124151
rect 451464 124108 451516 124117
rect 466736 124108 466788 124160
rect 309508 122816 309560 122868
rect 321744 122859 321796 122868
rect 321744 122825 321753 122859
rect 321753 122825 321787 122859
rect 321787 122825 321796 122859
rect 321744 122816 321796 122825
rect 324412 122859 324464 122868
rect 324412 122825 324421 122859
rect 324421 122825 324455 122859
rect 324455 122825 324464 122859
rect 324412 122816 324464 122825
rect 236368 122791 236420 122800
rect 236368 122757 236377 122791
rect 236377 122757 236411 122791
rect 236411 122757 236420 122791
rect 236368 122748 236420 122757
rect 294144 121456 294196 121508
rect 295616 121456 295668 121508
rect 294144 121363 294196 121372
rect 294144 121329 294153 121363
rect 294153 121329 294187 121363
rect 294187 121329 294196 121363
rect 294144 121320 294196 121329
rect 270776 120708 270828 120760
rect 305276 120708 305328 120760
rect 370136 120708 370188 120760
rect 375472 120708 375524 120760
rect 375748 120708 375800 120760
rect 270776 120572 270828 120624
rect 370136 120572 370188 120624
rect 298376 119391 298428 119400
rect 298376 119357 298385 119391
rect 298385 119357 298419 119391
rect 298419 119357 298428 119391
rect 298376 119348 298428 119357
rect 261024 118736 261076 118788
rect 295616 118736 295668 118788
rect 318984 118779 319036 118788
rect 318984 118745 318993 118779
rect 318993 118745 319027 118779
rect 319027 118745 319036 118779
rect 318984 118736 319036 118745
rect 321744 118736 321796 118788
rect 230756 118668 230808 118720
rect 336924 118736 336976 118788
rect 336832 118668 336884 118720
rect 408776 118736 408828 118788
rect 416872 118668 416924 118720
rect 472072 118668 472124 118720
rect 230848 118600 230900 118652
rect 261024 118600 261076 118652
rect 295616 118600 295668 118652
rect 321744 118600 321796 118652
rect 387984 118600 388036 118652
rect 388076 118600 388128 118652
rect 408684 118600 408736 118652
rect 416780 118600 416832 118652
rect 422392 118643 422444 118652
rect 422392 118609 422401 118643
rect 422401 118609 422435 118643
rect 422435 118609 422444 118643
rect 422392 118600 422444 118609
rect 427912 118643 427964 118652
rect 427912 118609 427921 118643
rect 427921 118609 427955 118643
rect 427955 118609 427964 118643
rect 427912 118600 427964 118609
rect 433616 118643 433668 118652
rect 433616 118609 433625 118643
rect 433625 118609 433659 118643
rect 433659 118609 433668 118643
rect 433616 118600 433668 118609
rect 471980 118600 472032 118652
rect 324228 117988 324280 118040
rect 324412 117988 324464 118040
rect 294144 116603 294196 116612
rect 294144 116569 294153 116603
rect 294153 116569 294187 116603
rect 294187 116569 294196 116603
rect 294144 116560 294196 116569
rect 272064 115948 272116 116000
rect 272156 115948 272208 116000
rect 283104 115991 283156 116000
rect 283104 115957 283113 115991
rect 283113 115957 283147 115991
rect 283147 115957 283156 115991
rect 283104 115948 283156 115957
rect 305184 115991 305236 116000
rect 305184 115957 305193 115991
rect 305193 115957 305227 115991
rect 305227 115957 305236 115991
rect 305184 115948 305236 115957
rect 310704 115991 310756 116000
rect 310704 115957 310713 115991
rect 310713 115957 310747 115991
rect 310747 115957 310756 115991
rect 310704 115948 310756 115957
rect 346584 115991 346636 116000
rect 346584 115957 346593 115991
rect 346593 115957 346627 115991
rect 346627 115957 346636 115991
rect 346584 115948 346636 115957
rect 353576 115991 353628 116000
rect 353576 115957 353585 115991
rect 353585 115957 353619 115991
rect 353619 115957 353628 115991
rect 353576 115948 353628 115957
rect 364524 115991 364576 116000
rect 364524 115957 364533 115991
rect 364533 115957 364567 115991
rect 364567 115957 364576 115991
rect 364524 115948 364576 115957
rect 376944 115991 376996 116000
rect 376944 115957 376953 115991
rect 376953 115957 376987 115991
rect 376987 115957 376996 115991
rect 376944 115948 376996 115957
rect 393228 115991 393280 116000
rect 393228 115957 393237 115991
rect 393237 115957 393271 115991
rect 393271 115957 393280 115991
rect 393228 115948 393280 115957
rect 230848 115880 230900 115932
rect 231032 115880 231084 115932
rect 254124 115923 254176 115932
rect 254124 115889 254133 115923
rect 254133 115889 254167 115923
rect 254167 115889 254176 115923
rect 254124 115880 254176 115889
rect 259644 115880 259696 115932
rect 259828 115880 259880 115932
rect 265164 115880 265216 115932
rect 265256 115880 265308 115932
rect 342444 115923 342496 115932
rect 342444 115889 342453 115923
rect 342453 115889 342487 115923
rect 342487 115889 342496 115923
rect 342444 115880 342496 115889
rect 347964 115880 348016 115932
rect 348056 115880 348108 115932
rect 356428 115880 356480 115932
rect 356612 115880 356664 115932
rect 375472 115880 375524 115932
rect 375748 115880 375800 115932
rect 381084 115880 381136 115932
rect 381268 115880 381320 115932
rect 386604 115880 386656 115932
rect 386788 115880 386840 115932
rect 392124 115880 392176 115932
rect 392308 115880 392360 115932
rect 393228 115812 393280 115864
rect 393320 115812 393372 115864
rect 298192 114520 298244 114572
rect 334440 114520 334492 114572
rect 353576 114563 353628 114572
rect 353576 114529 353585 114563
rect 353585 114529 353619 114563
rect 353619 114529 353628 114563
rect 353576 114520 353628 114529
rect 400312 114563 400364 114572
rect 400312 114529 400321 114563
rect 400321 114529 400355 114563
rect 400355 114529 400364 114563
rect 400312 114520 400364 114529
rect 451556 114520 451608 114572
rect 466644 114563 466696 114572
rect 466644 114529 466653 114563
rect 466653 114529 466687 114563
rect 466687 114529 466696 114563
rect 466644 114520 466696 114529
rect 267096 114452 267148 114504
rect 327172 114495 327224 114504
rect 327172 114461 327181 114495
rect 327181 114461 327215 114495
rect 327215 114461 327224 114495
rect 327172 114452 327224 114461
rect 356612 114452 356664 114504
rect 387984 114495 388036 114504
rect 387984 114461 387993 114495
rect 387993 114461 388027 114495
rect 388027 114461 388036 114495
rect 387984 114452 388036 114461
rect 298192 114427 298244 114436
rect 298192 114393 298201 114427
rect 298201 114393 298235 114427
rect 298235 114393 298244 114427
rect 298192 114384 298244 114393
rect 236460 113160 236512 113212
rect 309324 113160 309376 113212
rect 309508 113160 309560 113212
rect 334348 113203 334400 113212
rect 334348 113169 334357 113203
rect 334357 113169 334391 113203
rect 334391 113169 334400 113203
rect 334348 113160 334400 113169
rect 292764 113135 292816 113144
rect 292764 113101 292773 113135
rect 292773 113101 292807 113135
rect 292807 113101 292816 113135
rect 292764 113092 292816 113101
rect 295616 111775 295668 111784
rect 295616 111741 295625 111775
rect 295625 111741 295659 111775
rect 295659 111741 295668 111775
rect 295616 111732 295668 111741
rect 529572 111732 529624 111784
rect 580172 111732 580224 111784
rect 397644 109080 397696 109132
rect 233332 109012 233384 109064
rect 233516 109012 233568 109064
rect 243084 109012 243136 109064
rect 370136 109055 370188 109064
rect 370136 109021 370145 109055
rect 370145 109021 370179 109055
rect 370179 109021 370188 109055
rect 370136 109012 370188 109021
rect 408684 109012 408736 109064
rect 422300 109012 422352 109064
rect 422484 109012 422536 109064
rect 427820 109012 427872 109064
rect 428004 109012 428056 109064
rect 243176 108944 243228 108996
rect 254124 108987 254176 108996
rect 254124 108953 254133 108987
rect 254133 108953 254167 108987
rect 254167 108953 254176 108987
rect 254124 108944 254176 108953
rect 342444 108987 342496 108996
rect 342444 108953 342453 108987
rect 342453 108953 342487 108987
rect 342487 108953 342496 108987
rect 342444 108944 342496 108953
rect 397644 108944 397696 108996
rect 466644 109012 466696 109064
rect 408776 108944 408828 108996
rect 466552 108944 466604 108996
rect 370136 106335 370188 106344
rect 370136 106301 370145 106335
rect 370145 106301 370179 106335
rect 370179 106301 370188 106335
rect 370136 106292 370188 106301
rect 241796 106224 241848 106276
rect 241980 106224 242032 106276
rect 254124 106224 254176 106276
rect 254216 106224 254268 106276
rect 281816 106224 281868 106276
rect 281908 106224 281960 106276
rect 283104 106267 283156 106276
rect 283104 106233 283113 106267
rect 283113 106233 283147 106267
rect 283147 106233 283156 106267
rect 283104 106224 283156 106233
rect 305184 106267 305236 106276
rect 305184 106233 305193 106267
rect 305193 106233 305227 106267
rect 305227 106233 305236 106267
rect 305184 106224 305236 106233
rect 308036 106224 308088 106276
rect 308220 106224 308272 106276
rect 310704 106267 310756 106276
rect 310704 106233 310713 106267
rect 310713 106233 310747 106267
rect 310747 106233 310756 106267
rect 310704 106224 310756 106233
rect 330024 106224 330076 106276
rect 330208 106224 330260 106276
rect 331404 106224 331456 106276
rect 331496 106224 331548 106276
rect 346584 106267 346636 106276
rect 346584 106233 346593 106267
rect 346593 106233 346627 106267
rect 346627 106233 346636 106267
rect 346584 106224 346636 106233
rect 352012 106224 352064 106276
rect 352196 106224 352248 106276
rect 353484 106224 353536 106276
rect 353576 106224 353628 106276
rect 364524 106224 364576 106276
rect 364616 106224 364668 106276
rect 376944 106267 376996 106276
rect 376944 106233 376953 106267
rect 376953 106233 376987 106267
rect 376987 106233 376996 106267
rect 376944 106224 376996 106233
rect 393228 106224 393280 106276
rect 393412 106224 393464 106276
rect 422392 106267 422444 106276
rect 422392 106233 422401 106267
rect 422401 106233 422435 106267
rect 422435 106233 422444 106267
rect 422392 106224 422444 106233
rect 427912 106267 427964 106276
rect 427912 106233 427921 106267
rect 427921 106233 427955 106267
rect 427955 106233 427964 106267
rect 427912 106224 427964 106233
rect 231952 106156 232004 106208
rect 232136 106156 232188 106208
rect 236276 106156 236328 106208
rect 236552 106156 236604 106208
rect 243176 106199 243228 106208
rect 243176 106165 243185 106199
rect 243185 106165 243219 106199
rect 243219 106165 243228 106199
rect 243176 106156 243228 106165
rect 252744 106199 252796 106208
rect 252744 106165 252753 106199
rect 252753 106165 252787 106199
rect 252787 106165 252796 106199
rect 252744 106156 252796 106165
rect 267004 104975 267056 104984
rect 267004 104941 267013 104975
rect 267013 104941 267047 104975
rect 267047 104941 267056 104975
rect 267004 104932 267056 104941
rect 356428 104975 356480 104984
rect 356428 104941 356437 104975
rect 356437 104941 356471 104975
rect 356471 104941 356480 104975
rect 356428 104932 356480 104941
rect 298376 104864 298428 104916
rect 318984 104907 319036 104916
rect 318984 104873 318993 104907
rect 318993 104873 319027 104907
rect 319027 104873 319036 104907
rect 318984 104864 319036 104873
rect 327264 104864 327316 104916
rect 334348 104864 334400 104916
rect 334440 104864 334492 104916
rect 387984 104907 388036 104916
rect 387984 104873 387993 104907
rect 387993 104873 388027 104907
rect 388027 104873 388036 104907
rect 387984 104864 388036 104873
rect 232136 104839 232188 104848
rect 232136 104805 232145 104839
rect 232145 104805 232179 104839
rect 232179 104805 232188 104839
rect 232136 104796 232188 104805
rect 267004 104839 267056 104848
rect 267004 104805 267013 104839
rect 267013 104805 267047 104839
rect 267047 104805 267056 104839
rect 267004 104796 267056 104805
rect 324412 104796 324464 104848
rect 324688 104796 324740 104848
rect 353484 104839 353536 104848
rect 353484 104805 353493 104839
rect 353493 104805 353527 104839
rect 353527 104805 353536 104839
rect 353484 104796 353536 104805
rect 356428 104839 356480 104848
rect 356428 104805 356437 104839
rect 356437 104805 356471 104839
rect 356471 104805 356480 104839
rect 356428 104796 356480 104805
rect 408776 104796 408828 104848
rect 451556 104839 451608 104848
rect 451556 104805 451565 104839
rect 451565 104805 451599 104839
rect 451599 104805 451608 104839
rect 451556 104796 451608 104805
rect 292764 103615 292816 103624
rect 292764 103581 292773 103615
rect 292773 103581 292807 103615
rect 292807 103581 292816 103615
rect 292764 103572 292816 103581
rect 292764 103436 292816 103488
rect 334440 103436 334492 103488
rect 295708 102144 295760 102196
rect 270868 102119 270920 102128
rect 270868 102085 270877 102119
rect 270877 102085 270911 102119
rect 270911 102085 270920 102119
rect 270868 102076 270920 102085
rect 260840 100036 260892 100088
rect 261024 100036 261076 100088
rect 327264 99492 327316 99544
rect 298376 99467 298428 99476
rect 298376 99433 298385 99467
rect 298385 99433 298419 99467
rect 298419 99433 298428 99467
rect 298376 99424 298428 99433
rect 321744 99424 321796 99476
rect 230756 99356 230808 99408
rect 277584 99356 277636 99408
rect 318984 99356 319036 99408
rect 230848 99288 230900 99340
rect 277676 99288 277728 99340
rect 416872 99356 416924 99408
rect 466552 99356 466604 99408
rect 472072 99356 472124 99408
rect 319076 99288 319128 99340
rect 321744 99288 321796 99340
rect 327264 99288 327316 99340
rect 416780 99288 416832 99340
rect 422392 99331 422444 99340
rect 422392 99297 422401 99331
rect 422401 99297 422435 99331
rect 422435 99297 422444 99331
rect 422392 99288 422444 99297
rect 427912 99331 427964 99340
rect 427912 99297 427921 99331
rect 427921 99297 427955 99331
rect 427955 99297 427964 99331
rect 427912 99288 427964 99297
rect 466460 99288 466512 99340
rect 471980 99288 472032 99340
rect 243176 96747 243228 96756
rect 243176 96713 243185 96747
rect 243185 96713 243219 96747
rect 243219 96713 243228 96747
rect 243176 96704 243228 96713
rect 252744 96679 252796 96688
rect 252744 96645 252753 96679
rect 252753 96645 252787 96679
rect 252787 96645 252796 96679
rect 252744 96636 252796 96645
rect 283104 96679 283156 96688
rect 283104 96645 283113 96679
rect 283113 96645 283147 96679
rect 283147 96645 283156 96679
rect 283104 96636 283156 96645
rect 305184 96679 305236 96688
rect 305184 96645 305193 96679
rect 305193 96645 305227 96679
rect 305227 96645 305236 96679
rect 305184 96636 305236 96645
rect 310704 96679 310756 96688
rect 310704 96645 310713 96679
rect 310713 96645 310747 96679
rect 310747 96645 310756 96679
rect 310704 96636 310756 96645
rect 346584 96679 346636 96688
rect 346584 96645 346593 96679
rect 346593 96645 346627 96679
rect 346627 96645 346636 96679
rect 346584 96636 346636 96645
rect 376944 96679 376996 96688
rect 376944 96645 376953 96679
rect 376953 96645 376987 96679
rect 376987 96645 376996 96679
rect 376944 96636 376996 96645
rect 230848 96611 230900 96620
rect 230848 96577 230857 96611
rect 230857 96577 230891 96611
rect 230891 96577 230900 96611
rect 230848 96568 230900 96577
rect 243084 96568 243136 96620
rect 243176 96568 243228 96620
rect 281816 96568 281868 96620
rect 282000 96568 282052 96620
rect 232228 95208 232280 95260
rect 267096 95208 267148 95260
rect 298376 95251 298428 95260
rect 298376 95217 298385 95251
rect 298385 95217 298419 95251
rect 298419 95217 298428 95251
rect 298376 95208 298428 95217
rect 353484 95251 353536 95260
rect 353484 95217 353493 95251
rect 353493 95217 353527 95251
rect 353527 95217 353536 95251
rect 353484 95208 353536 95217
rect 356612 95208 356664 95260
rect 408684 95251 408736 95260
rect 408684 95217 408693 95251
rect 408693 95217 408727 95251
rect 408727 95217 408736 95251
rect 408684 95208 408736 95217
rect 451556 95251 451608 95260
rect 451556 95217 451565 95251
rect 451565 95217 451599 95251
rect 451599 95217 451608 95251
rect 451556 95208 451608 95217
rect 265164 95183 265216 95192
rect 265164 95149 265173 95183
rect 265173 95149 265207 95183
rect 265207 95149 265216 95183
rect 265164 95140 265216 95149
rect 324504 95183 324556 95192
rect 324504 95149 324513 95183
rect 324513 95149 324547 95183
rect 324547 95149 324556 95183
rect 324504 95140 324556 95149
rect 327264 95183 327316 95192
rect 327264 95149 327273 95183
rect 327273 95149 327307 95183
rect 327307 95149 327316 95183
rect 327264 95140 327316 95149
rect 387984 95183 388036 95192
rect 387984 95149 387993 95183
rect 387993 95149 388027 95183
rect 388027 95149 388036 95183
rect 387984 95140 388036 95149
rect 393228 95183 393280 95192
rect 393228 95149 393237 95183
rect 393237 95149 393271 95183
rect 393271 95149 393280 95183
rect 393228 95140 393280 95149
rect 292672 93891 292724 93900
rect 292672 93857 292681 93891
rect 292681 93857 292715 93891
rect 292715 93857 292724 93891
rect 292672 93848 292724 93857
rect 334348 93891 334400 93900
rect 334348 93857 334357 93891
rect 334357 93857 334391 93891
rect 334391 93857 334400 93891
rect 334348 93848 334400 93857
rect 270960 92488 271012 92540
rect 233332 89700 233384 89752
rect 233516 89700 233568 89752
rect 298376 89743 298428 89752
rect 298376 89709 298385 89743
rect 298385 89709 298419 89743
rect 298419 89709 298428 89743
rect 298376 89700 298428 89709
rect 408684 89700 408736 89752
rect 422300 89700 422352 89752
rect 422484 89700 422536 89752
rect 427820 89700 427872 89752
rect 428004 89700 428056 89752
rect 230848 89675 230900 89684
rect 230848 89641 230857 89675
rect 230857 89641 230891 89675
rect 230891 89641 230900 89675
rect 230848 89632 230900 89641
rect 408776 89564 408828 89616
rect 241796 86955 241848 86964
rect 241796 86921 241805 86955
rect 241805 86921 241839 86955
rect 241839 86921 241848 86955
rect 241796 86912 241848 86921
rect 271972 86912 272024 86964
rect 272064 86912 272116 86964
rect 305184 86955 305236 86964
rect 305184 86921 305193 86955
rect 305193 86921 305227 86955
rect 305227 86921 305236 86955
rect 305184 86912 305236 86921
rect 308036 86955 308088 86964
rect 308036 86921 308045 86955
rect 308045 86921 308079 86955
rect 308079 86921 308088 86955
rect 308036 86912 308088 86921
rect 309324 86955 309376 86964
rect 309324 86921 309333 86955
rect 309333 86921 309367 86955
rect 309367 86921 309376 86955
rect 309324 86912 309376 86921
rect 310704 86955 310756 86964
rect 310704 86921 310713 86955
rect 310713 86921 310747 86955
rect 310747 86921 310756 86955
rect 310704 86912 310756 86921
rect 318984 86912 319036 86964
rect 342444 86955 342496 86964
rect 342444 86921 342453 86955
rect 342453 86921 342487 86955
rect 342487 86921 342496 86955
rect 342444 86912 342496 86921
rect 346584 86955 346636 86964
rect 346584 86921 346593 86955
rect 346593 86921 346627 86955
rect 346627 86921 346636 86955
rect 346584 86912 346636 86921
rect 352012 86912 352064 86964
rect 353484 86912 353536 86964
rect 353576 86912 353628 86964
rect 357624 86912 357676 86964
rect 357808 86912 357860 86964
rect 397644 86955 397696 86964
rect 397644 86921 397653 86955
rect 397653 86921 397687 86955
rect 397687 86921 397696 86955
rect 397644 86912 397696 86921
rect 400404 86912 400456 86964
rect 422392 86955 422444 86964
rect 422392 86921 422401 86955
rect 422401 86921 422435 86955
rect 422435 86921 422444 86955
rect 422392 86912 422444 86921
rect 427912 86955 427964 86964
rect 427912 86921 427921 86955
rect 427921 86921 427955 86955
rect 427955 86921 427964 86955
rect 427912 86912 427964 86921
rect 433524 86912 433576 86964
rect 243084 86844 243136 86896
rect 243268 86844 243320 86896
rect 252744 86887 252796 86896
rect 252744 86853 252753 86887
rect 252753 86853 252787 86887
rect 252787 86853 252796 86887
rect 252744 86844 252796 86853
rect 254124 86887 254176 86896
rect 254124 86853 254133 86887
rect 254133 86853 254167 86887
rect 254167 86853 254176 86887
rect 254124 86844 254176 86853
rect 259644 86887 259696 86896
rect 259644 86853 259653 86887
rect 259653 86853 259687 86887
rect 259687 86853 259696 86887
rect 259644 86844 259696 86853
rect 319076 86844 319128 86896
rect 331404 86887 331456 86896
rect 331404 86853 331413 86887
rect 331413 86853 331447 86887
rect 331447 86853 331456 86887
rect 331404 86844 331456 86853
rect 334348 86887 334400 86896
rect 334348 86853 334357 86887
rect 334357 86853 334391 86887
rect 334391 86853 334400 86887
rect 334348 86844 334400 86853
rect 352104 86844 352156 86896
rect 364524 86887 364576 86896
rect 364524 86853 364533 86887
rect 364533 86853 364567 86887
rect 364567 86853 364576 86887
rect 364524 86844 364576 86853
rect 370044 86887 370096 86896
rect 370044 86853 370053 86887
rect 370053 86853 370087 86887
rect 370087 86853 370096 86887
rect 370044 86844 370096 86853
rect 386604 86887 386656 86896
rect 386604 86853 386613 86887
rect 386613 86853 386647 86887
rect 386647 86853 386656 86887
rect 386604 86844 386656 86853
rect 392124 86887 392176 86896
rect 392124 86853 392133 86887
rect 392133 86853 392167 86887
rect 392167 86853 392176 86887
rect 392124 86844 392176 86853
rect 260748 85620 260800 85672
rect 261024 85552 261076 85604
rect 265164 85595 265216 85604
rect 265164 85561 265173 85595
rect 265173 85561 265207 85595
rect 265207 85561 265216 85595
rect 265164 85552 265216 85561
rect 298376 85595 298428 85604
rect 298376 85561 298385 85595
rect 298385 85561 298419 85595
rect 298419 85561 298428 85595
rect 298376 85552 298428 85561
rect 324504 85595 324556 85604
rect 324504 85561 324513 85595
rect 324513 85561 324547 85595
rect 324547 85561 324556 85595
rect 324504 85552 324556 85561
rect 327264 85595 327316 85604
rect 327264 85561 327273 85595
rect 327273 85561 327307 85595
rect 327307 85561 327316 85595
rect 327264 85552 327316 85561
rect 330024 85552 330076 85604
rect 330116 85552 330168 85604
rect 356428 85552 356480 85604
rect 356612 85552 356664 85604
rect 387984 85595 388036 85604
rect 387984 85561 387993 85595
rect 387993 85561 388027 85595
rect 388027 85561 388036 85595
rect 387984 85552 388036 85561
rect 393412 85552 393464 85604
rect 231952 85527 232004 85536
rect 231952 85493 231961 85527
rect 231961 85493 231995 85527
rect 231995 85493 232004 85527
rect 231952 85484 232004 85493
rect 236276 85527 236328 85536
rect 236276 85493 236285 85527
rect 236285 85493 236319 85527
rect 236319 85493 236328 85527
rect 236276 85484 236328 85493
rect 353484 85484 353536 85536
rect 451556 85484 451608 85536
rect 466552 85527 466604 85536
rect 466552 85493 466561 85527
rect 466561 85493 466595 85527
rect 466595 85493 466604 85527
rect 466552 85484 466604 85493
rect 353576 85416 353628 85468
rect 270960 82764 271012 82816
rect 359004 82807 359056 82816
rect 359004 82773 359013 82807
rect 359013 82773 359047 82807
rect 359047 82773 359056 82807
rect 359004 82764 359056 82773
rect 408776 82127 408828 82136
rect 408776 82093 408785 82127
rect 408785 82093 408819 82127
rect 408819 82093 408828 82127
rect 408776 82084 408828 82093
rect 298376 80724 298428 80776
rect 346492 80724 346544 80776
rect 472072 80767 472124 80776
rect 472072 80733 472081 80767
rect 472081 80733 472115 80767
rect 472115 80733 472124 80767
rect 472072 80724 472124 80733
rect 230940 80155 230992 80164
rect 230940 80121 230949 80155
rect 230949 80121 230983 80155
rect 230983 80121 230992 80155
rect 230940 80112 230992 80121
rect 244464 80044 244516 80096
rect 277492 80112 277544 80164
rect 294144 80112 294196 80164
rect 295524 80112 295576 80164
rect 295708 80112 295760 80164
rect 371424 80044 371476 80096
rect 376944 80044 376996 80096
rect 382464 80044 382516 80096
rect 277400 79976 277452 80028
rect 294144 79976 294196 80028
rect 244464 79908 244516 79960
rect 371424 79908 371476 79960
rect 376944 79908 376996 79960
rect 382464 79908 382516 79960
rect 2780 79840 2832 79892
rect 4804 79840 4856 79892
rect 281816 77324 281868 77376
rect 282000 77324 282052 77376
rect 230940 77299 230992 77308
rect 230940 77265 230949 77299
rect 230949 77265 230983 77299
rect 230983 77265 230992 77299
rect 230940 77256 230992 77265
rect 241796 77299 241848 77308
rect 241796 77265 241805 77299
rect 241805 77265 241839 77299
rect 241839 77265 241848 77299
rect 241796 77256 241848 77265
rect 252744 77299 252796 77308
rect 252744 77265 252753 77299
rect 252753 77265 252787 77299
rect 252787 77265 252796 77299
rect 252744 77256 252796 77265
rect 254124 77299 254176 77308
rect 254124 77265 254133 77299
rect 254133 77265 254167 77299
rect 254167 77265 254176 77299
rect 254124 77256 254176 77265
rect 259644 77299 259696 77308
rect 259644 77265 259653 77299
rect 259653 77265 259687 77299
rect 259687 77265 259696 77299
rect 259644 77256 259696 77265
rect 287152 77256 287204 77308
rect 287244 77256 287296 77308
rect 305184 77299 305236 77308
rect 305184 77265 305193 77299
rect 305193 77265 305227 77299
rect 305227 77265 305236 77299
rect 305184 77256 305236 77265
rect 308036 77299 308088 77308
rect 308036 77265 308045 77299
rect 308045 77265 308079 77299
rect 308079 77265 308088 77299
rect 308036 77256 308088 77265
rect 309324 77299 309376 77308
rect 309324 77265 309333 77299
rect 309333 77265 309367 77299
rect 309367 77265 309376 77299
rect 309324 77256 309376 77265
rect 310704 77299 310756 77308
rect 310704 77265 310713 77299
rect 310713 77265 310747 77299
rect 310747 77265 310756 77299
rect 310704 77256 310756 77265
rect 327264 77324 327316 77376
rect 347872 77324 347924 77376
rect 416780 77324 416832 77376
rect 416964 77324 417016 77376
rect 331404 77299 331456 77308
rect 331404 77265 331413 77299
rect 331413 77265 331447 77299
rect 331447 77265 331456 77299
rect 331404 77256 331456 77265
rect 334348 77299 334400 77308
rect 334348 77265 334357 77299
rect 334357 77265 334391 77299
rect 334391 77265 334400 77299
rect 334348 77256 334400 77265
rect 342444 77299 342496 77308
rect 342444 77265 342453 77299
rect 342453 77265 342487 77299
rect 342487 77265 342496 77299
rect 342444 77256 342496 77265
rect 364524 77299 364576 77308
rect 364524 77265 364533 77299
rect 364533 77265 364567 77299
rect 364567 77265 364576 77299
rect 364524 77256 364576 77265
rect 370044 77299 370096 77308
rect 370044 77265 370053 77299
rect 370053 77265 370087 77299
rect 370087 77265 370096 77299
rect 370044 77256 370096 77265
rect 381084 77256 381136 77308
rect 381176 77256 381228 77308
rect 386604 77299 386656 77308
rect 386604 77265 386613 77299
rect 386613 77265 386647 77299
rect 386647 77265 386656 77299
rect 386604 77256 386656 77265
rect 392124 77299 392176 77308
rect 392124 77265 392133 77299
rect 392133 77265 392167 77299
rect 392167 77265 392176 77299
rect 392124 77256 392176 77265
rect 397644 77299 397696 77308
rect 397644 77265 397653 77299
rect 397653 77265 397687 77299
rect 397687 77265 397696 77299
rect 397644 77256 397696 77265
rect 400312 77299 400364 77308
rect 400312 77265 400321 77299
rect 400321 77265 400355 77299
rect 400355 77265 400364 77299
rect 400312 77256 400364 77265
rect 408776 77299 408828 77308
rect 408776 77265 408785 77299
rect 408785 77265 408819 77299
rect 408819 77265 408828 77299
rect 408776 77256 408828 77265
rect 422484 77256 422536 77308
rect 428004 77256 428056 77308
rect 433432 77299 433484 77308
rect 433432 77265 433441 77299
rect 433441 77265 433475 77299
rect 433475 77265 433484 77299
rect 433432 77256 433484 77265
rect 277400 77231 277452 77240
rect 277400 77197 277409 77231
rect 277409 77197 277443 77231
rect 277443 77197 277452 77231
rect 277400 77188 277452 77197
rect 327172 77188 327224 77240
rect 347872 77188 347924 77240
rect 416964 77188 417016 77240
rect 330024 76032 330076 76084
rect 231952 75939 232004 75948
rect 231952 75905 231961 75939
rect 231961 75905 231995 75939
rect 231995 75905 232004 75939
rect 231952 75896 232004 75905
rect 236276 75939 236328 75948
rect 236276 75905 236285 75939
rect 236285 75905 236319 75939
rect 236319 75905 236328 75939
rect 236276 75896 236328 75905
rect 261024 75964 261076 76016
rect 330116 75896 330168 75948
rect 466644 75896 466696 75948
rect 230940 75871 230992 75880
rect 230940 75837 230949 75871
rect 230949 75837 230983 75871
rect 230983 75837 230992 75871
rect 230940 75828 230992 75837
rect 260840 75828 260892 75880
rect 327172 75871 327224 75880
rect 327172 75837 327181 75871
rect 327181 75837 327215 75871
rect 327215 75837 327224 75871
rect 327172 75828 327224 75837
rect 346492 75828 346544 75880
rect 346584 75828 346636 75880
rect 353576 75871 353628 75880
rect 353576 75837 353585 75871
rect 353585 75837 353619 75871
rect 353619 75837 353628 75871
rect 353576 75828 353628 75837
rect 387984 75828 388036 75880
rect 388168 75828 388220 75880
rect 267096 74536 267148 74588
rect 267280 74536 267332 74588
rect 357624 74468 357676 74520
rect 359004 73219 359056 73228
rect 359004 73185 359013 73219
rect 359013 73185 359047 73219
rect 359047 73185 359056 73219
rect 359004 73176 359056 73185
rect 272064 73108 272116 73160
rect 281816 72428 281868 72480
rect 282000 72428 282052 72480
rect 240232 70456 240284 70508
rect 243084 70388 243136 70440
rect 236276 70363 236328 70372
rect 236276 70329 236285 70363
rect 236285 70329 236319 70363
rect 236319 70329 236328 70363
rect 236276 70320 236328 70329
rect 240232 70320 240284 70372
rect 266544 70456 266596 70508
rect 408776 70431 408828 70440
rect 408776 70397 408785 70431
rect 408785 70397 408819 70431
rect 408819 70397 408828 70431
rect 408776 70388 408828 70397
rect 266452 70320 266504 70372
rect 277492 70320 277544 70372
rect 243176 70252 243228 70304
rect 292764 69028 292816 69080
rect 292764 68892 292816 68944
rect 231860 67600 231912 67652
rect 231952 67600 232004 67652
rect 236276 67643 236328 67652
rect 236276 67609 236285 67643
rect 236285 67609 236319 67643
rect 236319 67609 236328 67643
rect 236276 67600 236328 67609
rect 267280 67668 267332 67720
rect 386604 67668 386656 67720
rect 392124 67668 392176 67720
rect 298376 67600 298428 67652
rect 319076 67643 319128 67652
rect 319076 67609 319085 67643
rect 319085 67609 319119 67643
rect 319119 67609 319128 67643
rect 319076 67600 319128 67609
rect 324412 67600 324464 67652
rect 324504 67600 324556 67652
rect 347872 67600 347924 67652
rect 348056 67600 348108 67652
rect 386696 67600 386748 67652
rect 392216 67600 392268 67652
rect 408776 67643 408828 67652
rect 408776 67609 408785 67643
rect 408785 67609 408819 67643
rect 408819 67609 408828 67643
rect 408776 67600 408828 67609
rect 416872 67643 416924 67652
rect 416872 67609 416881 67643
rect 416881 67609 416915 67643
rect 416915 67609 416924 67643
rect 416872 67600 416924 67609
rect 433432 67600 433484 67652
rect 433524 67600 433576 67652
rect 451464 67643 451516 67652
rect 451464 67609 451473 67643
rect 451473 67609 451507 67643
rect 451507 67609 451516 67643
rect 451464 67600 451516 67609
rect 472072 67643 472124 67652
rect 472072 67609 472081 67643
rect 472081 67609 472115 67643
rect 472115 67609 472124 67643
rect 472072 67600 472124 67609
rect 267188 67532 267240 67584
rect 305184 67532 305236 67584
rect 305276 67532 305328 67584
rect 308036 67575 308088 67584
rect 308036 67541 308045 67575
rect 308045 67541 308079 67575
rect 308079 67541 308088 67575
rect 308036 67532 308088 67541
rect 356520 67532 356572 67584
rect 393228 67575 393280 67584
rect 393228 67541 393237 67575
rect 393237 67541 393271 67575
rect 393271 67541 393280 67575
rect 393228 67532 393280 67541
rect 397644 67575 397696 67584
rect 397644 67541 397653 67575
rect 397653 67541 397687 67575
rect 397687 67541 397696 67575
rect 397644 67532 397696 67541
rect 260840 66308 260892 66360
rect 261024 66308 261076 66360
rect 231032 66240 231084 66292
rect 319076 66283 319128 66292
rect 319076 66249 319085 66283
rect 319085 66249 319119 66283
rect 319119 66249 319128 66283
rect 319076 66240 319128 66249
rect 327264 66240 327316 66292
rect 330024 66283 330076 66292
rect 330024 66249 330033 66283
rect 330033 66249 330067 66283
rect 330067 66249 330076 66283
rect 330024 66240 330076 66249
rect 353668 66240 353720 66292
rect 236276 66172 236328 66224
rect 281724 66215 281776 66224
rect 281724 66181 281733 66215
rect 281733 66181 281767 66215
rect 281767 66181 281776 66215
rect 281724 66172 281776 66181
rect 309416 66172 309468 66224
rect 336832 66172 336884 66224
rect 336924 66172 336976 66224
rect 387984 66215 388036 66224
rect 387984 66181 387993 66215
rect 387993 66181 388027 66215
rect 388027 66181 388036 66215
rect 387984 66172 388036 66181
rect 451464 66215 451516 66224
rect 451464 66181 451473 66215
rect 451473 66181 451507 66215
rect 451507 66181 451516 66215
rect 451464 66172 451516 66181
rect 466460 66215 466512 66224
rect 466460 66181 466469 66215
rect 466469 66181 466503 66215
rect 466503 66181 466512 66215
rect 466460 66172 466512 66181
rect 330024 64991 330076 65000
rect 330024 64957 330033 64991
rect 330033 64957 330067 64991
rect 330067 64957 330076 64991
rect 330024 64948 330076 64957
rect 270684 64923 270736 64932
rect 270684 64889 270693 64923
rect 270693 64889 270727 64923
rect 270727 64889 270736 64923
rect 270684 64880 270736 64889
rect 357532 64923 357584 64932
rect 357532 64889 357541 64923
rect 357541 64889 357575 64923
rect 357575 64889 357584 64923
rect 357532 64880 357584 64889
rect 243176 64812 243228 64864
rect 261024 64812 261076 64864
rect 292488 64812 292540 64864
rect 292764 64812 292816 64864
rect 332784 64812 332836 64864
rect 332876 64812 332928 64864
rect 529480 64812 529532 64864
rect 580172 64812 580224 64864
rect 271972 63563 272024 63572
rect 271972 63529 271981 63563
rect 271981 63529 272015 63563
rect 272015 63529 272024 63563
rect 271972 63520 272024 63529
rect 330024 63452 330076 63504
rect 332876 63495 332928 63504
rect 332876 63461 332885 63495
rect 332885 63461 332919 63495
rect 332919 63461 332928 63495
rect 332876 63452 332928 63461
rect 359096 63495 359148 63504
rect 359096 63461 359105 63495
rect 359105 63461 359139 63495
rect 359139 63461 359148 63495
rect 359096 63452 359148 63461
rect 408776 62815 408828 62824
rect 408776 62781 408785 62815
rect 408785 62781 408819 62815
rect 408819 62781 408828 62815
rect 408776 62772 408828 62781
rect 392216 61684 392268 61736
rect 392400 61684 392452 61736
rect 370044 61115 370096 61124
rect 370044 61081 370053 61115
rect 370053 61081 370087 61115
rect 370087 61081 370096 61115
rect 370044 61072 370096 61081
rect 375564 61115 375616 61124
rect 375564 61081 375573 61115
rect 375573 61081 375607 61115
rect 375607 61081 375616 61115
rect 375564 61072 375616 61081
rect 416780 60664 416832 60716
rect 416964 60664 417016 60716
rect 433524 60664 433576 60716
rect 433708 60664 433760 60716
rect 451648 60664 451700 60716
rect 471980 60664 472032 60716
rect 472164 60664 472216 60716
rect 371424 60639 371476 60648
rect 371424 60605 371433 60639
rect 371433 60605 371467 60639
rect 371467 60605 371476 60639
rect 371424 60596 371476 60605
rect 318984 60027 319036 60036
rect 318984 59993 318993 60027
rect 318993 59993 319027 60027
rect 319027 59993 319036 60027
rect 318984 59984 319036 59993
rect 259644 59755 259696 59764
rect 259644 59721 259653 59755
rect 259653 59721 259687 59755
rect 259687 59721 259696 59755
rect 259644 59712 259696 59721
rect 271972 58599 272024 58608
rect 271972 58565 271981 58599
rect 271981 58565 272015 58599
rect 272015 58565 272024 58599
rect 271972 58556 272024 58565
rect 352012 58123 352064 58132
rect 352012 58089 352021 58123
rect 352021 58089 352055 58123
rect 352055 58089 352064 58123
rect 352012 58080 352064 58089
rect 266452 57944 266504 57996
rect 266544 57944 266596 57996
rect 267096 57944 267148 57996
rect 267188 57944 267240 57996
rect 293960 57944 294012 57996
rect 294144 57944 294196 57996
rect 295524 57944 295576 57996
rect 308036 57987 308088 57996
rect 308036 57953 308045 57987
rect 308045 57953 308079 57987
rect 308079 57953 308088 57987
rect 308036 57944 308088 57953
rect 347964 57944 348016 57996
rect 348056 57944 348108 57996
rect 356428 57987 356480 57996
rect 356428 57953 356437 57987
rect 356437 57953 356471 57987
rect 356471 57953 356480 57987
rect 356428 57944 356480 57953
rect 386604 57944 386656 57996
rect 386696 57944 386748 57996
rect 393228 57987 393280 57996
rect 393228 57953 393237 57987
rect 393237 57953 393271 57987
rect 393271 57953 393280 57987
rect 393228 57944 393280 57953
rect 397736 57944 397788 57996
rect 408776 57987 408828 57996
rect 408776 57953 408785 57987
rect 408785 57953 408819 57987
rect 408819 57953 408828 57987
rect 408776 57944 408828 57953
rect 277584 57876 277636 57928
rect 288624 57876 288676 57928
rect 277676 57808 277728 57860
rect 324412 57919 324464 57928
rect 324412 57885 324421 57919
rect 324421 57885 324455 57919
rect 324455 57885 324464 57919
rect 324412 57876 324464 57885
rect 376944 57876 376996 57928
rect 377036 57876 377088 57928
rect 382464 57876 382516 57928
rect 416964 57876 417016 57928
rect 433708 57876 433760 57928
rect 472164 57876 472216 57928
rect 295616 57808 295668 57860
rect 270684 57536 270736 57588
rect 371424 56695 371476 56704
rect 371424 56661 371433 56695
rect 371433 56661 371467 56695
rect 371467 56661 371476 56695
rect 371424 56652 371476 56661
rect 281724 56627 281776 56636
rect 281724 56593 281733 56627
rect 281733 56593 281767 56627
rect 281767 56593 281776 56627
rect 281724 56584 281776 56593
rect 388076 56584 388128 56636
rect 466828 56584 466880 56636
rect 244464 56516 244516 56568
rect 249984 56559 250036 56568
rect 249984 56525 249993 56559
rect 249993 56525 250027 56559
rect 250027 56525 250036 56559
rect 249984 56516 250036 56525
rect 255504 56516 255556 56568
rect 277492 56516 277544 56568
rect 277676 56516 277728 56568
rect 283104 56516 283156 56568
rect 298284 56559 298336 56568
rect 298284 56525 298293 56559
rect 298293 56525 298327 56559
rect 298327 56525 298336 56559
rect 298284 56516 298336 56525
rect 336924 56559 336976 56568
rect 336924 56525 336933 56559
rect 336933 56525 336967 56559
rect 336967 56525 336976 56559
rect 336924 56516 336976 56525
rect 371424 56559 371476 56568
rect 371424 56525 371433 56559
rect 371433 56525 371467 56559
rect 371467 56525 371476 56559
rect 371424 56516 371476 56525
rect 392308 56516 392360 56568
rect 451648 56559 451700 56568
rect 451648 56525 451657 56559
rect 451657 56525 451691 56559
rect 451691 56525 451700 56559
rect 451648 56516 451700 56525
rect 331404 55675 331456 55684
rect 331404 55641 331413 55675
rect 331413 55641 331447 55675
rect 331447 55641 331456 55675
rect 331404 55632 331456 55641
rect 334348 55675 334400 55684
rect 334348 55641 334357 55675
rect 334357 55641 334391 55675
rect 334391 55641 334400 55675
rect 334348 55632 334400 55641
rect 242992 55267 243044 55276
rect 242992 55233 243001 55267
rect 243001 55233 243035 55267
rect 243035 55233 243044 55267
rect 242992 55224 243044 55233
rect 260840 55267 260892 55276
rect 260840 55233 260849 55267
rect 260849 55233 260883 55267
rect 260883 55233 260892 55267
rect 260840 55224 260892 55233
rect 292764 55199 292816 55208
rect 292764 55165 292773 55199
rect 292773 55165 292807 55199
rect 292807 55165 292816 55199
rect 292764 55156 292816 55165
rect 332876 55199 332928 55208
rect 332876 55165 332885 55199
rect 332885 55165 332919 55199
rect 332919 55165 332928 55199
rect 332876 55156 332928 55165
rect 329932 53839 329984 53848
rect 329932 53805 329941 53839
rect 329941 53805 329975 53839
rect 329975 53805 329984 53839
rect 329932 53796 329984 53805
rect 352012 53839 352064 53848
rect 352012 53805 352021 53839
rect 352021 53805 352055 53839
rect 352055 53805 352064 53839
rect 352012 53796 352064 53805
rect 359188 53796 359240 53848
rect 400496 51144 400548 51196
rect 408776 51187 408828 51196
rect 408776 51153 408785 51187
rect 408785 51153 408819 51187
rect 408819 51153 408828 51187
rect 408776 51144 408828 51153
rect 342444 51076 342496 51128
rect 342444 50940 342496 50992
rect 254124 48356 254176 48408
rect 309416 48399 309468 48408
rect 309416 48365 309425 48399
rect 309425 48365 309459 48399
rect 309459 48365 309468 48399
rect 309416 48356 309468 48365
rect 327264 48356 327316 48408
rect 400404 48399 400456 48408
rect 400404 48365 400413 48399
rect 400413 48365 400447 48399
rect 400447 48365 400456 48399
rect 400404 48356 400456 48365
rect 408684 48356 408736 48408
rect 416872 48399 416924 48408
rect 416872 48365 416881 48399
rect 416881 48365 416915 48399
rect 416915 48365 416924 48399
rect 416872 48356 416924 48365
rect 254216 48288 254268 48340
rect 259736 48288 259788 48340
rect 265164 48288 265216 48340
rect 265348 48288 265400 48340
rect 281724 48288 281776 48340
rect 281816 48288 281868 48340
rect 288532 48331 288584 48340
rect 288532 48297 288541 48331
rect 288541 48297 288575 48331
rect 288575 48297 288584 48331
rect 288532 48288 288584 48297
rect 327172 48288 327224 48340
rect 331496 48288 331548 48340
rect 334440 48288 334492 48340
rect 370136 48288 370188 48340
rect 375656 48288 375708 48340
rect 382372 48331 382424 48340
rect 382372 48297 382381 48331
rect 382381 48297 382415 48331
rect 382415 48297 382424 48331
rect 382372 48288 382424 48297
rect 386604 48288 386656 48340
rect 386696 48288 386748 48340
rect 387892 48288 387944 48340
rect 388076 48288 388128 48340
rect 422392 48288 422444 48340
rect 422484 48288 422536 48340
rect 433616 48331 433668 48340
rect 433616 48297 433625 48331
rect 433625 48297 433659 48331
rect 433659 48297 433668 48331
rect 433616 48288 433668 48297
rect 466644 48288 466696 48340
rect 466828 48288 466880 48340
rect 472072 48331 472124 48340
rect 472072 48297 472081 48331
rect 472081 48297 472115 48331
rect 472115 48297 472124 48331
rect 472072 48288 472124 48297
rect 295616 48220 295668 48272
rect 295708 48220 295760 48272
rect 308128 48263 308180 48272
rect 308128 48229 308137 48263
rect 308137 48229 308171 48263
rect 308171 48229 308180 48263
rect 308128 48220 308180 48229
rect 381176 48220 381228 48272
rect 381268 48220 381320 48272
rect 400404 48220 400456 48272
rect 400772 48220 400824 48272
rect 416872 48220 416924 48272
rect 417056 48220 417108 48272
rect 236276 46996 236328 47048
rect 282920 47039 282972 47048
rect 282920 47005 282929 47039
rect 282929 47005 282963 47039
rect 282963 47005 282972 47039
rect 282920 46996 282972 47005
rect 371332 46996 371384 47048
rect 392124 47039 392176 47048
rect 392124 47005 392133 47039
rect 392133 47005 392167 47039
rect 392167 47005 392176 47039
rect 392124 46996 392176 47005
rect 244372 46971 244424 46980
rect 244372 46937 244381 46971
rect 244381 46937 244415 46971
rect 244415 46937 244424 46971
rect 244372 46928 244424 46937
rect 249984 46971 250036 46980
rect 249984 46937 249993 46971
rect 249993 46937 250027 46971
rect 250027 46937 250036 46971
rect 249984 46928 250036 46937
rect 255412 46971 255464 46980
rect 255412 46937 255421 46971
rect 255421 46937 255455 46971
rect 255455 46937 255464 46971
rect 255412 46928 255464 46937
rect 270592 46971 270644 46980
rect 270592 46937 270601 46971
rect 270601 46937 270635 46971
rect 270635 46937 270644 46971
rect 270592 46928 270644 46937
rect 298376 46928 298428 46980
rect 318984 46971 319036 46980
rect 318984 46937 318993 46971
rect 318993 46937 319027 46971
rect 319027 46937 319036 46971
rect 318984 46928 319036 46937
rect 332876 46928 332928 46980
rect 336924 46971 336976 46980
rect 336924 46937 336933 46971
rect 336933 46937 336967 46971
rect 336967 46937 336976 46971
rect 336924 46928 336976 46937
rect 451832 46928 451884 46980
rect 231860 46860 231912 46912
rect 232044 46860 232096 46912
rect 236276 46860 236328 46912
rect 236460 46860 236512 46912
rect 243176 46860 243228 46912
rect 243268 46860 243320 46912
rect 267004 46860 267056 46912
rect 267188 46860 267240 46912
rect 282920 46860 282972 46912
rect 283104 46860 283156 46912
rect 310612 46860 310664 46912
rect 342444 46903 342496 46912
rect 342444 46869 342453 46903
rect 342453 46869 342487 46903
rect 342487 46869 342496 46903
rect 342444 46860 342496 46869
rect 359004 46860 359056 46912
rect 359188 46860 359240 46912
rect 371332 46860 371384 46912
rect 387892 46903 387944 46912
rect 387892 46869 387901 46903
rect 387901 46869 387935 46903
rect 387935 46869 387944 46903
rect 387892 46860 387944 46869
rect 392124 46860 392176 46912
rect 408776 46903 408828 46912
rect 408776 46869 408785 46903
rect 408785 46869 408819 46903
rect 408819 46869 408828 46903
rect 408776 46860 408828 46869
rect 332876 46792 332928 46844
rect 371516 46792 371568 46844
rect 392124 46724 392176 46776
rect 272064 45568 272116 45620
rect 292948 45568 293000 45620
rect 324504 45611 324556 45620
rect 324504 45577 324513 45611
rect 324513 45577 324547 45611
rect 324547 45577 324556 45611
rect 324504 45568 324556 45577
rect 243268 45500 243320 45552
rect 267188 45500 267240 45552
rect 277584 45543 277636 45552
rect 277584 45509 277593 45543
rect 277593 45509 277627 45543
rect 277627 45509 277636 45543
rect 277584 45500 277636 45509
rect 283104 45500 283156 45552
rect 332876 45500 332928 45552
rect 352012 45500 352064 45552
rect 352380 45500 352432 45552
rect 359004 45543 359056 45552
rect 359004 45509 359013 45543
rect 359013 45509 359047 45543
rect 359047 45509 359056 45543
rect 359004 45500 359056 45509
rect 255412 44820 255464 44872
rect 230664 43460 230716 43512
rect 230848 43460 230900 43512
rect 298376 42075 298428 42084
rect 298376 42041 298385 42075
rect 298385 42041 298419 42075
rect 298419 42041 298428 42075
rect 298376 42032 298428 42041
rect 309416 42032 309468 42084
rect 375656 41556 375708 41608
rect 370136 41420 370188 41472
rect 310612 41352 310664 41404
rect 471980 41352 472032 41404
rect 472164 41352 472216 41404
rect 433616 41327 433668 41336
rect 433616 41293 433625 41327
rect 433625 41293 433659 41327
rect 433659 41293 433668 41327
rect 433616 41284 433668 41293
rect 397644 40332 397696 40384
rect 405648 40332 405700 40384
rect 475936 40196 475988 40248
rect 478236 40196 478288 40248
rect 514576 40196 514628 40248
rect 514852 40196 514904 40248
rect 540980 40060 541032 40112
rect 545856 40060 545908 40112
rect 302148 39992 302200 40044
rect 307300 39992 307352 40044
rect 272064 38743 272116 38752
rect 272064 38709 272073 38743
rect 272073 38709 272107 38743
rect 272107 38709 272116 38743
rect 272064 38700 272116 38709
rect 382372 38700 382424 38752
rect 281632 38632 281684 38684
rect 281816 38632 281868 38684
rect 308128 38675 308180 38684
rect 308128 38641 308137 38675
rect 308137 38641 308171 38675
rect 308171 38641 308180 38675
rect 308128 38632 308180 38641
rect 376944 38632 376996 38684
rect 377036 38632 377088 38684
rect 294144 38607 294196 38616
rect 294144 38573 294153 38607
rect 294153 38573 294187 38607
rect 294187 38573 294196 38607
rect 294144 38564 294196 38573
rect 369952 38607 370004 38616
rect 369952 38573 369961 38607
rect 369961 38573 369995 38607
rect 369995 38573 370004 38607
rect 369952 38564 370004 38573
rect 382372 38564 382424 38616
rect 416964 38564 417016 38616
rect 422484 38607 422536 38616
rect 422484 38573 422493 38607
rect 422493 38573 422527 38607
rect 422527 38573 422536 38607
rect 422484 38564 422536 38573
rect 472164 38564 472216 38616
rect 408868 38496 408920 38548
rect 295708 38292 295760 38344
rect 295708 38156 295760 38208
rect 252744 37383 252796 37392
rect 252744 37349 252753 37383
rect 252753 37349 252787 37383
rect 252787 37349 252796 37383
rect 252744 37340 252796 37349
rect 331496 37340 331548 37392
rect 334440 37340 334492 37392
rect 386696 37340 386748 37392
rect 433524 37340 433576 37392
rect 331404 37272 331456 37324
rect 334348 37272 334400 37324
rect 342536 37272 342588 37324
rect 375472 37315 375524 37324
rect 375472 37281 375481 37315
rect 375481 37281 375515 37315
rect 375515 37281 375524 37315
rect 375472 37272 375524 37281
rect 386788 37272 386840 37324
rect 387892 37315 387944 37324
rect 387892 37281 387901 37315
rect 387901 37281 387935 37315
rect 387935 37281 387944 37315
rect 387892 37272 387944 37281
rect 230664 37204 230716 37256
rect 230756 37204 230808 37256
rect 272064 37247 272116 37256
rect 272064 37213 272073 37247
rect 272073 37213 272107 37247
rect 272107 37213 272116 37247
rect 272064 37204 272116 37213
rect 433616 37247 433668 37256
rect 433616 37213 433625 37247
rect 433625 37213 433659 37247
rect 433659 37213 433668 37247
rect 433616 37204 433668 37213
rect 292948 37136 293000 37188
rect 242992 35955 243044 35964
rect 242992 35921 243001 35955
rect 243001 35921 243035 35955
rect 243035 35921 243044 35955
rect 242992 35912 243044 35921
rect 267004 35955 267056 35964
rect 267004 35921 267013 35955
rect 267013 35921 267047 35955
rect 267047 35921 267056 35955
rect 267004 35912 267056 35921
rect 277584 35955 277636 35964
rect 277584 35921 277593 35955
rect 277593 35921 277627 35955
rect 277627 35921 277636 35955
rect 277584 35912 277636 35921
rect 292764 35955 292816 35964
rect 292764 35921 292773 35955
rect 292773 35921 292807 35955
rect 292807 35921 292816 35955
rect 292764 35912 292816 35921
rect 332692 35955 332744 35964
rect 332692 35921 332701 35955
rect 332701 35921 332735 35955
rect 332735 35921 332744 35955
rect 332692 35912 332744 35921
rect 359004 35955 359056 35964
rect 359004 35921 359013 35955
rect 359013 35921 359047 35955
rect 359047 35921 359056 35955
rect 359004 35912 359056 35921
rect 3424 35844 3476 35896
rect 72424 35844 72476 35896
rect 334348 35887 334400 35896
rect 334348 35853 334357 35887
rect 334357 35853 334391 35887
rect 334391 35853 334400 35887
rect 334348 35844 334400 35853
rect 369952 33804 370004 33856
rect 370228 33804 370280 33856
rect 298192 32376 298244 32428
rect 319076 31764 319128 31816
rect 233332 31696 233384 31748
rect 233516 31696 233568 31748
rect 281632 31696 281684 31748
rect 281816 31696 281868 31748
rect 346584 31764 346636 31816
rect 400680 31807 400732 31816
rect 400680 31773 400689 31807
rect 400689 31773 400723 31807
rect 400723 31773 400732 31807
rect 400680 31764 400732 31773
rect 427912 31764 427964 31816
rect 346492 31696 346544 31748
rect 427820 31696 427872 31748
rect 451648 31696 451700 31748
rect 451832 31696 451884 31748
rect 319076 31628 319128 31680
rect 270684 29044 270736 29096
rect 294144 29087 294196 29096
rect 294144 29053 294153 29087
rect 294153 29053 294187 29087
rect 294187 29053 294196 29087
rect 294144 29044 294196 29053
rect 400680 29087 400732 29096
rect 400680 29053 400689 29087
rect 400689 29053 400723 29087
rect 400723 29053 400732 29087
rect 400680 29044 400732 29053
rect 236276 28976 236328 29028
rect 236368 28976 236420 29028
rect 252836 28976 252888 29028
rect 270776 28976 270828 29028
rect 309324 29019 309376 29028
rect 309324 28985 309333 29019
rect 309333 28985 309367 29019
rect 309367 28985 309376 29019
rect 309324 28976 309376 28985
rect 381176 28976 381228 29028
rect 381268 28976 381320 29028
rect 386696 28976 386748 29028
rect 416872 29019 416924 29028
rect 231860 28908 231912 28960
rect 232044 28908 232096 28960
rect 244464 28908 244516 28960
rect 244556 28908 244608 28960
rect 254032 28908 254084 28960
rect 254216 28908 254268 28960
rect 259736 28908 259788 28960
rect 259828 28908 259880 28960
rect 265164 28908 265216 28960
rect 265256 28908 265308 28960
rect 266360 28908 266412 28960
rect 266544 28908 266596 28960
rect 292764 28908 292816 28960
rect 292856 28908 292908 28960
rect 293960 28908 294012 28960
rect 294144 28908 294196 28960
rect 295524 28908 295576 28960
rect 295616 28908 295668 28960
rect 308128 28908 308180 28960
rect 348056 28908 348108 28960
rect 348148 28908 348200 28960
rect 353576 28908 353628 28960
rect 353668 28908 353720 28960
rect 356428 28908 356480 28960
rect 356520 28908 356572 28960
rect 416872 28985 416881 29019
rect 416881 28985 416915 29019
rect 416915 28985 416924 29019
rect 416872 28976 416924 28985
rect 466552 28976 466604 29028
rect 466644 28976 466696 29028
rect 472072 29019 472124 29028
rect 472072 28985 472081 29019
rect 472081 28985 472115 29019
rect 472115 28985 472124 29019
rect 472072 28976 472124 28985
rect 392032 28908 392084 28960
rect 392216 28908 392268 28960
rect 393228 28951 393280 28960
rect 393228 28917 393237 28951
rect 393237 28917 393271 28951
rect 393271 28917 393280 28951
rect 393228 28908 393280 28917
rect 451832 28908 451884 28960
rect 386788 28840 386840 28892
rect 387892 27752 387944 27804
rect 277584 27684 277636 27736
rect 277676 27684 277728 27736
rect 282920 27659 282972 27668
rect 282920 27625 282929 27659
rect 282929 27625 282963 27659
rect 282963 27625 282972 27659
rect 282920 27616 282972 27625
rect 327172 27616 327224 27668
rect 327264 27616 327316 27668
rect 387800 27659 387852 27668
rect 387800 27625 387809 27659
rect 387809 27625 387843 27659
rect 387843 27625 387852 27659
rect 387800 27616 387852 27625
rect 422392 27616 422444 27668
rect 433708 27616 433760 27668
rect 230756 27548 230808 27600
rect 230848 27548 230900 27600
rect 252836 27591 252888 27600
rect 252836 27557 252845 27591
rect 252845 27557 252879 27591
rect 252879 27557 252888 27591
rect 252836 27548 252888 27557
rect 255320 27548 255372 27600
rect 259828 27591 259880 27600
rect 259828 27557 259837 27591
rect 259837 27557 259871 27591
rect 259871 27557 259880 27591
rect 259828 27548 259880 27557
rect 267004 27548 267056 27600
rect 267096 27548 267148 27600
rect 272064 27548 272116 27600
rect 293960 27591 294012 27600
rect 293960 27557 293969 27591
rect 293969 27557 294003 27591
rect 294003 27557 294012 27591
rect 293960 27548 294012 27557
rect 321652 27591 321704 27600
rect 321652 27557 321661 27591
rect 321661 27557 321695 27591
rect 321695 27557 321704 27591
rect 321652 27548 321704 27557
rect 336924 27548 336976 27600
rect 346492 27548 346544 27600
rect 353668 27591 353720 27600
rect 353668 27557 353677 27591
rect 353677 27557 353711 27591
rect 353711 27557 353720 27591
rect 353668 27548 353720 27557
rect 359004 27591 359056 27600
rect 359004 27557 359013 27591
rect 359013 27557 359047 27591
rect 359047 27557 359056 27591
rect 359004 27548 359056 27557
rect 400588 27591 400640 27600
rect 400588 27557 400597 27591
rect 400597 27557 400631 27591
rect 400631 27557 400640 27591
rect 400588 27548 400640 27557
rect 324504 26324 324556 26376
rect 324412 26256 324464 26308
rect 334532 26256 334584 26308
rect 230756 26188 230808 26240
rect 277584 26188 277636 26240
rect 334348 26120 334400 26172
rect 334532 26120 334584 26172
rect 346492 22720 346544 22772
rect 348148 22720 348200 22772
rect 270776 22584 270828 22636
rect 305276 22176 305328 22228
rect 281816 22108 281868 22160
rect 364524 22108 364576 22160
rect 281724 22040 281776 22092
rect 408776 22108 408828 22160
rect 408684 22040 408736 22092
rect 416780 22040 416832 22092
rect 416964 22040 417016 22092
rect 364524 21972 364576 22024
rect 236276 19320 236328 19372
rect 260932 19320 260984 19372
rect 261024 19320 261076 19372
rect 282920 19320 282972 19372
rect 283196 19320 283248 19372
rect 288440 19320 288492 19372
rect 288624 19320 288676 19372
rect 305092 19363 305144 19372
rect 305092 19329 305101 19363
rect 305101 19329 305135 19363
rect 305135 19329 305144 19363
rect 305092 19320 305144 19329
rect 308036 19363 308088 19372
rect 308036 19329 308045 19363
rect 308045 19329 308079 19363
rect 308079 19329 308088 19363
rect 308036 19320 308088 19329
rect 310428 19320 310480 19372
rect 310704 19320 310756 19372
rect 324412 19320 324464 19372
rect 324504 19320 324556 19372
rect 352012 19320 352064 19372
rect 352196 19320 352248 19372
rect 357532 19320 357584 19372
rect 357624 19320 357676 19372
rect 370044 19320 370096 19372
rect 370228 19320 370280 19372
rect 371332 19320 371384 19372
rect 371516 19320 371568 19372
rect 375564 19320 375616 19372
rect 375748 19320 375800 19372
rect 381084 19320 381136 19372
rect 381268 19320 381320 19372
rect 382280 19320 382332 19372
rect 382464 19320 382516 19372
rect 393228 19363 393280 19372
rect 393228 19329 393237 19363
rect 393237 19329 393271 19363
rect 393271 19329 393280 19363
rect 393228 19320 393280 19329
rect 451740 19363 451792 19372
rect 451740 19329 451749 19363
rect 451749 19329 451783 19363
rect 451783 19329 451792 19363
rect 451740 19320 451792 19329
rect 231860 19252 231912 19304
rect 233332 19252 233384 19304
rect 233424 19252 233476 19304
rect 231952 19184 232004 19236
rect 353668 19295 353720 19304
rect 353668 19261 353677 19295
rect 353677 19261 353711 19295
rect 353711 19261 353720 19295
rect 353668 19252 353720 19261
rect 416964 19295 417016 19304
rect 416964 19261 416973 19295
rect 416973 19261 417007 19295
rect 417007 19261 417016 19295
rect 416964 19252 417016 19261
rect 236368 19184 236420 19236
rect 422116 19184 422168 19236
rect 422484 19184 422536 19236
rect 386788 18980 386840 19032
rect 386788 18844 386840 18896
rect 252836 18003 252888 18012
rect 252836 17969 252845 18003
rect 252845 17969 252879 18003
rect 252879 17969 252888 18003
rect 252836 17960 252888 17969
rect 259828 18003 259880 18012
rect 259828 17969 259837 18003
rect 259837 17969 259871 18003
rect 259871 17969 259880 18003
rect 259828 17960 259880 17969
rect 271972 18003 272024 18012
rect 271972 17969 271981 18003
rect 271981 17969 272015 18003
rect 272015 17969 272024 18003
rect 271972 17960 272024 17969
rect 293960 18003 294012 18012
rect 293960 17969 293969 18003
rect 293969 17969 294003 18003
rect 294003 17969 294012 18003
rect 293960 17960 294012 17969
rect 321744 17960 321796 18012
rect 336832 18003 336884 18012
rect 336832 17969 336841 18003
rect 336841 17969 336875 18003
rect 336875 17969 336884 18003
rect 336832 17960 336884 17969
rect 359004 18003 359056 18012
rect 359004 17969 359013 18003
rect 359013 17969 359047 18003
rect 359047 17969 359056 18003
rect 359004 17960 359056 17969
rect 400588 18003 400640 18012
rect 400588 17969 400597 18003
rect 400597 17969 400631 18003
rect 400631 17969 400640 18003
rect 400588 17960 400640 17969
rect 381084 17892 381136 17944
rect 382464 17892 382516 17944
rect 400588 17824 400640 17876
rect 278780 16872 278832 16924
rect 288348 16872 288400 16924
rect 408408 16804 408460 16856
rect 410708 16804 410760 16856
rect 475936 16804 475988 16856
rect 477500 16804 477552 16856
rect 347688 16668 347740 16720
rect 355968 16668 356020 16720
rect 521660 16668 521712 16720
rect 524512 16668 524564 16720
rect 277492 16643 277544 16652
rect 277492 16609 277501 16643
rect 277501 16609 277535 16643
rect 277535 16609 277544 16643
rect 277492 16600 277544 16609
rect 125416 16328 125468 16380
rect 292764 16328 292816 16380
rect 121368 16260 121420 16312
rect 291292 16260 291344 16312
rect 114468 16192 114520 16244
rect 287244 16192 287296 16244
rect 110328 16124 110380 16176
rect 285772 16124 285824 16176
rect 107568 16056 107620 16108
rect 284392 16056 284444 16108
rect 103428 15988 103480 16040
rect 281724 15988 281776 16040
rect 28908 15920 28960 15972
rect 243084 15920 243136 15972
rect 31668 15852 31720 15904
rect 245752 15852 245804 15904
rect 129648 15104 129700 15156
rect 295524 15104 295576 15156
rect 99288 15036 99340 15088
rect 280252 15036 280304 15088
rect 96528 14968 96580 15020
rect 278872 14968 278924 15020
rect 92388 14900 92440 14952
rect 276112 14900 276164 14952
rect 89628 14832 89680 14884
rect 274732 14832 274784 14884
rect 85488 14764 85540 14816
rect 273352 14764 273404 14816
rect 82728 14696 82780 14748
rect 78588 14628 78640 14680
rect 269212 14628 269264 14680
rect 74448 14560 74500 14612
rect 267832 14560 267884 14612
rect 71688 14492 71740 14544
rect 265164 14492 265216 14544
rect 329932 14492 329984 14544
rect 330116 14492 330168 14544
rect 23388 14424 23440 14476
rect 241704 14424 241756 14476
rect 244188 14424 244240 14476
rect 354772 14424 354824 14476
rect 160008 14356 160060 14408
rect 311992 14356 312044 14408
rect 157248 14288 157300 14340
rect 309416 14288 309468 14340
rect 165528 14220 165580 14272
rect 313464 14220 313516 14272
rect 168288 14152 168340 14204
rect 316132 14152 316184 14204
rect 117228 14084 117280 14136
rect 246304 14084 246356 14136
rect 240048 14016 240100 14068
rect 352012 14016 352064 14068
rect 202788 13744 202840 13796
rect 334164 13744 334216 13796
rect 159916 13676 159968 13728
rect 310704 13676 310756 13728
rect 155868 13608 155920 13660
rect 309140 13608 309192 13660
rect 153108 13540 153160 13592
rect 307852 13540 307904 13592
rect 148968 13472 149020 13524
rect 305092 13472 305144 13524
rect 150348 13404 150400 13456
rect 306472 13404 306524 13456
rect 151728 13336 151780 13388
rect 307944 13336 307996 13388
rect 146208 13268 146260 13320
rect 303620 13268 303672 13320
rect 144828 13200 144880 13252
rect 303712 13200 303764 13252
rect 132408 13132 132460 13184
rect 296904 13132 296956 13184
rect 19248 13064 19300 13116
rect 238852 13064 238904 13116
rect 200028 12996 200080 13048
rect 331404 12996 331456 13048
rect 206928 12928 206980 12980
rect 335452 12928 335504 12980
rect 213828 12860 213880 12912
rect 339684 12860 339736 12912
rect 211068 12792 211120 12844
rect 336832 12792 336884 12844
rect 217968 12724 218020 12776
rect 340972 12724 341024 12776
rect 220728 12656 220780 12708
rect 342352 12656 342404 12708
rect 261024 12520 261076 12572
rect 236184 12452 236236 12504
rect 293960 12495 294012 12504
rect 293960 12461 293969 12495
rect 293969 12461 294003 12495
rect 294003 12461 294012 12495
rect 293960 12452 294012 12461
rect 397644 12452 397696 12504
rect 184848 12384 184900 12436
rect 323124 12384 323176 12436
rect 347872 12427 347924 12436
rect 347872 12393 347881 12427
rect 347881 12393 347915 12427
rect 347915 12393 347924 12427
rect 347872 12384 347924 12393
rect 397552 12384 397604 12436
rect 180708 12316 180760 12368
rect 321744 12316 321796 12368
rect 427912 12316 427964 12368
rect 428096 12316 428148 12368
rect 176568 12248 176620 12300
rect 320272 12248 320324 12300
rect 416964 12291 417016 12300
rect 416964 12257 416973 12291
rect 416973 12257 417007 12291
rect 417007 12257 417016 12291
rect 416964 12248 417016 12257
rect 173808 12180 173860 12232
rect 317604 12180 317656 12232
rect 169668 12112 169720 12164
rect 316040 12112 316092 12164
rect 166908 12044 166960 12096
rect 314752 12044 314804 12096
rect 162768 11976 162820 12028
rect 313372 11976 313424 12028
rect 142068 11908 142120 11960
rect 302424 11908 302476 11960
rect 126888 11840 126940 11892
rect 128268 11772 128320 11824
rect 295340 11772 295392 11824
rect 13636 11704 13688 11756
rect 260932 11747 260984 11756
rect 260932 11713 260941 11747
rect 260941 11713 260975 11747
rect 260975 11713 260984 11747
rect 260932 11704 260984 11713
rect 187608 11636 187660 11688
rect 325792 11636 325844 11688
rect 191748 11568 191800 11620
rect 327264 11568 327316 11620
rect 194508 11500 194560 11552
rect 328644 11500 328696 11552
rect 198648 11432 198700 11484
rect 331220 11432 331272 11484
rect 201500 11364 201552 11416
rect 332784 11364 332836 11416
rect 205548 11296 205600 11348
rect 334440 11296 334492 11348
rect 143448 10956 143500 11008
rect 302332 10956 302384 11008
rect 140688 10888 140740 10940
rect 301044 10888 301096 10940
rect 124128 10820 124180 10872
rect 292580 10820 292632 10872
rect 119988 10752 120040 10804
rect 291200 10752 291252 10804
rect 117136 10684 117188 10736
rect 288348 10684 288400 10736
rect 113088 10616 113140 10668
rect 287060 10616 287112 10668
rect 289820 10616 289872 10668
rect 367192 10616 367244 10668
rect 108764 10548 108816 10600
rect 285680 10548 285732 10600
rect 289912 10548 289964 10600
rect 367284 10548 367336 10600
rect 105176 10480 105228 10532
rect 283196 10480 283248 10532
rect 287612 10480 287664 10532
rect 365628 10480 365680 10532
rect 101588 10412 101640 10464
rect 281540 10412 281592 10464
rect 299664 10412 299716 10464
rect 379612 10412 379664 10464
rect 99196 10344 99248 10396
rect 280160 10344 280212 10396
rect 300952 10344 301004 10396
rect 383752 10344 383804 10396
rect 64788 10276 64840 10328
rect 262312 10276 262364 10328
rect 292948 10276 293000 10328
rect 378324 10276 378376 10328
rect 147588 10208 147640 10260
rect 305000 10208 305052 10260
rect 151636 10140 151688 10192
rect 306380 10140 306432 10192
rect 154488 10072 154540 10124
rect 307852 10072 307904 10124
rect 158628 10004 158680 10056
rect 310520 10004 310572 10056
rect 161388 9936 161440 9988
rect 311900 9936 311952 9988
rect 246764 9868 246816 9920
rect 356244 9868 356296 9920
rect 250352 9800 250404 9852
rect 357624 9800 357676 9852
rect 253848 9732 253900 9784
rect 360292 9732 360344 9784
rect 244280 9664 244332 9716
rect 244556 9664 244608 9716
rect 249984 9664 250036 9716
rect 250076 9664 250128 9716
rect 257436 9664 257488 9716
rect 361764 9664 361816 9716
rect 386512 9664 386564 9716
rect 386788 9664 386840 9716
rect 387892 9664 387944 9716
rect 388076 9664 388128 9716
rect 422300 9664 422352 9716
rect 422484 9664 422536 9716
rect 203892 9596 203944 9648
rect 333980 9596 334032 9648
rect 346492 9639 346544 9648
rect 346492 9605 346501 9639
rect 346501 9605 346535 9639
rect 346535 9605 346544 9639
rect 346492 9596 346544 9605
rect 393044 9639 393096 9648
rect 393044 9605 393053 9639
rect 393053 9605 393087 9639
rect 393087 9605 393096 9639
rect 393044 9596 393096 9605
rect 200396 9528 200448 9580
rect 332600 9528 332652 9580
rect 196808 9460 196860 9512
rect 330024 9460 330076 9512
rect 193220 9392 193272 9444
rect 328736 9392 328788 9444
rect 189632 9324 189684 9376
rect 327080 9324 327132 9376
rect 186044 9256 186096 9308
rect 324412 9256 324464 9308
rect 182548 9188 182600 9240
rect 323216 9188 323268 9240
rect 178960 9120 179012 9172
rect 321560 9120 321612 9172
rect 322572 9120 322624 9172
rect 361672 9256 361724 9308
rect 327080 9188 327132 9240
rect 392032 9188 392084 9240
rect 325516 9120 325568 9172
rect 390652 9120 390704 9172
rect 175372 9052 175424 9104
rect 318892 9052 318944 9104
rect 328552 9052 328604 9104
rect 394792 9052 394844 9104
rect 171784 8984 171836 9036
rect 317696 8984 317748 9036
rect 323584 8984 323636 9036
rect 389272 8984 389324 9036
rect 132592 8916 132644 8968
rect 296812 8916 296864 8968
rect 334716 8916 334768 8968
rect 401692 8916 401744 8968
rect 210976 8848 211028 8900
rect 338212 8848 338264 8900
rect 207480 8780 207532 8832
rect 335360 8780 335412 8832
rect 214656 8712 214708 8764
rect 339776 8712 339828 8764
rect 221740 8644 221792 8696
rect 343732 8644 343784 8696
rect 218152 8576 218204 8628
rect 340880 8576 340932 8628
rect 225328 8508 225380 8560
rect 345204 8508 345256 8560
rect 228916 8440 228968 8492
rect 232504 8372 232556 8424
rect 349252 8372 349304 8424
rect 230664 8347 230716 8356
rect 230664 8313 230673 8347
rect 230673 8313 230707 8347
rect 230707 8313 230716 8347
rect 230664 8304 230716 8313
rect 236000 8304 236052 8356
rect 350724 8304 350776 8356
rect 380992 8347 381044 8356
rect 380992 8313 381001 8347
rect 381001 8313 381035 8347
rect 381035 8313 381044 8347
rect 380992 8304 381044 8313
rect 382372 8347 382424 8356
rect 382372 8313 382381 8347
rect 382381 8313 382415 8347
rect 382415 8313 382424 8347
rect 382372 8304 382424 8313
rect 400404 8347 400456 8356
rect 400404 8313 400413 8347
rect 400413 8313 400447 8347
rect 400447 8313 400456 8347
rect 400404 8304 400456 8313
rect 56416 8236 56468 8288
rect 258356 8236 258408 8288
rect 274088 8236 274140 8288
rect 370136 8236 370188 8288
rect 52828 8168 52880 8220
rect 256792 8168 256844 8220
rect 270500 8168 270552 8220
rect 368572 8168 368624 8220
rect 49332 8100 49384 8152
rect 254032 8100 254084 8152
rect 267004 8100 267056 8152
rect 367100 8100 367152 8152
rect 44548 8032 44600 8084
rect 252652 8032 252704 8084
rect 263416 8032 263468 8084
rect 364524 8032 364576 8084
rect 40960 7964 41012 8016
rect 249984 7964 250036 8016
rect 259828 7964 259880 8016
rect 363052 7964 363104 8016
rect 37372 7896 37424 7948
rect 248512 7896 248564 7948
rect 256240 7896 256292 7948
rect 361580 7896 361632 7948
rect 33876 7828 33928 7880
rect 247224 7828 247276 7880
rect 252652 7828 252704 7880
rect 359004 7828 359056 7880
rect 30288 7760 30340 7812
rect 244280 7760 244332 7812
rect 249156 7760 249208 7812
rect 357440 7760 357492 7812
rect 26700 7692 26752 7744
rect 242900 7692 242952 7744
rect 245568 7692 245620 7744
rect 356152 7692 356204 7744
rect 8852 7624 8904 7676
rect 233332 7624 233384 7676
rect 234804 7624 234856 7676
rect 350632 7624 350684 7676
rect 3976 7556 4028 7608
rect 230664 7556 230716 7608
rect 231308 7556 231360 7608
rect 347872 7556 347924 7608
rect 351828 7556 351880 7608
rect 405832 7556 405884 7608
rect 87328 7488 87380 7540
rect 274640 7488 274692 7540
rect 277676 7488 277728 7540
rect 372712 7488 372764 7540
rect 90916 7420 90968 7472
rect 276020 7420 276072 7472
rect 281264 7420 281316 7472
rect 374092 7420 374144 7472
rect 94504 7352 94556 7404
rect 277584 7352 277636 7404
rect 284760 7352 284812 7404
rect 375564 7352 375616 7404
rect 138480 7284 138532 7336
rect 300860 7284 300912 7336
rect 347964 7284 348016 7336
rect 397552 7284 397604 7336
rect 141976 7216 142028 7268
rect 302516 7216 302568 7268
rect 346492 7216 346544 7268
rect 396172 7216 396224 7268
rect 224132 7148 224184 7200
rect 345112 7148 345164 7200
rect 227720 7080 227772 7132
rect 346400 7080 346452 7132
rect 238392 7012 238444 7064
rect 351920 7012 351972 7064
rect 241980 6944 242032 6996
rect 353392 6944 353444 6996
rect 163504 6808 163556 6860
rect 313556 6808 313608 6860
rect 349068 6808 349120 6860
rect 408776 6808 408828 6860
rect 83832 6740 83884 6792
rect 271880 6740 271932 6792
rect 320180 6740 320232 6792
rect 325608 6740 325660 6792
rect 386512 6740 386564 6792
rect 80244 6672 80296 6724
rect 270592 6672 270644 6724
rect 318800 6672 318852 6724
rect 380992 6672 381044 6724
rect 76656 6604 76708 6656
rect 269120 6604 269172 6656
rect 320180 6604 320232 6656
rect 385132 6604 385184 6656
rect 73068 6536 73120 6588
rect 266360 6536 266412 6588
rect 312176 6536 312228 6588
rect 389364 6536 389416 6588
rect 69480 6468 69532 6520
rect 264980 6468 265032 6520
rect 308588 6468 308640 6520
rect 387892 6468 387944 6520
rect 62396 6400 62448 6452
rect 260932 6400 260984 6452
rect 305000 6400 305052 6452
rect 386420 6400 386472 6452
rect 65984 6332 66036 6384
rect 263692 6332 263744 6384
rect 290740 6332 290792 6384
rect 378232 6332 378284 6384
rect 58808 6264 58860 6316
rect 259460 6264 259512 6316
rect 287152 6264 287204 6316
rect 376944 6264 376996 6316
rect 55220 6196 55272 6248
rect 258264 6196 258316 6248
rect 283656 6196 283708 6248
rect 375380 6196 375432 6248
rect 379980 6196 380032 6248
rect 425152 6196 425204 6248
rect 51632 6128 51684 6180
rect 255320 6128 255372 6180
rect 279976 6128 280028 6180
rect 372804 6128 372856 6180
rect 372896 6128 372948 6180
rect 421104 6128 421156 6180
rect 167092 6060 167144 6112
rect 314568 6060 314620 6112
rect 314660 6060 314712 6112
rect 371332 6060 371384 6112
rect 170588 5992 170640 6044
rect 317420 5992 317472 6044
rect 322940 5992 322992 6044
rect 354956 5992 355008 6044
rect 411352 5992 411404 6044
rect 174176 5924 174228 5976
rect 177764 5856 177816 5908
rect 316592 5924 316644 5976
rect 369860 5924 369912 5976
rect 318892 5856 318944 5908
rect 325332 5856 325384 5908
rect 360200 5856 360252 5908
rect 362132 5856 362184 5908
rect 415584 5856 415636 5908
rect 181352 5788 181404 5840
rect 322664 5788 322716 5840
rect 364340 5788 364392 5840
rect 369216 5788 369268 5840
rect 419632 5788 419684 5840
rect 184848 5720 184900 5772
rect 324320 5720 324372 5772
rect 188436 5652 188488 5704
rect 325700 5652 325752 5704
rect 192024 5584 192076 5636
rect 328460 5584 328512 5636
rect 195612 5516 195664 5568
rect 329840 5516 329892 5568
rect 137284 5448 137336 5500
rect 299480 5448 299532 5500
rect 315764 5448 315816 5500
rect 391940 5448 391992 5500
rect 401324 5448 401376 5500
rect 436192 5448 436244 5500
rect 133788 5380 133840 5432
rect 298100 5380 298152 5432
rect 301412 5380 301464 5432
rect 383844 5380 383896 5432
rect 397828 5380 397880 5432
rect 433616 5380 433668 5432
rect 130200 5312 130252 5364
rect 296720 5312 296772 5364
rect 297916 5312 297968 5364
rect 382372 5312 382424 5364
rect 394240 5312 394292 5364
rect 432144 5312 432196 5364
rect 67180 5244 67232 5296
rect 263784 5244 263836 5296
rect 294328 5244 294380 5296
rect 380900 5244 380952 5296
rect 390652 5244 390704 5296
rect 430672 5244 430724 5296
rect 21916 5176 21968 5228
rect 240232 5176 240284 5228
rect 251456 5176 251508 5228
rect 358820 5176 358872 5228
rect 387064 5176 387116 5228
rect 427912 5176 427964 5228
rect 17316 5108 17368 5160
rect 237472 5108 237524 5160
rect 247960 5108 248012 5160
rect 356428 5108 356480 5160
rect 383568 5108 383620 5160
rect 426716 5108 426768 5160
rect 12440 5040 12492 5092
rect 236092 5040 236144 5092
rect 244372 5040 244424 5092
rect 354680 5040 354732 5092
rect 376392 5040 376444 5092
rect 422300 5040 422352 5092
rect 7656 4972 7708 5024
rect 233240 4972 233292 5024
rect 240784 4972 240836 5024
rect 353300 4972 353352 5024
rect 365720 4972 365772 5024
rect 416964 4972 417016 5024
rect 2872 4904 2924 4956
rect 230480 4904 230532 4956
rect 237196 4904 237248 4956
rect 350540 4904 350592 4956
rect 358544 4904 358596 4956
rect 414112 4904 414164 4956
rect 503536 4904 503588 4956
rect 529664 4904 529716 4956
rect 572 4836 624 4888
rect 229100 4836 229152 4888
rect 230112 4836 230164 4888
rect 347780 4836 347832 4888
rect 347872 4836 347924 4888
rect 408500 4836 408552 4888
rect 509148 4836 509200 4888
rect 540520 4836 540572 4888
rect 1676 4768 1728 4820
rect 230572 4768 230624 4820
rect 233700 4768 233752 4820
rect 349160 4768 349212 4820
rect 351368 4768 351420 4820
rect 410064 4768 410116 4820
rect 506296 4768 506348 4820
rect 536932 4768 536984 4820
rect 215852 4700 215904 4752
rect 339500 4700 339552 4752
rect 340696 4700 340748 4752
rect 404544 4700 404596 4752
rect 404912 4700 404964 4752
rect 437756 4700 437808 4752
rect 222936 4632 222988 4684
rect 343640 4632 343692 4684
rect 344284 4632 344336 4684
rect 405924 4632 405976 4684
rect 226524 4564 226576 4616
rect 345020 4564 345072 4616
rect 356060 4564 356112 4616
rect 362960 4564 363012 4616
rect 208676 4496 208728 4548
rect 283564 4496 283616 4548
rect 319260 4496 319312 4548
rect 393504 4496 393556 4548
rect 212264 4428 212316 4480
rect 284944 4428 284996 4480
rect 322848 4428 322900 4480
rect 394884 4428 394936 4480
rect 326436 4360 326488 4412
rect 397460 4360 397512 4412
rect 330024 4292 330076 4344
rect 399024 4292 399076 4344
rect 333612 4224 333664 4276
rect 400404 4224 400456 4276
rect 408684 4224 408736 4276
rect 124220 4156 124272 4208
rect 125416 4156 125468 4208
rect 140872 4156 140924 4208
rect 142068 4156 142120 4208
rect 150440 4156 150492 4208
rect 151636 4156 151688 4208
rect 158720 4156 158772 4208
rect 159916 4156 159968 4208
rect 209872 4156 209924 4208
rect 211068 4156 211120 4208
rect 42156 4088 42208 4140
rect 50344 4088 50396 4140
rect 57612 4088 57664 4140
rect 255964 4088 256016 4140
rect 275284 4088 275336 4140
rect 276664 4088 276716 4140
rect 278872 4088 278924 4140
rect 280068 4088 280120 4140
rect 314660 4156 314712 4208
rect 337108 4156 337160 4208
rect 403072 4156 403124 4208
rect 405004 4156 405056 4208
rect 314568 4088 314620 4140
rect 316684 4088 316736 4140
rect 321652 4088 321704 4140
rect 322756 4088 322808 4140
rect 331220 4088 331272 4140
rect 332508 4088 332560 4140
rect 346676 4088 346728 4140
rect 50528 4020 50580 4072
rect 253204 4020 253256 4072
rect 262220 4020 262272 4072
rect 322664 4020 322716 4072
rect 339500 4020 339552 4072
rect 400220 4088 400272 4140
rect 408408 4088 408460 4140
rect 408592 4156 408644 4208
rect 410524 4088 410576 4140
rect 403532 4020 403584 4072
rect 34980 3952 35032 4004
rect 46204 3952 46256 4004
rect 46940 3952 46992 4004
rect 252744 3952 252796 4004
rect 271696 3952 271748 4004
rect 283472 3952 283524 4004
rect 300308 3952 300360 4004
rect 363604 3952 363656 4004
rect 364524 3952 364576 4004
rect 366364 3952 366416 4004
rect 371608 3952 371660 4004
rect 372528 3952 372580 4004
rect 409144 4020 409196 4072
rect 411904 4088 411956 4140
rect 412088 4088 412140 4140
rect 412548 4088 412600 4140
rect 414480 4088 414532 4140
rect 416044 4088 416096 4140
rect 419172 4088 419224 4140
rect 420184 4088 420236 4140
rect 420368 4088 420420 4140
rect 420828 4088 420880 4140
rect 422760 4088 422812 4140
rect 423588 4088 423640 4140
rect 423956 4088 424008 4140
rect 424968 4088 425020 4140
rect 429292 4088 429344 4140
rect 429936 4088 429988 4140
rect 430488 4088 430540 4140
rect 431132 4088 431184 4140
rect 431868 4088 431920 4140
rect 433524 4088 433576 4140
rect 434628 4088 434680 4140
rect 437020 4088 437072 4140
rect 442356 4088 442408 4140
rect 451280 4088 451332 4140
rect 453304 4088 453356 4140
rect 454868 4088 454920 4140
rect 456064 4088 456116 4140
rect 469128 4088 469180 4140
rect 469864 4088 469916 4140
rect 472164 4088 472216 4140
rect 472716 4088 472768 4140
rect 473360 4088 473412 4140
rect 473912 4088 473964 4140
rect 474648 4088 474700 4140
rect 475108 4088 475160 4140
rect 493968 4088 494020 4140
rect 512000 4088 512052 4140
rect 518808 4088 518860 4140
rect 559564 4088 559616 4140
rect 410892 4020 410944 4072
rect 413284 4020 413336 4072
rect 438952 4020 439004 4072
rect 440608 4020 440660 4072
rect 445024 4020 445076 4072
rect 492496 4020 492548 4072
rect 509608 4020 509660 4072
rect 520096 4020 520148 4072
rect 561956 4020 562008 4072
rect 408684 3952 408736 4004
rect 420276 3952 420328 4004
rect 424416 3952 424468 4004
rect 427544 3952 427596 4004
rect 45744 3884 45796 3936
rect 251824 3884 251876 3936
rect 258632 3884 258684 3936
rect 322572 3884 322624 3936
rect 325240 3884 325292 3936
rect 391112 3884 391164 3936
rect 400864 3884 400916 3936
rect 408592 3884 408644 3936
rect 425152 3884 425204 3936
rect 448520 3952 448572 4004
rect 458456 3952 458508 4004
rect 464436 3952 464488 4004
rect 493876 3952 493928 4004
rect 513196 3952 513248 4004
rect 520188 3952 520240 4004
rect 564348 3952 564400 4004
rect 565084 3952 565136 4004
rect 579804 3952 579856 4004
rect 442264 3884 442316 3936
rect 496084 3884 496136 3936
rect 39764 3816 39816 3868
rect 249800 3816 249852 3868
rect 255044 3816 255096 3868
rect 38568 3748 38620 3800
rect 248420 3748 248472 3800
rect 272892 3748 272944 3800
rect 316592 3748 316644 3800
rect 32680 3680 32732 3732
rect 245660 3680 245712 3732
rect 264612 3680 264664 3732
rect 287704 3680 287756 3732
rect 299112 3680 299164 3732
rect 300952 3680 301004 3732
rect 307392 3680 307444 3732
rect 309784 3680 309836 3732
rect 316960 3816 317012 3868
rect 327080 3816 327132 3868
rect 332416 3816 332468 3868
rect 318064 3748 318116 3800
rect 389824 3748 389876 3800
rect 396724 3816 396776 3868
rect 403716 3816 403768 3868
rect 437664 3816 437716 3868
rect 448980 3816 449032 3868
rect 453396 3816 453448 3868
rect 482928 3816 482980 3868
rect 490564 3816 490616 3868
rect 496728 3816 496780 3868
rect 509884 3884 509936 3936
rect 520280 3884 520332 3936
rect 521568 3884 521620 3936
rect 566740 3884 566792 3936
rect 515588 3816 515640 3868
rect 516784 3816 516836 3868
rect 395344 3748 395396 3800
rect 399024 3748 399076 3800
rect 434812 3748 434864 3800
rect 438216 3748 438268 3800
rect 447784 3748 447836 3800
rect 325332 3680 325384 3732
rect 352564 3680 352616 3732
rect 353208 3680 353260 3732
rect 385868 3680 385920 3732
rect 25504 3612 25556 3664
rect 239588 3612 239640 3664
rect 240048 3612 240100 3664
rect 243176 3612 243228 3664
rect 244188 3612 244240 3664
rect 269304 3612 269356 3664
rect 289820 3612 289872 3664
rect 291936 3612 291988 3664
rect 299664 3612 299716 3664
rect 303804 3612 303856 3664
rect 382924 3612 382976 3664
rect 388260 3612 388312 3664
rect 389088 3612 389140 3664
rect 391848 3612 391900 3664
rect 408316 3612 408368 3664
rect 408500 3612 408552 3664
rect 408592 3612 408644 3664
rect 18328 3544 18380 3596
rect 19248 3544 19300 3596
rect 19524 3544 19576 3596
rect 24124 3544 24176 3596
rect 24308 3544 24360 3596
rect 241520 3544 241572 3596
rect 14832 3476 14884 3528
rect 236368 3476 236420 3528
rect 241796 3476 241848 3528
rect 265808 3476 265860 3528
rect 287612 3476 287664 3528
rect 289544 3544 289596 3596
rect 296720 3544 296772 3596
rect 381544 3544 381596 3596
rect 389456 3544 389508 3596
rect 434536 3680 434588 3732
rect 446496 3680 446548 3732
rect 455604 3748 455656 3800
rect 489184 3748 489236 3800
rect 497740 3748 497792 3800
rect 498844 3748 498896 3800
rect 519084 3748 519136 3800
rect 450176 3680 450228 3732
rect 451188 3680 451240 3732
rect 457260 3680 457312 3732
rect 465356 3680 465408 3732
rect 466828 3680 466880 3732
rect 467748 3680 467800 3732
rect 485688 3680 485740 3732
rect 495348 3680 495400 3732
rect 499488 3680 499540 3732
rect 522672 3680 522724 3732
rect 525064 3816 525116 3868
rect 525616 3816 525668 3868
rect 572628 3816 572680 3868
rect 522948 3748 523000 3800
rect 569040 3748 569092 3800
rect 432604 3612 432656 3664
rect 443000 3612 443052 3664
rect 456892 3612 456944 3664
rect 478788 3612 478840 3664
rect 482284 3612 482336 3664
rect 484216 3612 484268 3664
rect 492956 3612 493008 3664
rect 500776 3612 500828 3664
rect 289912 3476 289964 3528
rect 378416 3476 378468 3528
rect 382372 3476 382424 3528
rect 433340 3544 433392 3596
rect 439412 3544 439464 3596
rect 447784 3544 447836 3596
rect 448428 3544 448480 3596
rect 467932 3544 467984 3596
rect 470784 3544 470836 3596
rect 484308 3544 484360 3596
rect 494152 3544 494204 3596
rect 499396 3544 499448 3596
rect 523868 3544 523920 3596
rect 524328 3680 524380 3732
rect 571432 3680 571484 3732
rect 525524 3612 525576 3664
rect 573824 3612 573876 3664
rect 527456 3544 527508 3596
rect 529848 3544 529900 3596
rect 582196 3544 582248 3596
rect 426348 3476 426400 3528
rect 428464 3476 428516 3528
rect 432328 3476 432380 3528
rect 451556 3476 451608 3528
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 16028 3408 16080 3460
rect 237564 3408 237616 3460
rect 261024 3408 261076 3460
rect 356060 3408 356112 3460
rect 368020 3408 368072 3460
rect 402520 3408 402572 3460
rect 36176 3340 36228 3392
rect 39304 3340 39356 3392
rect 11244 3272 11296 3324
rect 17224 3272 17276 3324
rect 20720 3272 20772 3324
rect 28264 3272 28316 3324
rect 43352 3204 43404 3256
rect 54024 3272 54076 3324
rect 57244 3272 57296 3324
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 63592 3340 63644 3392
rect 64788 3340 64840 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 61384 3272 61436 3324
rect 64788 3204 64840 3256
rect 257344 3340 257396 3392
rect 268108 3340 268160 3392
rect 282460 3340 282512 3392
rect 294604 3340 294656 3392
rect 295524 3340 295576 3392
rect 318800 3340 318852 3392
rect 324044 3340 324096 3392
rect 346492 3340 346544 3392
rect 353760 3340 353812 3392
rect 396632 3340 396684 3392
rect 408500 3408 408552 3460
rect 409788 3408 409840 3460
rect 412640 3408 412692 3460
rect 413468 3408 413520 3460
rect 71872 3272 71924 3324
rect 258724 3272 258776 3324
rect 276480 3272 276532 3324
rect 306196 3272 306248 3324
rect 325608 3272 325660 3324
rect 347964 3272 348016 3324
rect 366456 3272 366508 3324
rect 77852 3204 77904 3256
rect 78588 3204 78640 3256
rect 81440 3204 81492 3256
rect 82728 3204 82780 3256
rect 27896 3136 27948 3188
rect 28908 3136 28960 3188
rect 29092 3136 29144 3188
rect 32404 3136 32456 3188
rect 61200 3136 61252 3188
rect 66904 3136 66956 3188
rect 82636 3136 82688 3188
rect 84844 3204 84896 3256
rect 84936 3204 84988 3256
rect 85488 3204 85540 3256
rect 88524 3204 88576 3256
rect 89628 3204 89680 3256
rect 261484 3204 261536 3256
rect 288348 3204 288400 3256
rect 292948 3204 293000 3256
rect 302608 3204 302660 3256
rect 320180 3204 320232 3256
rect 328828 3204 328880 3256
rect 363696 3204 363748 3256
rect 89812 3136 89864 3188
rect 262864 3136 262916 3188
rect 285956 3136 286008 3188
rect 286968 3136 287020 3188
rect 293132 3136 293184 3188
rect 293868 3136 293920 3188
rect 309784 3136 309836 3188
rect 323584 3136 323636 3188
rect 327632 3136 327684 3188
rect 343088 3136 343140 3188
rect 95700 3068 95752 3120
rect 96528 3068 96580 3120
rect 10048 3000 10100 3052
rect 15844 3000 15896 3052
rect 68284 3000 68336 3052
rect 71044 3000 71096 3052
rect 93308 3000 93360 3052
rect 97264 3068 97316 3120
rect 98092 3068 98144 3120
rect 99196 3068 99248 3120
rect 102784 3068 102836 3120
rect 103428 3068 103480 3120
rect 103980 3068 104032 3120
rect 104808 3068 104860 3120
rect 106372 3068 106424 3120
rect 107568 3068 107620 3120
rect 111156 3068 111208 3120
rect 111708 3068 111760 3120
rect 96896 3000 96948 3052
rect 264244 3068 264296 3120
rect 313372 3068 313424 3120
rect 325516 3068 325568 3120
rect 335912 3068 335964 3120
rect 363328 3068 363380 3120
rect 370412 3204 370464 3256
rect 407120 3272 407172 3324
rect 407304 3272 407356 3324
rect 417424 3340 417476 3392
rect 417976 3340 418028 3392
rect 435364 3340 435416 3392
rect 444196 3408 444248 3460
rect 446404 3408 446456 3460
rect 446588 3408 446640 3460
rect 459744 3476 459796 3528
rect 487068 3476 487120 3528
rect 498936 3476 498988 3528
rect 500868 3476 500920 3528
rect 526260 3476 526312 3528
rect 528468 3476 528520 3528
rect 578608 3476 578660 3528
rect 452476 3408 452528 3460
rect 457444 3408 457496 3460
rect 462044 3408 462096 3460
rect 466460 3408 466512 3460
rect 488448 3408 488500 3460
rect 501236 3408 501288 3460
rect 502248 3408 502300 3460
rect 528652 3408 528704 3460
rect 529756 3408 529808 3460
rect 581000 3408 581052 3460
rect 444564 3340 444616 3392
rect 459652 3340 459704 3392
rect 464344 3340 464396 3392
rect 482836 3340 482888 3392
rect 489368 3340 489420 3392
rect 492588 3340 492640 3392
rect 508412 3340 508464 3392
rect 516784 3340 516836 3392
rect 517428 3340 517480 3392
rect 557172 3340 557224 3392
rect 558184 3340 558236 3392
rect 409696 3272 409748 3324
rect 431224 3272 431276 3324
rect 441804 3272 441856 3324
rect 449164 3272 449216 3324
rect 464436 3272 464488 3324
rect 464988 3272 465040 3324
rect 481548 3272 481600 3324
rect 486976 3272 487028 3324
rect 488356 3272 488408 3324
rect 502432 3272 502484 3324
rect 514668 3272 514720 3324
rect 552388 3272 552440 3324
rect 556804 3272 556856 3324
rect 565544 3272 565596 3324
rect 381176 3136 381228 3188
rect 79048 2932 79100 2984
rect 86132 2932 86184 2984
rect 75460 2864 75512 2916
rect 106924 2932 106976 2984
rect 100484 2864 100536 2916
rect 264336 3000 264388 3052
rect 320456 3000 320508 3052
rect 328552 3000 328604 3052
rect 338304 3000 338356 3052
rect 339408 3000 339460 3052
rect 350264 3000 350316 3052
rect 374644 3068 374696 3120
rect 375196 3068 375248 3120
rect 413376 3204 413428 3256
rect 416872 3204 416924 3256
rect 438124 3204 438176 3256
rect 485044 3204 485096 3256
rect 488172 3204 488224 3256
rect 489828 3204 489880 3256
rect 504824 3204 504876 3256
rect 511816 3204 511868 3256
rect 540244 3204 540296 3256
rect 541716 3204 541768 3256
rect 547144 3204 547196 3256
rect 550088 3204 550140 3256
rect 403624 3068 403676 3120
rect 374000 3000 374052 3052
rect 375288 3000 375340 3052
rect 378876 3000 378928 3052
rect 414664 3068 414716 3120
rect 415676 3068 415728 3120
rect 416688 3068 416740 3120
rect 430580 3136 430632 3188
rect 493324 3136 493376 3188
rect 496544 3136 496596 3188
rect 510528 3136 510580 3188
rect 424324 3068 424376 3120
rect 470324 3068 470376 3120
rect 470692 3068 470744 3120
rect 501604 3068 501656 3120
rect 506020 3068 506072 3120
rect 511908 3068 511960 3120
rect 540336 3136 540388 3188
rect 544108 3136 544160 3188
rect 112352 2932 112404 2984
rect 113088 2932 113140 2984
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 115940 2932 115992 2984
rect 116952 2932 117004 2984
rect 119436 2932 119488 2984
rect 119988 2932 120040 2984
rect 120632 2932 120684 2984
rect 121368 2932 121420 2984
rect 114744 2864 114796 2916
rect 105544 2796 105596 2848
rect 107568 2796 107620 2848
rect 266912 2932 266964 2984
rect 341892 2932 341944 2984
rect 351828 2932 351880 2984
rect 360936 2932 360988 2984
rect 377588 2932 377640 2984
rect 406108 2932 406160 2984
rect 409144 2932 409196 2984
rect 268384 2864 268436 2916
rect 376024 2864 376076 2916
rect 384672 2864 384724 2916
rect 412640 3000 412692 3052
rect 409420 2932 409472 2984
rect 427084 3000 427136 3052
rect 445392 3000 445444 3052
rect 451924 3000 451976 3052
rect 477408 3000 477460 3052
rect 479892 3000 479944 3052
rect 507768 3000 507820 3052
rect 538128 3000 538180 3052
rect 545304 3068 545356 3120
rect 545764 3068 545816 3120
rect 554780 3068 554832 3120
rect 546500 3000 546552 3052
rect 547236 3000 547288 3052
rect 548892 3000 548944 3052
rect 549904 3000 549956 3052
rect 558368 3204 558420 3256
rect 569224 3340 569276 3392
rect 570236 3340 570288 3392
rect 576216 3204 576268 3256
rect 571984 3000 572036 3052
rect 577412 3000 577464 3052
rect 426624 2932 426676 2984
rect 506388 2932 506440 2984
rect 535736 2932 535788 2984
rect 547696 2932 547748 2984
rect 416044 2864 416096 2916
rect 421564 2864 421616 2916
rect 422208 2864 422260 2916
rect 465632 2864 465684 2916
rect 466368 2864 466420 2916
rect 505008 2864 505060 2916
rect 533436 2864 533488 2916
rect 121828 2796 121880 2848
rect 269764 2796 269816 2848
rect 310980 2796 311032 2848
rect 385684 2796 385736 2848
rect 395436 2796 395488 2848
rect 460204 2796 460256 2848
rect 463240 2796 463292 2848
rect 463608 2796 463660 2848
rect 471520 2796 471572 2848
rect 471888 2796 471940 2848
rect 503720 2796 503772 2848
rect 531044 2796 531096 2848
rect 543004 2796 543056 2848
rect 551192 2932 551244 2984
rect 456064 2728 456116 2780
rect 345480 688 345532 740
rect 346308 688 346360 740
rect 139676 552 139728 604
rect 140688 552 140740 604
rect 172980 552 173032 604
rect 173808 552 173860 604
rect 180156 552 180208 604
rect 180708 552 180760 604
rect 205088 552 205140 604
rect 205548 552 205600 604
rect 206284 552 206336 604
rect 206928 552 206980 604
rect 220544 552 220596 604
rect 220728 552 220780 604
rect 393044 595 393096 604
rect 393044 561 393053 595
rect 393053 561 393087 595
rect 393087 561 393096 595
rect 393044 552 393096 561
rect 413284 552 413336 604
rect 435824 552 435876 604
rect 436008 552 436060 604
rect 453672 552 453724 604
rect 453948 552 454000 604
rect 477776 552 477828 604
rect 478696 552 478748 604
rect 480352 552 480404 604
rect 481088 552 481140 604
rect 499764 552 499816 604
rect 500132 552 500184 604
rect 506664 552 506716 604
rect 507216 552 507268 604
rect 513564 552 513616 604
rect 514392 552 514444 604
rect 520372 552 520424 604
rect 521476 552 521528 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 105464 700602 105492 703520
rect 137848 700670 137876 703520
rect 154132 700738 154160 703520
rect 170324 700806 170352 703520
rect 202800 700874 202828 703520
rect 218992 701010 219020 703520
rect 218980 701004 219032 701010
rect 218980 700946 219032 700952
rect 202788 700868 202840 700874
rect 202788 700810 202840 700816
rect 170312 700800 170364 700806
rect 170312 700742 170364 700748
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 105452 700596 105504 700602
rect 105452 700538 105504 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 235184 699718 235212 703520
rect 267660 700194 267688 703520
rect 267648 700188 267700 700194
rect 267648 700130 267700 700136
rect 283852 699990 283880 703520
rect 283840 699984 283892 699990
rect 283840 699926 283892 699932
rect 300136 699718 300164 703520
rect 332520 699922 332548 703520
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 348804 699786 348832 703520
rect 355968 700936 356020 700942
rect 355968 700878 356020 700884
rect 353208 700256 353260 700262
rect 353208 700198 353260 700204
rect 348792 699780 348844 699786
rect 348792 699722 348844 699728
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 235920 643822 235948 699654
rect 269028 670744 269080 670750
rect 269028 670686 269080 670692
rect 235908 643816 235960 643822
rect 235908 643758 235960 643764
rect 3514 643104 3570 643113
rect 3514 643039 3570 643048
rect 3332 639736 3384 639742
rect 3332 639678 3384 639684
rect 3240 624912 3292 624918
rect 3238 624880 3240 624889
rect 3292 624880 3294 624889
rect 3238 624815 3294 624824
rect 2780 610632 2832 610638
rect 2780 610574 2832 610580
rect 2792 610473 2820 610574
rect 2778 610464 2834 610473
rect 2778 610399 2834 610408
rect 3240 596080 3292 596086
rect 3238 596048 3240 596057
rect 3292 596048 3294 596057
rect 3238 595983 3294 595992
rect 3240 567792 3292 567798
rect 3240 567734 3292 567740
rect 3252 567361 3280 567734
rect 3238 567352 3294 567361
rect 3238 567287 3294 567296
rect 2780 553104 2832 553110
rect 2778 553072 2780 553081
rect 2832 553072 2834 553081
rect 2778 553007 2834 553016
rect 3240 539572 3292 539578
rect 3240 539514 3292 539520
rect 3252 538665 3280 539514
rect 3238 538656 3294 538665
rect 3238 538591 3294 538600
rect 3240 510400 3292 510406
rect 3240 510342 3292 510348
rect 3252 509969 3280 510342
rect 3238 509960 3294 509969
rect 3238 509895 3294 509904
rect 2780 496732 2832 496738
rect 2780 496674 2832 496680
rect 2792 495553 2820 496674
rect 2778 495544 2834 495553
rect 2778 495479 2834 495488
rect 3240 481160 3292 481166
rect 3238 481128 3240 481137
rect 3292 481128 3294 481137
rect 3238 481063 3294 481072
rect 3148 452464 3200 452470
rect 3146 452432 3148 452441
rect 3200 452432 3202 452441
rect 3146 452367 3202 452376
rect 3148 438796 3200 438802
rect 3148 438738 3200 438744
rect 3160 438025 3188 438738
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 3344 423745 3372 639678
rect 3422 639568 3478 639577
rect 3422 639503 3478 639512
rect 3330 423736 3386 423745
rect 3330 423671 3386 423680
rect 3148 395480 3200 395486
rect 3148 395422 3200 395428
rect 3160 395049 3188 395422
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 2780 380656 2832 380662
rect 2778 380624 2780 380633
rect 2832 380624 2834 380633
rect 2778 380559 2834 380568
rect 3332 366512 3384 366518
rect 3332 366454 3384 366460
rect 3344 366217 3372 366454
rect 3330 366208 3386 366217
rect 3330 366143 3386 366152
rect 3240 337952 3292 337958
rect 3240 337894 3292 337900
rect 3252 337521 3280 337894
rect 3238 337512 3294 337521
rect 3238 337447 3294 337456
rect 2780 323604 2832 323610
rect 2780 323546 2832 323552
rect 2792 323105 2820 323546
rect 2778 323096 2834 323105
rect 2778 323031 2834 323040
rect 3332 294432 3384 294438
rect 3330 294400 3332 294409
rect 3384 294400 3386 294409
rect 3330 294335 3386 294344
rect 3148 280152 3200 280158
rect 3146 280120 3148 280129
rect 3200 280120 3202 280129
rect 3146 280055 3202 280064
rect 3332 266348 3384 266354
rect 3332 266290 3384 266296
rect 3344 265713 3372 266290
rect 3330 265704 3386 265713
rect 3330 265639 3386 265648
rect 3146 252512 3202 252521
rect 3146 252447 3202 252456
rect 3160 251297 3188 252447
rect 3146 251288 3202 251297
rect 3146 251223 3202 251232
rect 2780 237312 2832 237318
rect 2780 237254 2832 237260
rect 2792 237017 2820 237254
rect 2778 237008 2834 237017
rect 2778 236943 2834 236952
rect 3148 194336 3200 194342
rect 3148 194278 3200 194284
rect 3160 193905 3188 194278
rect 3146 193896 3202 193905
rect 3146 193831 3202 193840
rect 2780 179512 2832 179518
rect 2778 179480 2780 179489
rect 2832 179480 2834 179489
rect 2778 179415 2834 179424
rect 2780 79892 2832 79898
rect 2780 79834 2832 79840
rect 2792 78985 2820 79834
rect 2778 78976 2834 78985
rect 2778 78911 2834 78920
rect 3436 50153 3464 639503
rect 3528 64569 3556 643039
rect 259918 642968 259974 642977
rect 259918 642903 259974 642912
rect 258722 642832 258778 642841
rect 258722 642767 258778 642776
rect 236276 642592 236328 642598
rect 236276 642534 236328 642540
rect 86224 642320 86276 642326
rect 86224 642262 86276 642268
rect 5448 642252 5500 642258
rect 5448 642194 5500 642200
rect 5356 642184 5408 642190
rect 5356 642126 5408 642132
rect 5264 642048 5316 642054
rect 4894 642016 4950 642025
rect 5264 641990 5316 641996
rect 4894 641951 4950 641960
rect 3698 641880 3754 641889
rect 3698 641815 3754 641824
rect 3606 639024 3662 639033
rect 3606 638959 3662 638968
rect 3620 107681 3648 638959
rect 3606 107672 3662 107681
rect 3606 107607 3662 107616
rect 3712 93265 3740 641815
rect 3976 641028 4028 641034
rect 3976 640970 4028 640976
rect 3882 639704 3938 639713
rect 3882 639639 3938 639648
rect 3790 638208 3846 638217
rect 3790 638143 3846 638152
rect 3804 122097 3832 638143
rect 3896 136377 3924 639639
rect 3988 150793 4016 640970
rect 4804 640348 4856 640354
rect 4804 640290 4856 640296
rect 4158 639840 4214 639849
rect 4158 639775 4214 639784
rect 4068 639668 4120 639674
rect 4068 639610 4120 639616
rect 4080 222601 4108 639610
rect 4066 222592 4122 222601
rect 4066 222527 4122 222536
rect 3974 150784 4030 150793
rect 3974 150719 4030 150728
rect 3882 136368 3938 136377
rect 3882 136303 3938 136312
rect 3790 122088 3846 122097
rect 3790 122023 3846 122032
rect 3698 93256 3754 93265
rect 3698 93191 3754 93200
rect 3514 64560 3570 64569
rect 3514 64495 3570 64504
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3976 7608 4028 7614
rect 3976 7550 4028 7556
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4898
rect 3988 626 4016 7550
rect 4066 7168 4122 7177
rect 4172 7154 4200 639775
rect 4816 79898 4844 640290
rect 4908 179518 4936 641951
rect 5172 641912 5224 641918
rect 5172 641854 5224 641860
rect 5080 641844 5132 641850
rect 5080 641786 5132 641792
rect 4988 641776 5040 641782
rect 4988 641718 5040 641724
rect 5000 237318 5028 641718
rect 5092 323610 5120 641786
rect 5184 380662 5212 641854
rect 5276 496738 5304 641990
rect 5368 553110 5396 642126
rect 5460 610638 5488 642194
rect 72422 642152 72478 642161
rect 7932 642116 7984 642122
rect 72422 642087 72478 642096
rect 7932 642058 7984 642064
rect 7656 641980 7708 641986
rect 7656 641922 7708 641928
rect 6552 640688 6604 640694
rect 6552 640630 6604 640636
rect 6460 640620 6512 640626
rect 6460 640562 6512 640568
rect 6368 640484 6420 640490
rect 6368 640426 6420 640432
rect 5538 639568 5594 639577
rect 5538 639503 5540 639512
rect 5592 639503 5594 639512
rect 5540 639474 5592 639480
rect 6276 639464 6328 639470
rect 6276 639406 6328 639412
rect 6182 639160 6238 639169
rect 6182 639095 6238 639104
rect 5448 610632 5500 610638
rect 5448 610574 5500 610580
rect 5356 553104 5408 553110
rect 5356 553046 5408 553052
rect 5264 496732 5316 496738
rect 5264 496674 5316 496680
rect 5172 380656 5224 380662
rect 5172 380598 5224 380604
rect 5080 323604 5132 323610
rect 5080 323546 5132 323552
rect 4988 237312 5040 237318
rect 4988 237254 5040 237260
rect 6196 194342 6224 639095
rect 6288 280158 6316 639406
rect 6380 337958 6408 640426
rect 6472 452470 6500 640562
rect 6564 510406 6592 640630
rect 7564 640416 7616 640422
rect 7564 640358 7616 640364
rect 6552 510400 6604 510406
rect 6552 510342 6604 510348
rect 6460 452464 6512 452470
rect 6460 452406 6512 452412
rect 6368 337952 6420 337958
rect 6368 337894 6420 337900
rect 7576 294438 7604 640358
rect 7668 366518 7696 641922
rect 7748 640552 7800 640558
rect 7748 640494 7800 640500
rect 7760 395486 7788 640494
rect 7840 639600 7892 639606
rect 7840 639542 7892 639548
rect 7852 438802 7880 639542
rect 7944 481166 7972 642058
rect 41602 641608 41658 641617
rect 41602 641543 41658 641552
rect 53102 641608 53158 641617
rect 53102 641543 53158 641552
rect 60922 641608 60978 641617
rect 60922 641543 60978 641552
rect 68466 641608 68522 641617
rect 68466 641543 68522 641552
rect 41616 640937 41644 641543
rect 53116 640937 53144 641543
rect 60936 640937 60964 641543
rect 68480 640937 68508 641543
rect 41602 640928 41658 640937
rect 8208 640892 8260 640898
rect 41602 640863 41658 640872
rect 53102 640928 53158 640937
rect 53102 640863 53158 640872
rect 60922 640928 60978 640937
rect 60922 640863 60978 640872
rect 68466 640928 68522 640937
rect 68466 640863 68522 640872
rect 8208 640834 8260 640840
rect 8116 640824 8168 640830
rect 8116 640766 8168 640772
rect 8024 640756 8076 640762
rect 8024 640698 8076 640704
rect 8036 567798 8064 640698
rect 8128 596086 8156 640766
rect 8220 624918 8248 640834
rect 23386 639568 23442 639577
rect 23308 639538 23386 639554
rect 23296 639532 23386 639538
rect 23348 639526 23386 639532
rect 23386 639503 23442 639512
rect 23296 639474 23348 639480
rect 50802 639432 50858 639441
rect 51078 639432 51134 639441
rect 50858 639390 51078 639418
rect 50802 639367 50858 639376
rect 51078 639367 51134 639376
rect 60646 639432 60702 639441
rect 60646 639367 60702 639376
rect 70122 639432 70178 639441
rect 70398 639432 70454 639441
rect 70178 639390 70398 639418
rect 70122 639367 70178 639376
rect 70398 639367 70454 639376
rect 60660 639266 60688 639367
rect 66166 639296 66222 639305
rect 60648 639260 60700 639266
rect 66166 639231 66168 639240
rect 60648 639202 60700 639208
rect 66220 639231 66222 639240
rect 66168 639202 66220 639208
rect 8208 624912 8260 624918
rect 8208 624854 8260 624860
rect 8116 596080 8168 596086
rect 8116 596022 8168 596028
rect 8024 567792 8076 567798
rect 8024 567734 8076 567740
rect 7932 481160 7984 481166
rect 7932 481102 7984 481108
rect 7840 438796 7892 438802
rect 7840 438738 7892 438744
rect 7748 395480 7800 395486
rect 7748 395422 7800 395428
rect 7656 366512 7708 366518
rect 7656 366454 7708 366460
rect 71044 338088 71096 338094
rect 71044 338030 71096 338036
rect 66904 338020 66956 338026
rect 66904 337962 66956 337968
rect 57244 337952 57296 337958
rect 57244 337894 57296 337900
rect 50344 337884 50396 337890
rect 50344 337826 50396 337832
rect 46204 337816 46256 337822
rect 46204 337758 46256 337764
rect 39304 337748 39356 337754
rect 39304 337690 39356 337696
rect 32404 337680 32456 337686
rect 32404 337622 32456 337628
rect 28264 337612 28316 337618
rect 28264 337554 28316 337560
rect 17224 337544 17276 337550
rect 17224 337486 17276 337492
rect 15844 337408 15896 337414
rect 10322 337376 10378 337385
rect 15844 337350 15896 337356
rect 10322 337311 10378 337320
rect 7564 294432 7616 294438
rect 7564 294374 7616 294380
rect 6276 280152 6328 280158
rect 6276 280094 6328 280100
rect 6184 194336 6236 194342
rect 6184 194278 6236 194284
rect 4896 179512 4948 179518
rect 4896 179454 4948 179460
rect 4804 79892 4856 79898
rect 4804 79834 4856 79840
rect 8852 7676 8904 7682
rect 8852 7618 8904 7624
rect 4122 7126 4200 7154
rect 4066 7103 4122 7112
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 3988 598 4108 626
rect 4080 480 4108 598
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8864 480 8892 7618
rect 10336 3466 10364 337311
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11244 3324 11296 3330
rect 11244 3266 11296 3272
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10060 480 10088 2994
rect 11256 480 11284 3266
rect 12452 480 12480 5034
rect 13648 480 13676 11698
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14844 480 14872 3470
rect 15856 3058 15884 337350
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 16040 480 16068 3402
rect 17236 3330 17264 337486
rect 24124 337476 24176 337482
rect 24124 337418 24176 337424
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 19248 13116 19300 13122
rect 19248 13058 19300 13064
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17224 3324 17276 3330
rect 17224 3266 17276 3272
rect 17328 1034 17356 5102
rect 19260 3602 19288 13058
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 17236 1006 17356 1034
rect 17236 480 17264 1006
rect 18340 480 18368 3538
rect 19536 480 19564 3538
rect 20720 3324 20772 3330
rect 20720 3266 20772 3272
rect 20732 480 20760 3266
rect 21928 480 21956 5170
rect 23400 3482 23428 14418
rect 24136 3602 24164 337418
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 25504 3664 25556 3670
rect 25504 3606 25556 3612
rect 24124 3596 24176 3602
rect 24124 3538 24176 3544
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 23124 3454 23428 3482
rect 23124 480 23152 3454
rect 24320 480 24348 3538
rect 25516 480 25544 3606
rect 26712 480 26740 7686
rect 28276 3330 28304 337554
rect 28908 15972 28960 15978
rect 28908 15914 28960 15920
rect 28264 3324 28316 3330
rect 28264 3266 28316 3272
rect 28920 3194 28948 15914
rect 31668 15904 31720 15910
rect 31668 15846 31720 15852
rect 30288 7812 30340 7818
rect 30288 7754 30340 7760
rect 27896 3188 27948 3194
rect 27896 3130 27948 3136
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 27908 480 27936 3130
rect 29104 480 29132 3130
rect 30300 480 30328 7754
rect 31680 626 31708 15846
rect 32416 3194 32444 337622
rect 37372 7948 37424 7954
rect 37372 7890 37424 7896
rect 33876 7880 33928 7886
rect 33876 7822 33928 7828
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 32404 3188 32456 3194
rect 32404 3130 32456 3136
rect 31496 598 31708 626
rect 31496 480 31524 598
rect 32692 480 32720 3674
rect 33888 480 33916 7822
rect 34980 4004 35032 4010
rect 34980 3946 35032 3952
rect 34992 480 35020 3946
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36188 480 36216 3334
rect 37384 480 37412 7890
rect 38568 3800 38620 3806
rect 38568 3742 38620 3748
rect 38580 480 38608 3742
rect 39316 3398 39344 337690
rect 44548 8084 44600 8090
rect 44548 8026 44600 8032
rect 40960 8016 41012 8022
rect 40960 7958 41012 7964
rect 39764 3868 39816 3874
rect 39764 3810 39816 3816
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 39776 480 39804 3810
rect 40972 480 41000 7958
rect 42156 4140 42208 4146
rect 42156 4082 42208 4088
rect 42168 480 42196 4082
rect 43352 3256 43404 3262
rect 43352 3198 43404 3204
rect 43364 480 43392 3198
rect 44560 480 44588 8026
rect 46216 4010 46244 337758
rect 49332 8152 49384 8158
rect 49332 8094 49384 8100
rect 48134 6216 48190 6225
rect 48134 6151 48190 6160
rect 46204 4004 46256 4010
rect 46204 3946 46256 3952
rect 46940 4004 46992 4010
rect 46940 3946 46992 3952
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45756 480 45784 3878
rect 46952 480 46980 3946
rect 48148 480 48176 6151
rect 49344 480 49372 8094
rect 50356 4146 50384 337826
rect 56416 8288 56468 8294
rect 56416 8230 56468 8236
rect 52828 8220 52880 8226
rect 52828 8162 52880 8168
rect 51632 6180 51684 6186
rect 51632 6122 51684 6128
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 50528 4072 50580 4078
rect 50528 4014 50580 4020
rect 50540 480 50568 4014
rect 51644 480 51672 6122
rect 52840 480 52868 8162
rect 55220 6248 55272 6254
rect 55220 6190 55272 6196
rect 54024 3324 54076 3330
rect 54024 3266 54076 3272
rect 54036 480 54064 3266
rect 55232 480 55260 6190
rect 56428 480 56456 8230
rect 57256 3330 57284 337894
rect 61384 337340 61436 337346
rect 61384 337282 61436 337288
rect 60646 10296 60702 10305
rect 60646 10231 60702 10240
rect 58808 6316 58860 6322
rect 58808 6258 58860 6264
rect 57612 4140 57664 4146
rect 57612 4082 57664 4088
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57624 480 57652 4082
rect 58820 480 58848 6258
rect 60660 3398 60688 10231
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60016 480 60044 3334
rect 61396 3330 61424 337282
rect 64788 10328 64840 10334
rect 64788 10270 64840 10276
rect 62396 6452 62448 6458
rect 62396 6394 62448 6400
rect 61384 3324 61436 3330
rect 61384 3266 61436 3272
rect 61200 3188 61252 3194
rect 61200 3130 61252 3136
rect 61212 480 61240 3130
rect 62408 480 62436 6394
rect 64800 3398 64828 10270
rect 65984 6384 66036 6390
rect 65984 6326 66036 6332
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 63604 480 63632 3334
rect 64788 3256 64840 3262
rect 64788 3198 64840 3204
rect 64800 480 64828 3198
rect 65996 480 66024 6326
rect 66916 3194 66944 337962
rect 69480 6520 69532 6526
rect 69480 6462 69532 6468
rect 67180 5296 67232 5302
rect 67180 5238 67232 5244
rect 66904 3188 66956 3194
rect 66904 3130 66956 3136
rect 67192 480 67220 5238
rect 68284 3052 68336 3058
rect 68284 2994 68336 3000
rect 68296 480 68324 2994
rect 69492 480 69520 6462
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 70688 480 70716 3334
rect 71056 3058 71084 338030
rect 72436 35902 72464 642087
rect 79966 639432 80022 639441
rect 80150 639432 80206 639441
rect 80022 639390 80150 639418
rect 79966 639367 80022 639376
rect 80150 639367 80206 639376
rect 86236 539578 86264 642262
rect 91742 641608 91798 641617
rect 91742 641543 91798 641552
rect 99562 641608 99618 641617
rect 99562 641543 99618 641552
rect 118882 641608 118938 641617
rect 118882 641543 118938 641552
rect 130382 641608 130438 641617
rect 130382 641543 130438 641552
rect 146114 641608 146170 641617
rect 146114 641543 146170 641552
rect 157522 641608 157578 641617
rect 157522 641543 157578 641552
rect 176842 641608 176898 641617
rect 176842 641543 176898 641552
rect 188342 641608 188398 641617
rect 188342 641543 188398 641552
rect 193954 641608 194010 641617
rect 193954 641543 194010 641552
rect 207662 641608 207718 641617
rect 207662 641543 207718 641552
rect 91756 640937 91784 641543
rect 99576 640937 99604 641543
rect 118896 640937 118924 641543
rect 130396 640937 130424 641543
rect 146128 640937 146156 641543
rect 157536 640937 157564 641543
rect 176856 640937 176884 641543
rect 188356 640937 188384 641543
rect 193968 640937 193996 641543
rect 207676 640937 207704 641543
rect 91742 640928 91798 640937
rect 91742 640863 91798 640872
rect 99562 640928 99618 640937
rect 99562 640863 99618 640872
rect 118882 640928 118938 640937
rect 118882 640863 118938 640872
rect 130382 640928 130438 640937
rect 130382 640863 130438 640872
rect 146114 640928 146170 640937
rect 146114 640863 146170 640872
rect 157522 640928 157578 640937
rect 157522 640863 157578 640872
rect 176842 640928 176898 640937
rect 176842 640863 176898 640872
rect 188342 640928 188398 640937
rect 188342 640863 188398 640872
rect 193954 640928 194010 640937
rect 193954 640863 194010 640872
rect 207662 640928 207718 640937
rect 207662 640863 207718 640872
rect 229744 640008 229796 640014
rect 231398 639976 231454 639985
rect 229744 639950 229796 639956
rect 220912 639940 220964 639946
rect 220912 639882 220964 639888
rect 109682 639840 109738 639849
rect 109682 639775 109738 639784
rect 119342 639840 119398 639849
rect 119342 639775 119398 639784
rect 162858 639840 162914 639849
rect 162858 639775 162914 639784
rect 177302 639840 177358 639849
rect 177302 639775 177358 639784
rect 89442 639432 89498 639441
rect 89718 639432 89774 639441
rect 89498 639390 89718 639418
rect 89442 639367 89498 639376
rect 89718 639367 89774 639376
rect 109696 639305 109724 639775
rect 119356 639441 119384 639775
rect 147770 639568 147826 639577
rect 147600 639526 147770 639554
rect 147600 639441 147628 639526
rect 147770 639503 147826 639512
rect 156326 639568 156382 639577
rect 156326 639503 156328 639512
rect 156380 639503 156382 639512
rect 162676 639532 162728 639538
rect 156328 639474 156380 639480
rect 162676 639474 162728 639480
rect 119342 639432 119398 639441
rect 119342 639367 119398 639376
rect 147586 639432 147642 639441
rect 162688 639418 162716 639474
rect 162872 639418 162900 639775
rect 177316 639441 177344 639775
rect 186318 639568 186374 639577
rect 220818 639568 220874 639577
rect 186318 639503 186374 639512
rect 201500 639532 201552 639538
rect 162688 639390 162900 639418
rect 177302 639432 177358 639441
rect 147586 639367 147642 639376
rect 177302 639367 177358 639376
rect 186042 639432 186098 639441
rect 186332 639418 186360 639503
rect 201500 639474 201552 639480
rect 211068 639532 211120 639538
rect 220818 639503 220874 639512
rect 211068 639474 211120 639480
rect 201512 639441 201540 639474
rect 186098 639390 186360 639418
rect 201498 639432 201554 639441
rect 186042 639367 186098 639376
rect 201498 639367 201554 639376
rect 211080 639305 211108 639474
rect 220832 639418 220860 639503
rect 220924 639418 220952 639882
rect 220832 639390 220952 639418
rect 109682 639296 109738 639305
rect 109682 639231 109738 639240
rect 211066 639296 211122 639305
rect 211066 639231 211122 639240
rect 86224 539572 86276 539578
rect 86224 539514 86276 539520
rect 228180 337544 228232 337550
rect 228180 337486 228232 337492
rect 228192 337414 228220 337486
rect 228180 337408 228232 337414
rect 228180 337350 228232 337356
rect 84844 337272 84896 337278
rect 84844 337214 84896 337220
rect 72424 35896 72476 35902
rect 72424 35838 72476 35844
rect 82728 14748 82780 14754
rect 82728 14690 82780 14696
rect 78588 14680 78640 14686
rect 78588 14622 78640 14628
rect 74448 14612 74500 14618
rect 74448 14554 74500 14560
rect 71688 14544 71740 14550
rect 71688 14486 71740 14492
rect 71700 3398 71728 14486
rect 73068 6588 73120 6594
rect 73068 6530 73120 6536
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 71872 3324 71924 3330
rect 71872 3266 71924 3272
rect 71044 3052 71096 3058
rect 71044 2994 71096 3000
rect 71884 480 71912 3266
rect 73080 480 73108 6530
rect 74460 3380 74488 14554
rect 76656 6656 76708 6662
rect 76656 6598 76708 6604
rect 74276 3352 74488 3380
rect 74276 480 74304 3352
rect 75460 2916 75512 2922
rect 75460 2858 75512 2864
rect 75472 480 75500 2858
rect 76668 480 76696 6598
rect 78600 3262 78628 14622
rect 80244 6724 80296 6730
rect 80244 6666 80296 6672
rect 77852 3256 77904 3262
rect 77852 3198 77904 3204
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 77864 480 77892 3198
rect 79048 2984 79100 2990
rect 79048 2926 79100 2932
rect 79060 480 79088 2926
rect 80256 480 80284 6666
rect 82740 3262 82768 14690
rect 83832 6792 83884 6798
rect 83832 6734 83884 6740
rect 81440 3256 81492 3262
rect 81440 3198 81492 3204
rect 82728 3256 82780 3262
rect 82728 3198 82780 3204
rect 81452 480 81480 3198
rect 82636 3188 82688 3194
rect 82636 3130 82688 3136
rect 82648 480 82676 3130
rect 83844 480 83872 6734
rect 84856 3262 84884 337214
rect 97264 337204 97316 337210
rect 97264 337146 97316 337152
rect 96528 15020 96580 15026
rect 96528 14962 96580 14968
rect 92388 14952 92440 14958
rect 92388 14894 92440 14900
rect 89628 14884 89680 14890
rect 89628 14826 89680 14832
rect 85488 14816 85540 14822
rect 85488 14758 85540 14764
rect 85500 3262 85528 14758
rect 87328 7540 87380 7546
rect 87328 7482 87380 7488
rect 84844 3256 84896 3262
rect 84844 3198 84896 3204
rect 84936 3256 84988 3262
rect 84936 3198 84988 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 84948 480 84976 3198
rect 86132 2984 86184 2990
rect 86132 2926 86184 2932
rect 86144 480 86172 2926
rect 87340 480 87368 7482
rect 89640 3262 89668 14826
rect 90916 7472 90968 7478
rect 90916 7414 90968 7420
rect 88524 3256 88576 3262
rect 88524 3198 88576 3204
rect 89628 3256 89680 3262
rect 89628 3198 89680 3204
rect 88536 480 88564 3198
rect 89812 3188 89864 3194
rect 89812 3130 89864 3136
rect 89824 1578 89852 3130
rect 89732 1550 89852 1578
rect 89732 480 89760 1550
rect 90928 480 90956 7414
rect 92400 3482 92428 14894
rect 94504 7404 94556 7410
rect 94504 7346 94556 7352
rect 92124 3454 92428 3482
rect 92124 480 92152 3454
rect 93308 3052 93360 3058
rect 93308 2994 93360 3000
rect 93320 480 93348 2994
rect 94516 480 94544 7346
rect 96540 3126 96568 14962
rect 97276 3126 97304 337146
rect 104808 337136 104860 337142
rect 104808 337078 104860 337084
rect 103428 16040 103480 16046
rect 103428 15982 103480 15988
rect 99288 15088 99340 15094
rect 99288 15030 99340 15036
rect 99196 10396 99248 10402
rect 99196 10338 99248 10344
rect 99208 3126 99236 10338
rect 95700 3120 95752 3126
rect 95700 3062 95752 3068
rect 96528 3120 96580 3126
rect 96528 3062 96580 3068
rect 97264 3120 97316 3126
rect 97264 3062 97316 3068
rect 98092 3120 98144 3126
rect 98092 3062 98144 3068
rect 99196 3120 99248 3126
rect 99196 3062 99248 3068
rect 95712 480 95740 3062
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 96908 480 96936 2994
rect 98104 480 98132 3062
rect 99300 480 99328 15030
rect 101588 10464 101640 10470
rect 101588 10406 101640 10412
rect 100484 2916 100536 2922
rect 100484 2858 100536 2864
rect 100496 480 100524 2858
rect 101600 480 101628 10406
rect 103440 3126 103468 15982
rect 104820 3126 104848 337078
rect 111708 337068 111760 337074
rect 111708 337010 111760 337016
rect 105544 336864 105596 336870
rect 105544 336806 105596 336812
rect 105176 10532 105228 10538
rect 105176 10474 105228 10480
rect 102784 3120 102836 3126
rect 102784 3062 102836 3068
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 103980 3120 104032 3126
rect 103980 3062 104032 3068
rect 104808 3120 104860 3126
rect 104808 3062 104860 3068
rect 102796 480 102824 3062
rect 103992 480 104020 3062
rect 105188 480 105216 10474
rect 105556 2854 105584 336806
rect 106924 336796 106976 336802
rect 106924 336738 106976 336744
rect 106372 3120 106424 3126
rect 106372 3062 106424 3068
rect 105544 2848 105596 2854
rect 105544 2790 105596 2796
rect 106384 480 106412 3062
rect 106936 2990 106964 336738
rect 110328 16176 110380 16182
rect 110328 16118 110380 16124
rect 107568 16108 107620 16114
rect 107568 16050 107620 16056
rect 107580 3126 107608 16050
rect 108764 10600 108816 10606
rect 108764 10542 108816 10548
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 106924 2984 106976 2990
rect 106924 2926 106976 2932
rect 107568 2848 107620 2854
rect 107568 2790 107620 2796
rect 107580 480 107608 2790
rect 108776 480 108804 10542
rect 110340 3346 110368 16118
rect 109972 3318 110368 3346
rect 109972 480 110000 3318
rect 111720 3126 111748 337010
rect 118608 337000 118660 337006
rect 118608 336942 118660 336948
rect 114468 16244 114520 16250
rect 114468 16186 114520 16192
rect 113088 10668 113140 10674
rect 113088 10610 113140 10616
rect 111156 3120 111208 3126
rect 111156 3062 111208 3068
rect 111708 3120 111760 3126
rect 111708 3062 111760 3068
rect 111168 480 111196 3062
rect 113100 2990 113128 10610
rect 114480 2990 114508 16186
rect 117228 14136 117280 14142
rect 117228 14078 117280 14084
rect 117136 10736 117188 10742
rect 117136 10678 117188 10684
rect 117148 3618 117176 10678
rect 116964 3590 117176 3618
rect 116964 2990 116992 3590
rect 117240 3482 117268 14078
rect 117148 3454 117268 3482
rect 112352 2984 112404 2990
rect 112352 2926 112404 2932
rect 113088 2984 113140 2990
rect 113088 2926 113140 2932
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 115940 2984 115992 2990
rect 115940 2926 115992 2932
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 112364 480 112392 2926
rect 113560 480 113588 2926
rect 114744 2916 114796 2922
rect 114744 2858 114796 2864
rect 114756 480 114784 2858
rect 115952 480 115980 2926
rect 117148 480 117176 3454
rect 118620 3346 118648 336942
rect 125508 336932 125560 336938
rect 125508 336874 125560 336880
rect 125416 16380 125468 16386
rect 125416 16322 125468 16328
rect 121368 16312 121420 16318
rect 121368 16254 121420 16260
rect 119988 10804 120040 10810
rect 119988 10746 120040 10752
rect 118252 3318 118648 3346
rect 118252 480 118280 3318
rect 120000 2990 120028 10746
rect 121380 2990 121408 16254
rect 124128 10872 124180 10878
rect 124128 10814 124180 10820
rect 124140 3482 124168 10814
rect 125428 4214 125456 16322
rect 124220 4208 124272 4214
rect 124220 4150 124272 4156
rect 125416 4208 125468 4214
rect 125416 4150 125468 4156
rect 123036 3454 124168 3482
rect 119436 2984 119488 2990
rect 119436 2926 119488 2932
rect 119988 2984 120040 2990
rect 119988 2926 120040 2932
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 121368 2984 121420 2990
rect 121368 2926 121420 2932
rect 119448 480 119476 2926
rect 120644 480 120672 2926
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 121840 480 121868 2790
rect 123036 480 123064 3454
rect 124232 480 124260 4150
rect 125520 3482 125548 336874
rect 229100 335640 229152 335646
rect 229100 335582 229152 335588
rect 129648 15156 129700 15162
rect 129648 15098 129700 15104
rect 126888 11892 126940 11898
rect 126888 11834 126940 11840
rect 126900 3482 126928 11834
rect 128268 11824 128320 11830
rect 128268 11766 128320 11772
rect 128280 3482 128308 11766
rect 129660 3482 129688 15098
rect 160008 14408 160060 14414
rect 160008 14350 160060 14356
rect 157248 14340 157300 14346
rect 157248 14282 157300 14288
rect 155868 13660 155920 13666
rect 155868 13602 155920 13608
rect 153108 13592 153160 13598
rect 153108 13534 153160 13540
rect 148968 13524 149020 13530
rect 148968 13466 149020 13472
rect 146208 13320 146260 13326
rect 146208 13262 146260 13268
rect 144828 13252 144880 13258
rect 144828 13194 144880 13200
rect 132408 13184 132460 13190
rect 132408 13126 132460 13132
rect 130200 5364 130252 5370
rect 130200 5306 130252 5312
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 127820 3454 128308 3482
rect 129016 3454 129688 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3454
rect 129016 480 129044 3454
rect 130212 480 130240 5306
rect 132420 3482 132448 13126
rect 142068 11960 142120 11966
rect 142068 11902 142120 11908
rect 140688 10940 140740 10946
rect 140688 10882 140740 10888
rect 132592 8968 132644 8974
rect 132592 8910 132644 8916
rect 136086 8936 136142 8945
rect 131408 3454 132448 3482
rect 131408 480 131436 3454
rect 132604 480 132632 8910
rect 136086 8871 136142 8880
rect 134890 7576 134946 7585
rect 134890 7511 134946 7520
rect 133788 5432 133840 5438
rect 133788 5374 133840 5380
rect 133800 480 133828 5374
rect 134904 480 134932 7511
rect 136100 480 136128 8871
rect 138480 7336 138532 7342
rect 138480 7278 138532 7284
rect 137284 5500 137336 5506
rect 137284 5442 137336 5448
rect 137296 480 137324 5442
rect 138492 480 138520 7278
rect 140700 610 140728 10882
rect 141976 7268 142028 7274
rect 141976 7210 142028 7216
rect 140872 4208 140924 4214
rect 140872 4150 140924 4156
rect 139676 604 139728 610
rect 139676 546 139728 552
rect 140688 604 140740 610
rect 140688 546 140740 552
rect 139688 480 139716 546
rect 140884 480 140912 4150
rect 141988 3482 142016 7210
rect 142080 4214 142108 11902
rect 143448 11008 143500 11014
rect 143448 10950 143500 10956
rect 142068 4208 142120 4214
rect 142068 4150 142120 4156
rect 141988 3454 142108 3482
rect 142080 480 142108 3454
rect 143460 3346 143488 10950
rect 144840 3346 144868 13194
rect 146220 3346 146248 13262
rect 147588 10260 147640 10266
rect 147588 10202 147640 10208
rect 147600 3346 147628 10202
rect 148980 3346 149008 13466
rect 150348 13456 150400 13462
rect 150348 13398 150400 13404
rect 150360 3346 150388 13398
rect 151728 13388 151780 13394
rect 151728 13330 151780 13336
rect 151636 10192 151688 10198
rect 151636 10134 151688 10140
rect 151648 4214 151676 10134
rect 150440 4208 150492 4214
rect 150440 4150 150492 4156
rect 151636 4208 151688 4214
rect 151636 4150 151688 4156
rect 143276 3318 143488 3346
rect 144472 3318 144868 3346
rect 145668 3318 146248 3346
rect 146864 3318 147628 3346
rect 148060 3318 149008 3346
rect 149256 3318 150388 3346
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3318
rect 146864 480 146892 3318
rect 148060 480 148088 3318
rect 149256 480 149284 3318
rect 150452 480 150480 4150
rect 151740 3482 151768 13330
rect 151556 3454 151768 3482
rect 151556 480 151584 3454
rect 153120 3346 153148 13534
rect 154488 10124 154540 10130
rect 154488 10066 154540 10072
rect 154500 3346 154528 10066
rect 155880 3346 155908 13602
rect 157260 3346 157288 14282
rect 159916 13728 159968 13734
rect 159916 13670 159968 13676
rect 158628 10056 158680 10062
rect 158628 9998 158680 10004
rect 158640 3346 158668 9998
rect 159928 4214 159956 13670
rect 158720 4208 158772 4214
rect 158720 4150 158772 4156
rect 159916 4208 159968 4214
rect 159916 4150 159968 4156
rect 152752 3318 153148 3346
rect 153948 3318 154528 3346
rect 155144 3318 155908 3346
rect 156340 3318 157288 3346
rect 157536 3318 158668 3346
rect 152752 480 152780 3318
rect 153948 480 153976 3318
rect 155144 480 155172 3318
rect 156340 480 156368 3318
rect 157536 480 157564 3318
rect 158732 480 158760 4150
rect 160020 3482 160048 14350
rect 165528 14272 165580 14278
rect 165528 14214 165580 14220
rect 162768 12028 162820 12034
rect 162768 11970 162820 11976
rect 161388 9988 161440 9994
rect 161388 9930 161440 9936
rect 159928 3454 160048 3482
rect 159928 480 159956 3454
rect 161400 3346 161428 9930
rect 162780 3346 162808 11970
rect 163504 6860 163556 6866
rect 163504 6802 163556 6808
rect 161124 3318 161428 3346
rect 162320 3318 162808 3346
rect 161124 480 161152 3318
rect 162320 480 162348 3318
rect 163516 480 163544 6802
rect 165540 3346 165568 14214
rect 168288 14204 168340 14210
rect 168288 14146 168340 14152
rect 166908 12096 166960 12102
rect 166908 12038 166960 12044
rect 166920 3346 166948 12038
rect 167092 6112 167144 6118
rect 167092 6054 167144 6060
rect 164712 3318 165568 3346
rect 165908 3318 166948 3346
rect 164712 480 164740 3318
rect 165908 480 165936 3318
rect 167104 480 167132 6054
rect 168300 3482 168328 14146
rect 202788 13796 202840 13802
rect 202788 13738 202840 13744
rect 200028 13048 200080 13054
rect 200028 12990 200080 12996
rect 184848 12436 184900 12442
rect 184848 12378 184900 12384
rect 180708 12368 180760 12374
rect 180708 12310 180760 12316
rect 176568 12300 176620 12306
rect 176568 12242 176620 12248
rect 173808 12232 173860 12238
rect 173808 12174 173860 12180
rect 169668 12164 169720 12170
rect 169668 12106 169720 12112
rect 168208 3454 168328 3482
rect 168208 480 168236 3454
rect 169680 3346 169708 12106
rect 171784 9036 171836 9042
rect 171784 8978 171836 8984
rect 170588 6044 170640 6050
rect 170588 5986 170640 5992
rect 169404 3318 169708 3346
rect 169404 480 169432 3318
rect 170600 480 170628 5986
rect 171796 480 171824 8978
rect 173820 610 173848 12174
rect 175372 9104 175424 9110
rect 175372 9046 175424 9052
rect 174176 5976 174228 5982
rect 174176 5918 174228 5924
rect 172980 604 173032 610
rect 172980 546 173032 552
rect 173808 604 173860 610
rect 173808 546 173860 552
rect 172992 480 173020 546
rect 174188 480 174216 5918
rect 175384 480 175412 9046
rect 176580 480 176608 12242
rect 178960 9172 179012 9178
rect 178960 9114 179012 9120
rect 177764 5908 177816 5914
rect 177764 5850 177816 5856
rect 177776 480 177804 5850
rect 178972 480 179000 9114
rect 180720 610 180748 12310
rect 182548 9240 182600 9246
rect 182548 9182 182600 9188
rect 181352 5840 181404 5846
rect 181352 5782 181404 5788
rect 180156 604 180208 610
rect 180156 546 180208 552
rect 180708 604 180760 610
rect 180708 546 180760 552
rect 180168 480 180196 546
rect 181364 480 181392 5782
rect 182560 480 182588 9182
rect 184860 5930 184888 12378
rect 187608 11688 187660 11694
rect 187608 11630 187660 11636
rect 186044 9308 186096 9314
rect 186044 9250 186096 9256
rect 183756 5902 184888 5930
rect 183756 480 183784 5902
rect 184848 5772 184900 5778
rect 184848 5714 184900 5720
rect 184860 480 184888 5714
rect 186056 480 186084 9250
rect 187620 3482 187648 11630
rect 191748 11620 191800 11626
rect 191748 11562 191800 11568
rect 189632 9376 189684 9382
rect 189632 9318 189684 9324
rect 188436 5704 188488 5710
rect 188436 5646 188488 5652
rect 187252 3454 187648 3482
rect 187252 480 187280 3454
rect 188448 480 188476 5646
rect 189644 480 189672 9318
rect 191760 3482 191788 11562
rect 194508 11552 194560 11558
rect 194508 11494 194560 11500
rect 193220 9444 193272 9450
rect 193220 9386 193272 9392
rect 192024 5636 192076 5642
rect 192024 5578 192076 5584
rect 190840 3454 191788 3482
rect 190840 480 190868 3454
rect 192036 480 192064 5578
rect 193232 480 193260 9386
rect 194520 3482 194548 11494
rect 198648 11484 198700 11490
rect 198648 11426 198700 11432
rect 196808 9512 196860 9518
rect 196808 9454 196860 9460
rect 195612 5568 195664 5574
rect 195612 5510 195664 5516
rect 194428 3454 194548 3482
rect 194428 480 194456 3454
rect 195624 480 195652 5510
rect 196820 480 196848 9454
rect 198660 3482 198688 11426
rect 200040 3482 200068 12990
rect 201500 11416 201552 11422
rect 201500 11358 201552 11364
rect 200396 9580 200448 9586
rect 200396 9522 200448 9528
rect 198016 3454 198688 3482
rect 199212 3454 200068 3482
rect 198016 480 198044 3454
rect 199212 480 199240 3454
rect 200408 480 200436 9522
rect 201512 480 201540 11358
rect 202800 3482 202828 13738
rect 206928 12980 206980 12986
rect 206928 12922 206980 12928
rect 205548 11348 205600 11354
rect 205548 11290 205600 11296
rect 203892 9648 203944 9654
rect 203892 9590 203944 9596
rect 202708 3454 202828 3482
rect 202708 480 202736 3454
rect 203904 480 203932 9590
rect 205560 610 205588 11290
rect 206940 610 206968 12922
rect 213828 12912 213880 12918
rect 213828 12854 213880 12860
rect 211068 12844 211120 12850
rect 211068 12786 211120 12792
rect 210976 8900 211028 8906
rect 210976 8842 211028 8848
rect 207480 8832 207532 8838
rect 207480 8774 207532 8780
rect 205088 604 205140 610
rect 205088 546 205140 552
rect 205548 604 205600 610
rect 205548 546 205600 552
rect 206284 604 206336 610
rect 206284 546 206336 552
rect 206928 604 206980 610
rect 206928 546 206980 552
rect 205100 480 205128 546
rect 206296 480 206324 546
rect 207492 480 207520 8774
rect 208676 4548 208728 4554
rect 208676 4490 208728 4496
rect 208688 480 208716 4490
rect 209872 4208 209924 4214
rect 209872 4150 209924 4156
rect 209884 480 209912 4150
rect 210988 3482 211016 8842
rect 211080 4214 211108 12786
rect 212264 4480 212316 4486
rect 212264 4422 212316 4428
rect 211068 4208 211120 4214
rect 211068 4150 211120 4156
rect 210988 3454 211108 3482
rect 211080 480 211108 3454
rect 212276 480 212304 4422
rect 213840 3482 213868 12854
rect 217968 12776 218020 12782
rect 217968 12718 218020 12724
rect 214656 8764 214708 8770
rect 214656 8706 214708 8712
rect 213472 3454 213868 3482
rect 213472 480 213500 3454
rect 214668 480 214696 8706
rect 215852 4752 215904 4758
rect 215852 4694 215904 4700
rect 215864 480 215892 4694
rect 217980 3482 218008 12718
rect 220728 12708 220780 12714
rect 220728 12650 220780 12656
rect 218152 8628 218204 8634
rect 218152 8570 218204 8576
rect 217060 3454 218008 3482
rect 217060 480 217088 3454
rect 218164 480 218192 8570
rect 219346 4856 219402 4865
rect 219346 4791 219402 4800
rect 219360 480 219388 4791
rect 220740 610 220768 12650
rect 221740 8696 221792 8702
rect 221740 8638 221792 8644
rect 220544 604 220596 610
rect 220544 546 220596 552
rect 220728 604 220780 610
rect 220728 546 220780 552
rect 220556 480 220584 546
rect 221752 480 221780 8638
rect 225328 8560 225380 8566
rect 225328 8502 225380 8508
rect 224132 7200 224184 7206
rect 224132 7142 224184 7148
rect 222936 4684 222988 4690
rect 222936 4626 222988 4632
rect 222948 480 222976 4626
rect 224144 480 224172 7142
rect 225340 480 225368 8502
rect 228916 8492 228968 8498
rect 228916 8434 228968 8440
rect 227720 7132 227772 7138
rect 227720 7074 227772 7080
rect 226524 4616 226576 4622
rect 226524 4558 226576 4564
rect 226536 480 226564 4558
rect 227732 480 227760 7074
rect 228928 480 228956 8434
rect 229112 4894 229140 335582
rect 229756 266354 229784 639950
rect 231058 639934 231398 639962
rect 236288 639948 236316 642534
rect 252008 642456 252060 642462
rect 252008 642398 252060 642404
rect 241518 642288 241574 642297
rect 241518 642223 241574 642232
rect 238852 640960 238904 640966
rect 238852 640902 238904 640908
rect 238864 639948 238892 640902
rect 241532 639948 241560 642223
rect 243542 641608 243598 641617
rect 243542 641543 243598 641552
rect 243556 640937 243584 641543
rect 246764 641096 246816 641102
rect 246764 641038 246816 641044
rect 243542 640928 243598 640937
rect 243542 640863 243598 640872
rect 244186 640112 244242 640121
rect 244186 640047 244242 640056
rect 244200 639948 244228 640047
rect 246776 639948 246804 641038
rect 252020 639948 252048 642398
rect 257344 642388 257396 642394
rect 257344 642330 257396 642336
rect 257356 639948 257384 642330
rect 258736 641034 258764 642767
rect 258724 641028 258776 641034
rect 258724 640970 258776 640976
rect 259932 639948 259960 642903
rect 265164 642864 265216 642870
rect 265164 642806 265216 642812
rect 263600 642456 263652 642462
rect 263600 642398 263652 642404
rect 262588 641164 262640 641170
rect 262588 641106 262640 641112
rect 262600 639948 262628 641106
rect 263612 639946 263640 642398
rect 265176 639948 265204 642806
rect 269040 642666 269068 670686
rect 300780 643958 300808 699654
rect 344928 696992 344980 696998
rect 344928 696934 344980 696940
rect 342168 673532 342220 673538
rect 342168 673474 342220 673480
rect 336648 650072 336700 650078
rect 336648 650014 336700 650020
rect 300768 643952 300820 643958
rect 300768 643894 300820 643900
rect 283656 643068 283708 643074
rect 283656 643010 283708 643016
rect 267832 642660 267884 642666
rect 267832 642602 267884 642608
rect 269028 642660 269080 642666
rect 269028 642602 269080 642608
rect 267844 639948 267872 642602
rect 270500 642524 270552 642530
rect 270500 642466 270552 642472
rect 270512 639948 270540 642466
rect 278320 642456 278372 642462
rect 278320 642398 278372 642404
rect 275282 641608 275338 641617
rect 275282 641543 275338 641552
rect 275296 640937 275324 641543
rect 275744 641232 275796 641238
rect 275744 641174 275796 641180
rect 275282 640928 275338 640937
rect 275282 640863 275338 640872
rect 275756 639948 275784 641174
rect 278332 639948 278360 642398
rect 283668 639948 283696 643010
rect 307300 643000 307352 643006
rect 307300 642942 307352 642948
rect 325698 642968 325754 642977
rect 288900 642728 288952 642734
rect 288900 642670 288952 642676
rect 286232 641300 286284 641306
rect 286232 641242 286284 641248
rect 286244 639948 286272 641242
rect 288912 639948 288940 642670
rect 304632 642660 304684 642666
rect 304632 642602 304684 642608
rect 290004 642592 290056 642598
rect 290004 642534 290056 642540
rect 294144 642592 294196 642598
rect 294144 642534 294196 642540
rect 231398 639911 231454 639920
rect 235264 639940 235316 639946
rect 235264 639882 235316 639888
rect 263600 639940 263652 639946
rect 263600 639882 263652 639888
rect 235276 639849 235304 639882
rect 281264 639872 281316 639878
rect 233974 639840 234030 639849
rect 233634 639798 233974 639826
rect 233974 639775 234030 639784
rect 235262 639840 235318 639849
rect 249522 639840 249578 639849
rect 249458 639798 249522 639826
rect 235262 639775 235318 639784
rect 254950 639840 255006 639849
rect 254702 639798 254950 639826
rect 249522 639775 249578 639784
rect 273102 639810 273208 639826
rect 281014 639820 281264 639826
rect 290016 639849 290044 642534
rect 291476 641028 291528 641034
rect 291476 640970 291528 640976
rect 291488 639948 291516 640970
rect 294156 639948 294184 642534
rect 299388 641368 299440 641374
rect 299388 641310 299440 641316
rect 296812 640144 296864 640150
rect 296812 640086 296864 640092
rect 296824 639948 296852 640086
rect 299400 639948 299428 641310
rect 302054 640112 302110 640121
rect 302054 640047 302110 640056
rect 302068 639948 302096 640047
rect 304644 639948 304672 642602
rect 307312 639948 307340 642942
rect 325698 642903 325754 642912
rect 331036 642932 331088 642938
rect 320824 642864 320876 642870
rect 320824 642806 320876 642812
rect 323124 642864 323176 642870
rect 323124 642806 323176 642812
rect 320456 642796 320508 642802
rect 320456 642738 320508 642744
rect 307668 642728 307720 642734
rect 307668 642670 307720 642676
rect 315212 642728 315264 642734
rect 315212 642670 315264 642676
rect 307680 640218 307708 642670
rect 312544 641504 312596 641510
rect 312544 641446 312596 641452
rect 309968 641436 310020 641442
rect 309968 641378 310020 641384
rect 307668 640212 307720 640218
rect 307668 640154 307720 640160
rect 309980 639948 310008 641378
rect 312556 639948 312584 641446
rect 315224 639948 315252 642670
rect 317788 641572 317840 641578
rect 317788 641514 317840 641520
rect 317800 639948 317828 641514
rect 320468 639948 320496 642738
rect 320836 640286 320864 642806
rect 320824 640280 320876 640286
rect 320824 640222 320876 640228
rect 323136 639948 323164 642806
rect 325712 639948 325740 642903
rect 331036 642874 331088 642880
rect 328182 639976 328238 639985
rect 328238 639934 328394 639962
rect 331048 639948 331076 642874
rect 333612 641640 333664 641646
rect 333612 641582 333664 641588
rect 333624 639948 333652 641582
rect 336660 639962 336688 650014
rect 339224 640076 339276 640082
rect 339224 640018 339276 640024
rect 339236 639962 339264 640018
rect 342180 639962 342208 673474
rect 344940 639962 344968 696934
rect 347688 685908 347740 685914
rect 347688 685850 347740 685856
rect 347700 640098 347728 685850
rect 349436 643748 349488 643754
rect 349436 643690 349488 643696
rect 336306 639934 336688 639962
rect 338882 639934 339264 639962
rect 341996 639934 342208 639962
rect 344756 639934 344968 639962
rect 347332 640070 347728 640098
rect 328182 639911 328238 639920
rect 281014 639814 281316 639820
rect 290002 639840 290058 639849
rect 273102 639804 273220 639810
rect 273102 639798 273168 639804
rect 254950 639775 255006 639784
rect 281014 639798 281304 639814
rect 290002 639775 290058 639784
rect 340786 639840 340842 639849
rect 340970 639840 341026 639849
rect 340842 639798 340970 639826
rect 340786 639775 340842 639784
rect 341996 639826 342024 639934
rect 344756 639826 344784 639934
rect 347332 639826 347360 640070
rect 349448 639948 349476 643690
rect 353220 640098 353248 700198
rect 355980 640098 356008 700878
rect 362868 700120 362920 700126
rect 362868 700062 362920 700068
rect 360108 700052 360160 700058
rect 360108 699994 360160 700000
rect 357348 643884 357400 643890
rect 357348 643826 357400 643832
rect 352576 640070 353248 640098
rect 355336 640070 356008 640098
rect 352576 639962 352604 640070
rect 355336 639962 355364 640070
rect 352038 639934 352604 639962
rect 354706 639934 355364 639962
rect 357360 639948 357388 643826
rect 360120 639962 360148 699994
rect 362880 639962 362908 700062
rect 364996 699718 365024 703520
rect 393320 701004 393372 701010
rect 393320 700946 393372 700952
rect 390560 700868 390612 700874
rect 390560 700810 390612 700816
rect 383660 700188 383712 700194
rect 383660 700130 383712 700136
rect 375380 699916 375432 699922
rect 375380 699858 375432 699864
rect 371148 699848 371200 699854
rect 371148 699790 371200 699796
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 365628 699712 365680 699718
rect 365628 699654 365680 699660
rect 368388 699712 368440 699718
rect 368388 699654 368440 699660
rect 365168 644020 365220 644026
rect 365168 643962 365220 643968
rect 359950 639934 360148 639962
rect 362618 639934 362908 639962
rect 365180 639948 365208 643962
rect 365640 643142 365668 699654
rect 365628 643136 365680 643142
rect 365628 643078 365680 643084
rect 368400 639826 368428 699654
rect 371160 639826 371188 699790
rect 373080 643136 373132 643142
rect 373080 643078 373132 643084
rect 373092 639948 373120 643078
rect 375392 639962 375420 699858
rect 378140 699780 378192 699786
rect 378140 699722 378192 699728
rect 378152 639962 378180 699722
rect 380992 643952 381044 643958
rect 380992 643894 381044 643900
rect 375392 639934 375774 639962
rect 378152 639934 378350 639962
rect 381004 639948 381032 643894
rect 383672 639948 383700 700130
rect 385040 699984 385092 699990
rect 385040 699926 385092 699932
rect 385052 640098 385080 699926
rect 388904 643816 388956 643822
rect 388904 643758 388956 643764
rect 385052 640070 385724 640098
rect 341550 639798 342024 639826
rect 344218 639798 344784 639826
rect 346794 639798 347360 639826
rect 367862 639798 368428 639826
rect 370530 639798 371188 639826
rect 385696 639826 385724 640070
rect 388916 639948 388944 643758
rect 390572 640098 390600 700810
rect 390572 640070 391244 640098
rect 391216 639962 391244 640070
rect 391216 639934 391506 639962
rect 393332 639826 393360 700946
rect 396080 700800 396132 700806
rect 396080 700742 396132 700748
rect 396092 639826 396120 700742
rect 397472 699718 397500 703520
rect 401600 700732 401652 700738
rect 401600 700674 401652 700680
rect 398840 700664 398892 700670
rect 398840 700606 398892 700612
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 398852 639826 398880 700606
rect 401612 639962 401640 700674
rect 404360 700596 404412 700602
rect 404360 700538 404412 700544
rect 404372 639962 404400 700538
rect 409880 700528 409932 700534
rect 409880 700470 409932 700476
rect 407120 700460 407172 700466
rect 407120 700402 407172 700408
rect 407132 639962 407160 700402
rect 409892 639962 409920 700470
rect 411260 700392 411312 700398
rect 411260 700334 411312 700340
rect 411272 645182 411300 700334
rect 413664 699854 413692 703520
rect 414018 700360 414074 700369
rect 414018 700295 414074 700304
rect 416780 700324 416832 700330
rect 413652 699848 413704 699854
rect 413652 699790 413704 699796
rect 411260 645176 411312 645182
rect 411260 645118 411312 645124
rect 412548 645176 412600 645182
rect 412548 645118 412600 645124
rect 401612 639934 402086 639962
rect 404372 639934 404662 639962
rect 407132 639934 407330 639962
rect 409892 639934 409998 639962
rect 412560 639948 412588 645118
rect 414032 639826 414060 700295
rect 416780 700266 416832 700272
rect 416792 639826 416820 700266
rect 429856 688634 429884 703520
rect 462332 700058 462360 703520
rect 478524 700126 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700120 478564 700126
rect 478512 700062 478564 700068
rect 462320 700052 462372 700058
rect 462320 699994 462372 700000
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 429396 685930 429424 688570
rect 494900 686089 494928 703446
rect 527192 700262 527220 703520
rect 543476 700942 543504 703520
rect 543464 700936 543516 700942
rect 543464 700878 543516 700884
rect 527180 700256 527232 700262
rect 527180 700198 527232 700204
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 429304 685902 429424 685930
rect 494242 685944 494298 685953
rect 429304 684486 429332 685902
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 419540 681760 419592 681766
rect 419540 681702 419592 681708
rect 419552 640098 419580 681702
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 577504 670744 577556 670750
rect 577504 670686 577556 670692
rect 425060 667956 425112 667962
rect 425060 667898 425112 667904
rect 422300 652792 422352 652798
rect 422300 652734 422352 652740
rect 422312 640234 422340 652734
rect 425072 640234 425100 667898
rect 429476 666596 429528 666602
rect 429476 666538 429528 666544
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 429488 659682 429516 666538
rect 429304 659654 429516 659682
rect 494164 659682 494192 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 429304 656878 429332 659654
rect 429292 656872 429344 656878
rect 429292 656814 429344 656820
rect 494256 654158 494284 659654
rect 559208 659654 559420 659682
rect 559208 656878 559236 659654
rect 559196 656872 559248 656878
rect 559196 656814 559248 656820
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 429200 647284 429252 647290
rect 429200 647226 429252 647232
rect 429212 644026 429240 647226
rect 429200 644020 429252 644026
rect 429200 643962 429252 643968
rect 494072 643890 494100 654094
rect 559288 647284 559340 647290
rect 559288 647226 559340 647232
rect 494060 643884 494112 643890
rect 494060 643826 494112 643832
rect 559300 643754 559328 647226
rect 559288 643748 559340 643754
rect 559288 643690 559340 643696
rect 520462 643104 520518 643113
rect 427820 643068 427872 643074
rect 427820 643010 427872 643016
rect 429016 643068 429068 643074
rect 520462 643039 520518 643048
rect 523132 643068 523184 643074
rect 429016 643010 429068 643016
rect 427832 641714 427860 643010
rect 429028 642161 429056 643010
rect 473360 643000 473412 643006
rect 473360 642942 473412 642948
rect 438860 642320 438912 642326
rect 438860 642262 438912 642268
rect 438952 642320 439004 642326
rect 438952 642262 439004 642268
rect 454684 642320 454736 642326
rect 454684 642262 454736 642268
rect 433616 642252 433668 642258
rect 433616 642194 433668 642200
rect 429014 642152 429070 642161
rect 429014 642087 429070 642096
rect 427820 641708 427872 641714
rect 427820 641650 427872 641656
rect 428372 640892 428424 640898
rect 428372 640834 428424 640840
rect 422312 640206 422800 640234
rect 425072 640206 425376 640234
rect 419552 640070 420132 640098
rect 420104 639962 420132 640070
rect 422772 639962 422800 640206
rect 425348 639962 425376 640206
rect 420104 639934 420486 639962
rect 422772 639934 423154 639962
rect 425348 639934 425730 639962
rect 428384 639948 428412 640834
rect 431040 640824 431092 640830
rect 431040 640766 431092 640772
rect 431052 639948 431080 640766
rect 433628 639948 433656 642194
rect 436284 640756 436336 640762
rect 436284 640698 436336 640704
rect 436296 639948 436324 640698
rect 438872 639948 438900 642262
rect 385696 639798 386262 639826
rect 393332 639798 394174 639826
rect 396092 639798 396842 639826
rect 398852 639798 399418 639826
rect 414032 639798 415242 639826
rect 416792 639798 417818 639826
rect 340970 639775 341026 639784
rect 273168 639746 273220 639752
rect 438964 639742 438992 642262
rect 441528 642184 441580 642190
rect 441528 642126 441580 642132
rect 441540 639948 441568 642126
rect 446772 642116 446824 642122
rect 446772 642058 446824 642064
rect 446864 642116 446916 642122
rect 446864 642058 446916 642064
rect 444196 640824 444248 640830
rect 444196 640766 444248 640772
rect 444208 639948 444236 640766
rect 446784 639948 446812 642058
rect 438952 639736 439004 639742
rect 340786 639704 340842 639713
rect 340970 639704 341026 639713
rect 340842 639662 340970 639690
rect 340786 639639 340842 639648
rect 438952 639678 439004 639684
rect 446876 639674 446904 642058
rect 449440 642048 449492 642054
rect 449440 641990 449492 641996
rect 449452 639948 449480 641990
rect 452016 640620 452068 640626
rect 452016 640562 452068 640568
rect 452028 639948 452056 640562
rect 454696 639948 454724 642262
rect 462596 641980 462648 641986
rect 462596 641922 462648 641928
rect 462964 641980 463016 641986
rect 462964 641922 463016 641928
rect 459928 640552 459980 640558
rect 459928 640494 459980 640500
rect 459940 639948 459968 640494
rect 462608 639948 462636 641922
rect 457076 639736 457128 639742
rect 462976 639713 463004 641922
rect 465172 641912 465224 641918
rect 465172 641854 465224 641860
rect 463422 640112 463478 640121
rect 463422 640047 463478 640056
rect 463238 639976 463294 639985
rect 463238 639911 463294 639920
rect 463252 639713 463280 639911
rect 463436 639713 463464 640047
rect 465184 639948 465212 641854
rect 473084 641844 473136 641850
rect 473084 641786 473136 641792
rect 467840 640484 467892 640490
rect 467840 640426 467892 640432
rect 467852 639948 467880 640426
rect 471058 639976 471114 639985
rect 473096 639948 473124 641786
rect 473372 640898 473400 642942
rect 504638 642832 504694 642841
rect 504638 642767 504694 642776
rect 483662 642696 483718 642705
rect 483662 642631 483718 642640
rect 473360 640892 473412 640898
rect 473360 640834 473412 640840
rect 475752 640416 475804 640422
rect 475752 640358 475804 640364
rect 475764 639948 475792 640358
rect 478052 640008 478104 640014
rect 478104 639956 478354 639962
rect 478052 639950 478354 639956
rect 478064 639934 478354 639950
rect 483676 639948 483704 642631
rect 491482 642560 491538 642569
rect 491482 642495 491538 642504
rect 486240 642116 486292 642122
rect 486240 642058 486292 642064
rect 485136 641844 485188 641850
rect 485136 641786 485188 641792
rect 471058 639911 471114 639920
rect 471072 639713 471100 639911
rect 485148 639713 485176 641786
rect 486252 639948 486280 642058
rect 488908 641776 488960 641782
rect 488908 641718 488960 641724
rect 488920 639948 488948 641718
rect 491496 639948 491524 642495
rect 499394 642424 499450 642433
rect 499394 642359 499450 642368
rect 494150 642016 494206 642025
rect 494150 641951 494206 641960
rect 494164 639948 494192 641951
rect 499408 639948 499436 642359
rect 502064 641980 502116 641986
rect 502064 641922 502116 641928
rect 502076 639948 502104 641922
rect 504652 639948 504680 642767
rect 507306 642152 507362 642161
rect 507306 642087 507362 642096
rect 507320 639948 507348 642087
rect 509974 641880 510030 641889
rect 509974 641815 510030 641824
rect 517796 641844 517848 641850
rect 509988 639948 510016 641815
rect 517796 641786 517848 641792
rect 515862 641744 515918 641753
rect 515862 641679 515918 641688
rect 515220 640348 515272 640354
rect 515220 640290 515272 640296
rect 515232 639948 515260 640290
rect 515876 640257 515904 641679
rect 515862 640248 515918 640257
rect 515862 640183 515918 640192
rect 517808 639948 517836 641786
rect 520476 639948 520504 643039
rect 523132 643010 523184 643016
rect 523144 639948 523172 643010
rect 532332 642932 532384 642938
rect 532332 642874 532384 642880
rect 532240 642864 532292 642870
rect 532240 642806 532292 642812
rect 530400 642796 530452 642802
rect 530400 642738 530452 642744
rect 525706 641744 525762 641753
rect 525706 641679 525762 641688
rect 525720 639948 525748 641679
rect 530216 641640 530268 641646
rect 530216 641582 530268 641588
rect 529848 641572 529900 641578
rect 529848 641514 529900 641520
rect 529756 641436 529808 641442
rect 529756 641378 529808 641384
rect 529572 641096 529624 641102
rect 529572 641038 529624 641044
rect 529480 640960 529532 640966
rect 529480 640902 529532 640908
rect 462962 639704 463018 639713
rect 457128 639684 457378 639690
rect 457076 639678 457378 639684
rect 340970 639639 341026 639648
rect 446864 639668 446916 639674
rect 457088 639662 457378 639678
rect 462962 639639 463018 639648
rect 463238 639704 463294 639713
rect 463238 639639 463294 639648
rect 463422 639704 463478 639713
rect 463422 639639 463478 639648
rect 470138 639704 470194 639713
rect 471058 639704 471114 639713
rect 470194 639662 470534 639690
rect 470138 639639 470194 639648
rect 485134 639704 485190 639713
rect 480640 639674 481022 639690
rect 471058 639639 471114 639648
rect 480628 639668 481022 639674
rect 446864 639610 446916 639616
rect 480680 639662 481022 639668
rect 485134 639639 485190 639648
rect 496634 639704 496690 639713
rect 512274 639704 512330 639713
rect 496690 639662 496846 639690
rect 496634 639639 496690 639648
rect 528098 639704 528154 639713
rect 512330 639662 512578 639690
rect 512274 639639 512330 639648
rect 528154 639662 528402 639690
rect 528098 639639 528154 639648
rect 480628 639610 480680 639616
rect 231320 340190 231794 340218
rect 243556 340190 244122 340218
rect 261312 340190 261878 340218
rect 265544 340190 266110 340218
rect 266832 340190 267306 340218
rect 271064 340190 271630 340218
rect 272352 340190 272826 340218
rect 283300 340190 283866 340218
rect 288820 340190 289386 340218
rect 331692 340190 332258 340218
rect 334820 340190 335294 340218
rect 337212 340190 337778 340218
rect 342732 340190 343298 340218
rect 348252 340190 348818 340218
rect 356808 340190 357374 340218
rect 366008 340190 366574 340218
rect 373368 340190 373842 340218
rect 375760 340190 376326 340218
rect 382660 340190 383042 340218
rect 384408 340190 384882 340218
rect 408880 340190 409354 340218
rect 451752 340190 452226 340218
rect 457272 340190 457746 340218
rect 514050 340190 514616 340218
rect 229848 340054 230046 340082
rect 229848 335646 229876 340054
rect 229836 335640 229888 335646
rect 229836 335582 229888 335588
rect 230480 335640 230532 335646
rect 230480 335582 230532 335588
rect 229744 266348 229796 266354
rect 229744 266290 229796 266296
rect 230492 4962 230520 335582
rect 230480 4956 230532 4962
rect 230480 4898 230532 4904
rect 229100 4888 229152 4894
rect 229100 4830 229152 4836
rect 230112 4888 230164 4894
rect 230112 4830 230164 4836
rect 230124 480 230152 4830
rect 230584 4826 230612 340068
rect 230952 340054 231242 340082
rect 230952 335646 230980 340054
rect 230940 335640 230992 335646
rect 230940 335582 230992 335588
rect 231320 335458 231348 340190
rect 232424 337385 232452 340068
rect 232792 340054 233082 340082
rect 233252 340054 233634 340082
rect 233804 340054 234278 340082
rect 232410 337376 232466 337385
rect 232410 337311 232466 337320
rect 230676 335430 231348 335458
rect 230676 325582 230704 335430
rect 232792 331294 232820 340054
rect 231952 331288 232004 331294
rect 231952 331230 232004 331236
rect 232780 331288 232832 331294
rect 232780 331230 232832 331236
rect 230664 325576 230716 325582
rect 230664 325518 230716 325524
rect 231964 321638 231992 331230
rect 231952 321632 232004 321638
rect 231952 321574 232004 321580
rect 232044 321496 232096 321502
rect 232044 321438 232096 321444
rect 230848 318844 230900 318850
rect 230848 318786 230900 318792
rect 230860 311914 230888 318786
rect 232056 315994 232084 321438
rect 232044 315988 232096 315994
rect 232044 315930 232096 315936
rect 230664 311908 230716 311914
rect 230664 311850 230716 311856
rect 230848 311908 230900 311914
rect 230848 311850 230900 311856
rect 230676 304298 230704 311850
rect 230664 304292 230716 304298
rect 230664 304234 230716 304240
rect 230848 299532 230900 299538
rect 230848 299474 230900 299480
rect 230860 292602 230888 299474
rect 232044 298172 232096 298178
rect 232044 298114 232096 298120
rect 232056 298058 232084 298114
rect 232056 298030 232176 298058
rect 230664 292596 230716 292602
rect 230664 292538 230716 292544
rect 230848 292596 230900 292602
rect 230848 292538 230900 292544
rect 230676 283014 230704 292538
rect 232148 292482 232176 298030
rect 231964 292454 232176 292482
rect 231964 285938 231992 292454
rect 231952 285932 232004 285938
rect 231952 285874 232004 285880
rect 232320 285932 232372 285938
rect 232320 285874 232372 285880
rect 230664 283008 230716 283014
rect 230664 282950 230716 282956
rect 230664 282872 230716 282878
rect 230664 282814 230716 282820
rect 230676 280158 230704 282814
rect 230664 280152 230716 280158
rect 230664 280094 230716 280100
rect 230848 273284 230900 273290
rect 230848 273226 230900 273232
rect 230860 263634 230888 273226
rect 232332 270570 232360 285874
rect 232044 270564 232096 270570
rect 232044 270506 232096 270512
rect 232320 270564 232372 270570
rect 232320 270506 232372 270512
rect 232056 269090 232084 270506
rect 231964 269062 232084 269090
rect 231964 263634 231992 269062
rect 230848 263628 230900 263634
rect 230848 263570 230900 263576
rect 231952 263628 232004 263634
rect 231952 263570 232004 263576
rect 230940 263492 230992 263498
rect 230940 263434 230992 263440
rect 230952 254454 230980 263434
rect 231860 259480 231912 259486
rect 231860 259422 231912 259428
rect 231872 254658 231900 259422
rect 231860 254652 231912 254658
rect 231860 254594 231912 254600
rect 232044 254652 232096 254658
rect 232044 254594 232096 254600
rect 230940 254448 230992 254454
rect 230940 254390 230992 254396
rect 232056 244390 232084 254594
rect 232044 244384 232096 244390
rect 232044 244326 232096 244332
rect 231952 244248 232004 244254
rect 231952 244190 232004 244196
rect 230940 244180 230992 244186
rect 230940 244122 230992 244128
rect 230952 234734 230980 244122
rect 231964 240106 231992 244190
rect 231952 240100 232004 240106
rect 231952 240042 232004 240048
rect 232228 240100 232280 240106
rect 232228 240042 232280 240048
rect 230940 234728 230992 234734
rect 230940 234670 230992 234676
rect 230848 234592 230900 234598
rect 230848 234534 230900 234540
rect 230860 231849 230888 234534
rect 230662 231840 230718 231849
rect 230662 231775 230718 231784
rect 230846 231840 230902 231849
rect 230846 231775 230902 231784
rect 230676 222222 230704 231775
rect 232240 222290 232268 240042
rect 231952 222284 232004 222290
rect 231952 222226 232004 222232
rect 232228 222284 232280 222290
rect 232228 222226 232280 222232
rect 230664 222216 230716 222222
rect 230664 222158 230716 222164
rect 230940 222216 230992 222222
rect 230940 222158 230992 222164
rect 230952 215422 230980 222158
rect 231964 220833 231992 222226
rect 231766 220824 231822 220833
rect 231766 220759 231822 220768
rect 231950 220824 232006 220833
rect 231950 220759 232006 220768
rect 230940 215416 230992 215422
rect 230940 215358 230992 215364
rect 231780 215286 231808 220759
rect 230848 215280 230900 215286
rect 230848 215222 230900 215228
rect 231768 215280 231820 215286
rect 231768 215222 231820 215228
rect 231952 215280 232004 215286
rect 231952 215222 232004 215228
rect 230860 212537 230888 215222
rect 230662 212528 230718 212537
rect 230662 212463 230718 212472
rect 230846 212528 230902 212537
rect 230846 212463 230902 212472
rect 230676 202910 230704 212463
rect 231964 211154 231992 215222
rect 231964 211126 232084 211154
rect 232056 202910 232084 211126
rect 230664 202904 230716 202910
rect 230664 202846 230716 202852
rect 230940 202904 230992 202910
rect 230940 202846 230992 202852
rect 231952 202904 232004 202910
rect 231952 202846 232004 202852
rect 232044 202904 232096 202910
rect 232044 202846 232096 202852
rect 230952 196110 230980 202846
rect 230940 196104 230992 196110
rect 230940 196046 230992 196052
rect 230848 195968 230900 195974
rect 230848 195910 230900 195916
rect 230860 193225 230888 195910
rect 230662 193216 230718 193225
rect 230662 193151 230718 193160
rect 230846 193216 230902 193225
rect 230846 193151 230902 193160
rect 230676 183598 230704 193151
rect 231964 186266 231992 202846
rect 231964 186238 232084 186266
rect 230664 183592 230716 183598
rect 230664 183534 230716 183540
rect 230940 183592 230992 183598
rect 230940 183534 230992 183540
rect 230952 174418 230980 183534
rect 232056 182186 232084 186238
rect 232056 182158 232176 182186
rect 232148 180810 232176 182158
rect 232136 180804 232188 180810
rect 232136 180746 232188 180752
rect 230756 174412 230808 174418
rect 230756 174354 230808 174360
rect 230940 174412 230992 174418
rect 230940 174354 230992 174360
rect 230768 167006 230796 174354
rect 230756 167000 230808 167006
rect 230756 166942 230808 166948
rect 230940 167000 230992 167006
rect 230940 166942 230992 166948
rect 230952 164218 230980 166942
rect 230664 164212 230716 164218
rect 230664 164154 230716 164160
rect 230940 164212 230992 164218
rect 230940 164154 230992 164160
rect 230676 154601 230704 164154
rect 232136 162920 232188 162926
rect 232136 162862 232188 162868
rect 232148 161430 232176 162862
rect 232136 161424 232188 161430
rect 232136 161366 232188 161372
rect 230662 154592 230718 154601
rect 230662 154527 230718 154536
rect 230846 154592 230902 154601
rect 230846 154527 230848 154536
rect 230900 154527 230902 154536
rect 231032 154556 231084 154562
rect 230848 154498 230900 154504
rect 231032 154498 231084 154504
rect 231044 144945 231072 154498
rect 232228 151836 232280 151842
rect 232228 151778 232280 151784
rect 230754 144936 230810 144945
rect 230754 144871 230810 144880
rect 231030 144936 231086 144945
rect 231030 144871 231086 144880
rect 230768 138038 230796 144871
rect 232240 143585 232268 151778
rect 231950 143576 232006 143585
rect 232226 143576 232282 143585
rect 231950 143511 231952 143520
rect 232004 143511 232006 143520
rect 232044 143540 232096 143546
rect 231952 143482 232004 143488
rect 232226 143511 232282 143520
rect 232044 143482 232096 143488
rect 232056 142118 232084 143482
rect 232044 142112 232096 142118
rect 232044 142054 232096 142060
rect 230756 138032 230808 138038
rect 230756 137974 230808 137980
rect 230848 137964 230900 137970
rect 230848 137906 230900 137912
rect 230860 135250 230888 137906
rect 230848 135244 230900 135250
rect 230848 135186 230900 135192
rect 231032 135244 231084 135250
rect 231032 135186 231084 135192
rect 231044 125633 231072 135186
rect 230754 125624 230810 125633
rect 230754 125559 230810 125568
rect 231030 125624 231086 125633
rect 231030 125559 231086 125568
rect 230768 118726 230796 125559
rect 231952 124228 232004 124234
rect 231952 124170 232004 124176
rect 230756 118720 230808 118726
rect 230756 118662 230808 118668
rect 230848 118652 230900 118658
rect 230848 118594 230900 118600
rect 230860 115938 230888 118594
rect 230848 115932 230900 115938
rect 230848 115874 230900 115880
rect 231032 115932 231084 115938
rect 231032 115874 231084 115880
rect 231044 106321 231072 115874
rect 230754 106312 230810 106321
rect 230754 106247 230810 106256
rect 231030 106312 231086 106321
rect 231030 106247 231086 106256
rect 230768 99414 230796 106247
rect 231964 106214 231992 124170
rect 231952 106208 232004 106214
rect 231952 106150 232004 106156
rect 232136 106208 232188 106214
rect 232136 106150 232188 106156
rect 232148 104854 232176 106150
rect 232136 104848 232188 104854
rect 232136 104790 232188 104796
rect 230756 99408 230808 99414
rect 230756 99350 230808 99356
rect 230848 99340 230900 99346
rect 230848 99282 230900 99288
rect 230860 96626 230888 99282
rect 230848 96620 230900 96626
rect 230848 96562 230900 96568
rect 232228 95260 232280 95266
rect 232228 95202 232280 95208
rect 230848 89684 230900 89690
rect 230848 89626 230900 89632
rect 230860 86986 230888 89626
rect 232240 87009 232268 95202
rect 231950 87000 232006 87009
rect 230860 86958 230980 86986
rect 230952 80170 230980 86958
rect 231950 86935 232006 86944
rect 232226 87000 232282 87009
rect 232226 86935 232282 86944
rect 231964 85542 231992 86935
rect 231952 85536 232004 85542
rect 231952 85478 232004 85484
rect 230940 80164 230992 80170
rect 230940 80106 230992 80112
rect 230940 77308 230992 77314
rect 230940 77250 230992 77256
rect 230952 75886 230980 77250
rect 231952 75948 232004 75954
rect 231952 75890 232004 75896
rect 230940 75880 230992 75886
rect 230940 75822 230992 75828
rect 231964 72570 231992 75890
rect 231872 72542 231992 72570
rect 231872 67658 231900 72542
rect 231860 67652 231912 67658
rect 231860 67594 231912 67600
rect 231952 67652 232004 67658
rect 231952 67594 232004 67600
rect 231032 66292 231084 66298
rect 231032 66234 231084 66240
rect 231044 61418 231072 66234
rect 230768 61390 231072 61418
rect 230768 51082 230796 61390
rect 231964 58018 231992 67594
rect 231964 57990 232084 58018
rect 232056 56658 232084 57990
rect 231872 56630 232084 56658
rect 230768 51054 230888 51082
rect 230860 43518 230888 51054
rect 231872 46918 231900 56630
rect 231860 46912 231912 46918
rect 231860 46854 231912 46860
rect 232044 46912 232096 46918
rect 232044 46854 232096 46860
rect 230664 43512 230716 43518
rect 230664 43454 230716 43460
rect 230848 43512 230900 43518
rect 230848 43454 230900 43460
rect 230676 37262 230704 43454
rect 230664 37256 230716 37262
rect 230664 37198 230716 37204
rect 230756 37256 230808 37262
rect 230756 37198 230808 37204
rect 230768 27690 230796 37198
rect 232056 28966 232084 46854
rect 231860 28960 231912 28966
rect 231860 28902 231912 28908
rect 232044 28960 232096 28966
rect 232044 28902 232096 28908
rect 230768 27662 230888 27690
rect 230860 27606 230888 27662
rect 230756 27600 230808 27606
rect 230756 27542 230808 27548
rect 230848 27600 230900 27606
rect 230848 27542 230900 27548
rect 230768 26246 230796 27542
rect 230756 26240 230808 26246
rect 230756 26182 230808 26188
rect 231872 19310 231900 28902
rect 231860 19304 231912 19310
rect 231860 19246 231912 19252
rect 231952 19236 232004 19242
rect 231952 19178 232004 19184
rect 230664 8356 230716 8362
rect 230664 8298 230716 8304
rect 230676 7614 230704 8298
rect 230664 7608 230716 7614
rect 230664 7550 230716 7556
rect 231308 7608 231360 7614
rect 231308 7550 231360 7556
rect 230572 4820 230624 4826
rect 230572 4762 230624 4768
rect 231320 480 231348 7550
rect 231964 3369 231992 19178
rect 232504 8424 232556 8430
rect 232504 8366 232556 8372
rect 231950 3360 232006 3369
rect 231950 3295 232006 3304
rect 232516 480 232544 8366
rect 233252 5030 233280 340054
rect 233804 331242 233832 340054
rect 234908 337550 234936 340068
rect 234896 337544 234948 337550
rect 234896 337486 234948 337492
rect 235460 337414 235488 340068
rect 235448 337408 235500 337414
rect 235448 337350 235500 337356
rect 233344 331214 233832 331242
rect 233344 280158 233372 331214
rect 233332 280152 233384 280158
rect 233332 280094 233384 280100
rect 233516 280152 233568 280158
rect 233516 280094 233568 280100
rect 233528 244322 233556 280094
rect 233332 244316 233384 244322
rect 233332 244258 233384 244264
rect 233516 244316 233568 244322
rect 233516 244258 233568 244264
rect 233344 244202 233372 244258
rect 233344 244174 233464 244202
rect 233436 234682 233464 244174
rect 233436 234654 233556 234682
rect 233528 225010 233556 234654
rect 233332 225004 233384 225010
rect 233332 224946 233384 224952
rect 233516 225004 233568 225010
rect 233516 224946 233568 224952
rect 233344 215286 233372 224946
rect 233332 215280 233384 215286
rect 233332 215222 233384 215228
rect 233516 215280 233568 215286
rect 233516 215222 233568 215228
rect 233528 205222 233556 215222
rect 233516 205216 233568 205222
rect 233516 205158 233568 205164
rect 233516 205080 233568 205086
rect 233516 205022 233568 205028
rect 233528 186386 233556 205022
rect 233332 186380 233384 186386
rect 233332 186322 233384 186328
rect 233516 186380 233568 186386
rect 233516 186322 233568 186328
rect 233344 176610 233372 186322
rect 233344 176582 233464 176610
rect 233436 173890 233464 176582
rect 233436 173862 233556 173890
rect 233528 154442 233556 173862
rect 233436 154414 233556 154442
rect 233436 149682 233464 154414
rect 233344 149654 233464 149682
rect 233344 137986 233372 149654
rect 233344 137958 233556 137986
rect 233528 128382 233556 137958
rect 233332 128376 233384 128382
rect 233332 128318 233384 128324
rect 233516 128376 233568 128382
rect 233516 128318 233568 128324
rect 233344 118674 233372 128318
rect 233344 118646 233556 118674
rect 233528 109070 233556 118646
rect 233332 109064 233384 109070
rect 233332 109006 233384 109012
rect 233516 109064 233568 109070
rect 233516 109006 233568 109012
rect 233344 99362 233372 109006
rect 233344 99334 233556 99362
rect 233528 89758 233556 99334
rect 233332 89752 233384 89758
rect 233332 89694 233384 89700
rect 233516 89752 233568 89758
rect 233516 89694 233568 89700
rect 233344 80050 233372 89694
rect 233344 80022 233556 80050
rect 233528 51082 233556 80022
rect 233528 51054 233648 51082
rect 233620 50810 233648 51054
rect 233528 50782 233648 50810
rect 233528 41426 233556 50782
rect 233344 41398 233556 41426
rect 233344 31754 233372 41398
rect 233332 31748 233384 31754
rect 233332 31690 233384 31696
rect 233516 31748 233568 31754
rect 233516 31690 233568 31696
rect 233528 19394 233556 31690
rect 233436 19366 233556 19394
rect 233436 19310 233464 19366
rect 233332 19304 233384 19310
rect 233332 19246 233384 19252
rect 233424 19304 233476 19310
rect 233424 19246 233476 19252
rect 233344 7682 233372 19246
rect 236000 8356 236052 8362
rect 236000 8298 236052 8304
rect 233332 7676 233384 7682
rect 233332 7618 233384 7624
rect 234804 7676 234856 7682
rect 234804 7618 234856 7624
rect 233240 5024 233292 5030
rect 233240 4966 233292 4972
rect 233700 4820 233752 4826
rect 233700 4762 233752 4768
rect 233712 480 233740 4762
rect 234816 480 234844 7618
rect 236012 480 236040 8298
rect 236104 5098 236132 340068
rect 236196 340054 236762 340082
rect 236932 340054 237314 340082
rect 237576 340054 237958 340082
rect 238312 340054 238602 340082
rect 238864 340054 239154 340082
rect 236196 12510 236224 340054
rect 236932 327146 236960 340054
rect 237472 333668 237524 333674
rect 237472 333610 237524 333616
rect 236276 327140 236328 327146
rect 236276 327082 236328 327088
rect 236920 327140 236972 327146
rect 236920 327082 236972 327088
rect 236288 321450 236316 327082
rect 236288 321422 236408 321450
rect 236380 309126 236408 321422
rect 236276 309120 236328 309126
rect 236276 309062 236328 309068
rect 236368 309120 236420 309126
rect 236368 309062 236420 309068
rect 236288 298110 236316 309062
rect 236276 298104 236328 298110
rect 236276 298046 236328 298052
rect 236460 289740 236512 289746
rect 236460 289682 236512 289688
rect 236472 288425 236500 289682
rect 236458 288416 236514 288425
rect 236458 288351 236514 288360
rect 236642 288416 236698 288425
rect 236642 288351 236698 288360
rect 236380 278798 236408 278829
rect 236656 278798 236684 288351
rect 236368 278792 236420 278798
rect 236288 278740 236368 278746
rect 236288 278734 236420 278740
rect 236644 278792 236696 278798
rect 236644 278734 236696 278740
rect 236288 278718 236408 278734
rect 236288 277386 236316 278718
rect 236288 277358 236408 277386
rect 236380 270570 236408 277358
rect 236368 270564 236420 270570
rect 236368 270506 236420 270512
rect 236276 270496 236328 270502
rect 236276 270438 236328 270444
rect 236288 263634 236316 270438
rect 236276 263628 236328 263634
rect 236276 263570 236328 263576
rect 236368 263560 236420 263566
rect 236368 263502 236420 263508
rect 236380 253910 236408 263502
rect 236368 253904 236420 253910
rect 236368 253846 236420 253852
rect 236276 253768 236328 253774
rect 236276 253710 236328 253716
rect 236288 244322 236316 253710
rect 236276 244316 236328 244322
rect 236276 244258 236328 244264
rect 236276 240236 236328 240242
rect 236276 240178 236328 240184
rect 236288 240106 236316 240178
rect 236276 240100 236328 240106
rect 236276 240042 236328 240048
rect 236276 230580 236328 230586
rect 236276 230522 236328 230528
rect 236288 230489 236316 230522
rect 236274 230480 236330 230489
rect 236274 230415 236330 230424
rect 236458 230480 236514 230489
rect 236458 230415 236514 230424
rect 236288 220862 236316 220893
rect 236472 220862 236500 230415
rect 236276 220856 236328 220862
rect 236460 220856 236512 220862
rect 236328 220804 236408 220810
rect 236276 220798 236408 220804
rect 236460 220798 236512 220804
rect 236288 220782 236408 220798
rect 236380 216034 236408 220782
rect 236368 216028 236420 216034
rect 236368 215970 236420 215976
rect 236552 216028 236604 216034
rect 236552 215970 236604 215976
rect 236564 211177 236592 215970
rect 236274 211168 236330 211177
rect 236274 211103 236330 211112
rect 236550 211168 236606 211177
rect 236550 211103 236606 211112
rect 236288 205630 236316 211103
rect 236276 205624 236328 205630
rect 236276 205566 236328 205572
rect 236276 202904 236328 202910
rect 236276 202846 236328 202852
rect 236288 198694 236316 202846
rect 236276 198688 236328 198694
rect 236276 198630 236328 198636
rect 236368 189100 236420 189106
rect 236368 189042 236420 189048
rect 236380 179382 236408 189042
rect 236368 179376 236420 179382
rect 236368 179318 236420 179324
rect 236368 161492 236420 161498
rect 236368 161434 236420 161440
rect 236380 153202 236408 161434
rect 236276 153196 236328 153202
rect 236276 153138 236328 153144
rect 236368 153196 236420 153202
rect 236368 153138 236420 153144
rect 236288 143546 236316 153138
rect 236276 143540 236328 143546
rect 236276 143482 236328 143488
rect 236460 143540 236512 143546
rect 236460 143482 236512 143488
rect 236472 142118 236500 143482
rect 236460 142112 236512 142118
rect 236460 142054 236512 142060
rect 236460 132524 236512 132530
rect 236460 132466 236512 132472
rect 236472 124302 236500 132466
rect 236368 124296 236420 124302
rect 236368 124238 236420 124244
rect 236460 124296 236512 124302
rect 236460 124238 236512 124244
rect 236380 122806 236408 124238
rect 236368 122800 236420 122806
rect 236368 122742 236420 122748
rect 236460 113212 236512 113218
rect 236460 113154 236512 113160
rect 236472 106321 236500 113154
rect 236274 106312 236330 106321
rect 236274 106247 236330 106256
rect 236458 106312 236514 106321
rect 236458 106247 236514 106256
rect 236288 106214 236316 106247
rect 236276 106208 236328 106214
rect 236276 106150 236328 106156
rect 236552 106208 236604 106214
rect 236552 106150 236604 106156
rect 236564 96665 236592 106150
rect 236366 96656 236422 96665
rect 236366 96591 236422 96600
rect 236550 96656 236606 96665
rect 236550 96591 236606 96600
rect 236380 87145 236408 96591
rect 236366 87136 236422 87145
rect 236366 87071 236422 87080
rect 236274 87000 236330 87009
rect 236274 86935 236330 86944
rect 236288 85542 236316 86935
rect 236276 85536 236328 85542
rect 236276 85478 236328 85484
rect 236276 75948 236328 75954
rect 236276 75890 236328 75896
rect 236288 70378 236316 75890
rect 236276 70372 236328 70378
rect 236276 70314 236328 70320
rect 236276 67652 236328 67658
rect 236276 67594 236328 67600
rect 236288 66230 236316 67594
rect 236276 66224 236328 66230
rect 236276 66166 236328 66172
rect 236276 47048 236328 47054
rect 236276 46990 236328 46996
rect 236288 46918 236316 46990
rect 236276 46912 236328 46918
rect 236276 46854 236328 46860
rect 236460 46912 236512 46918
rect 236460 46854 236512 46860
rect 236472 41290 236500 46854
rect 236380 41262 236500 41290
rect 236380 29034 236408 41262
rect 236276 29028 236328 29034
rect 236276 28970 236328 28976
rect 236368 29028 236420 29034
rect 236368 28970 236420 28976
rect 236288 19378 236316 28970
rect 236276 19372 236328 19378
rect 236276 19314 236328 19320
rect 236368 19236 236420 19242
rect 236368 19178 236420 19184
rect 236184 12504 236236 12510
rect 236184 12446 236236 12452
rect 236092 5092 236144 5098
rect 236092 5034 236144 5040
rect 236380 3534 236408 19178
rect 237484 5166 237512 333610
rect 237472 5160 237524 5166
rect 237472 5102 237524 5108
rect 237196 4956 237248 4962
rect 237196 4898 237248 4904
rect 236368 3528 236420 3534
rect 236368 3470 236420 3476
rect 237208 480 237236 4898
rect 237576 3466 237604 340054
rect 238312 333674 238340 340054
rect 238300 333668 238352 333674
rect 238300 333610 238352 333616
rect 238758 170368 238814 170377
rect 238758 170303 238760 170312
rect 238812 170303 238814 170312
rect 238760 170274 238812 170280
rect 238864 13122 238892 340054
rect 239784 337414 239812 340068
rect 240428 337754 240456 340068
rect 240612 340054 240994 340082
rect 241638 340054 241744 340082
rect 240416 337748 240468 337754
rect 240416 337690 240468 337696
rect 239772 337408 239824 337414
rect 239772 337350 239824 337356
rect 240612 331242 240640 340054
rect 241520 335640 241572 335646
rect 241520 335582 241572 335588
rect 240152 331214 240640 331242
rect 240152 331106 240180 331214
rect 240152 331078 240272 331106
rect 240244 302274 240272 331078
rect 240152 302246 240272 302274
rect 240152 302138 240180 302246
rect 240152 302110 240272 302138
rect 240244 282962 240272 302110
rect 240152 282934 240272 282962
rect 240152 282826 240180 282934
rect 240152 282798 240272 282826
rect 240244 263650 240272 282798
rect 240152 263622 240272 263650
rect 240152 263514 240180 263622
rect 240152 263486 240272 263514
rect 240244 244338 240272 263486
rect 240152 244310 240272 244338
rect 240152 244202 240180 244310
rect 240152 244174 240272 244202
rect 240244 225026 240272 244174
rect 240152 224998 240272 225026
rect 240152 224890 240180 224998
rect 240152 224862 240272 224890
rect 240244 205714 240272 224862
rect 240152 205686 240272 205714
rect 240152 205578 240180 205686
rect 240152 205550 240272 205578
rect 240244 186402 240272 205550
rect 240152 186374 240272 186402
rect 240152 186266 240180 186374
rect 240152 186238 240272 186266
rect 240244 167090 240272 186238
rect 240244 167062 240364 167090
rect 240336 164257 240364 167062
rect 240138 164248 240194 164257
rect 240138 164183 240140 164192
rect 240192 164183 240194 164192
rect 240322 164248 240378 164257
rect 240322 164183 240324 164192
rect 240140 164154 240192 164160
rect 240376 164183 240378 164192
rect 240324 164154 240376 164160
rect 240336 159202 240364 164154
rect 240244 159174 240364 159202
rect 240244 153202 240272 159174
rect 240140 153196 240192 153202
rect 240140 153138 240192 153144
rect 240232 153196 240284 153202
rect 240232 153138 240284 153144
rect 240152 143721 240180 153138
rect 240138 143712 240194 143721
rect 240138 143647 240194 143656
rect 240138 143576 240194 143585
rect 240138 143511 240194 143520
rect 240152 142118 240180 143511
rect 240140 142112 240192 142118
rect 240140 142054 240192 142060
rect 240324 132524 240376 132530
rect 240324 132466 240376 132472
rect 240336 128194 240364 132466
rect 240152 128166 240364 128194
rect 240152 119354 240180 128166
rect 240152 119326 240272 119354
rect 240244 89842 240272 119326
rect 240152 89814 240272 89842
rect 240152 89706 240180 89814
rect 240152 89678 240272 89706
rect 240244 70514 240272 89678
rect 240232 70508 240284 70514
rect 240232 70450 240284 70456
rect 240232 70372 240284 70378
rect 240232 70314 240284 70320
rect 240048 14068 240100 14074
rect 240048 14010 240100 14016
rect 238852 13116 238904 13122
rect 238852 13058 238904 13064
rect 238392 7064 238444 7070
rect 238392 7006 238444 7012
rect 237564 3460 237616 3466
rect 237564 3402 237616 3408
rect 238404 480 238432 7006
rect 240060 3670 240088 14010
rect 240244 5234 240272 70314
rect 240232 5228 240284 5234
rect 240232 5170 240284 5176
rect 240784 5024 240836 5030
rect 240784 4966 240836 4972
rect 239588 3664 239640 3670
rect 239588 3606 239640 3612
rect 240048 3664 240100 3670
rect 240048 3606 240100 3612
rect 239600 480 239628 3606
rect 240796 480 240824 4966
rect 241532 3602 241560 335582
rect 241716 14482 241744 340054
rect 241992 340054 242282 340082
rect 242452 340054 242834 340082
rect 242912 340054 243478 340082
rect 241992 335646 242020 340054
rect 241980 335640 242032 335646
rect 241980 335582 242032 335588
rect 242452 328506 242480 340054
rect 241796 328500 241848 328506
rect 241796 328442 241848 328448
rect 242440 328500 242492 328506
rect 242440 328442 242492 328448
rect 241808 299470 241836 328442
rect 241796 299464 241848 299470
rect 241796 299406 241848 299412
rect 241796 289876 241848 289882
rect 241796 289818 241848 289824
rect 241808 280158 241836 289818
rect 241796 280152 241848 280158
rect 241796 280094 241848 280100
rect 242808 280152 242860 280158
rect 242808 280094 242860 280100
rect 242820 270609 242848 280094
rect 242806 270600 242862 270609
rect 241796 270564 241848 270570
rect 242806 270535 242862 270544
rect 241796 270506 241848 270512
rect 241808 260846 241836 270506
rect 241796 260840 241848 260846
rect 241796 260782 241848 260788
rect 242808 260840 242860 260846
rect 242808 260782 242860 260788
rect 242820 251297 242848 260782
rect 242806 251288 242862 251297
rect 241796 251252 241848 251258
rect 242806 251223 242862 251232
rect 241796 251194 241848 251200
rect 241808 183569 241836 251194
rect 241794 183560 241850 183569
rect 241794 183495 241850 183504
rect 241978 183560 242034 183569
rect 241978 183495 242034 183504
rect 241992 173942 242020 183495
rect 241796 173936 241848 173942
rect 241796 173878 241848 173884
rect 241980 173936 242032 173942
rect 241980 173878 242032 173884
rect 241808 125594 241836 173878
rect 241796 125588 241848 125594
rect 241796 125530 241848 125536
rect 241980 125588 242032 125594
rect 241980 125530 242032 125536
rect 241992 115977 242020 125530
rect 241794 115968 241850 115977
rect 241794 115903 241850 115912
rect 241978 115968 242034 115977
rect 241978 115903 242034 115912
rect 241808 106282 241836 115903
rect 241796 106276 241848 106282
rect 241796 106218 241848 106224
rect 241980 106276 242032 106282
rect 241980 106218 242032 106224
rect 241992 96665 242020 106218
rect 241794 96656 241850 96665
rect 241794 96591 241850 96600
rect 241978 96656 242034 96665
rect 241978 96591 242034 96600
rect 241808 86970 241836 96591
rect 241796 86964 241848 86970
rect 241796 86906 241848 86912
rect 241796 77308 241848 77314
rect 241796 77250 241848 77256
rect 241704 14476 241756 14482
rect 241704 14418 241756 14424
rect 241520 3596 241572 3602
rect 241520 3538 241572 3544
rect 241808 3534 241836 77250
rect 242912 7750 242940 340054
rect 243556 327321 243584 340190
rect 244660 337550 244688 340068
rect 244844 340054 245318 340082
rect 245764 340054 245962 340082
rect 244648 337544 244700 337550
rect 244648 337486 244700 337492
rect 244844 331242 244872 340054
rect 245660 335572 245712 335578
rect 245660 335514 245712 335520
rect 244476 331214 244872 331242
rect 243542 327312 243598 327321
rect 243542 327247 243598 327256
rect 243082 327176 243138 327185
rect 243082 327111 243138 327120
rect 243096 307766 243124 327111
rect 244476 311930 244504 331214
rect 244384 311902 244504 311930
rect 244384 311794 244412 311902
rect 244384 311766 244504 311794
rect 243084 307760 243136 307766
rect 243084 307702 243136 307708
rect 242992 298172 243044 298178
rect 242992 298114 243044 298120
rect 243004 282878 243032 298114
rect 242992 282872 243044 282878
rect 242992 282814 243044 282820
rect 243176 282872 243228 282878
rect 243176 282814 243228 282820
rect 243188 280158 243216 282814
rect 244476 280158 244504 311766
rect 243176 280152 243228 280158
rect 243176 280094 243228 280100
rect 244464 280152 244516 280158
rect 244464 280094 244516 280100
rect 244556 280152 244608 280158
rect 244556 280094 244608 280100
rect 244568 273170 244596 280094
rect 244476 273142 244596 273170
rect 243174 270464 243230 270473
rect 243174 270399 243230 270408
rect 243188 263634 243216 270399
rect 243176 263628 243228 263634
rect 243176 263570 243228 263576
rect 243176 263492 243228 263498
rect 243176 263434 243228 263440
rect 243188 260846 243216 263434
rect 244476 260846 244504 273142
rect 243176 260840 243228 260846
rect 243176 260782 243228 260788
rect 244464 260840 244516 260846
rect 244464 260782 244516 260788
rect 244556 260772 244608 260778
rect 244556 260714 244608 260720
rect 244568 253858 244596 260714
rect 244476 253830 244596 253858
rect 242990 251152 243046 251161
rect 242990 251087 243046 251096
rect 243004 241534 243032 251087
rect 242992 241528 243044 241534
rect 242990 241496 242992 241505
rect 243176 241528 243228 241534
rect 243044 241496 243046 241505
rect 242990 241431 243046 241440
rect 243174 241496 243176 241505
rect 243228 241496 243230 241505
rect 243174 241431 243230 241440
rect 243004 231878 243032 241431
rect 242992 231872 243044 231878
rect 242992 231814 243044 231820
rect 243084 231872 243136 231878
rect 243136 231820 243216 231826
rect 243084 231814 243216 231820
rect 243096 231798 243216 231814
rect 243188 231742 243216 231798
rect 243176 231736 243228 231742
rect 243176 231678 243228 231684
rect 243360 224256 243412 224262
rect 243360 224198 243412 224204
rect 243372 219434 243400 224198
rect 243084 219428 243136 219434
rect 243084 219370 243136 219376
rect 243360 219428 243412 219434
rect 243360 219370 243412 219376
rect 243096 218006 243124 219370
rect 243084 218000 243136 218006
rect 243084 217942 243136 217948
rect 243084 201476 243136 201482
rect 243084 201418 243136 201424
rect 243096 200138 243124 201418
rect 243096 200110 243216 200138
rect 243188 196110 243216 200110
rect 243176 196104 243228 196110
rect 244476 196058 244504 253830
rect 243176 196046 243228 196052
rect 244384 196030 244504 196058
rect 243176 195968 243228 195974
rect 243176 195910 243228 195916
rect 244384 195922 244412 196030
rect 243188 180810 243216 195910
rect 244384 195894 244504 195922
rect 244476 186998 244504 195894
rect 244464 186992 244516 186998
rect 244464 186934 244516 186940
rect 244648 186992 244700 186998
rect 244648 186934 244700 186940
rect 244660 182209 244688 186934
rect 244462 182200 244518 182209
rect 244462 182135 244518 182144
rect 244646 182200 244702 182209
rect 244646 182135 244702 182144
rect 243176 180804 243228 180810
rect 243176 180746 243228 180752
rect 243360 180804 243412 180810
rect 243360 180746 243412 180752
rect 243372 171193 243400 180746
rect 243174 171184 243230 171193
rect 243096 171142 243174 171170
rect 243096 171086 243124 171142
rect 243174 171119 243230 171128
rect 243358 171184 243414 171193
rect 243358 171119 243414 171128
rect 243084 171080 243136 171086
rect 243084 171022 243136 171028
rect 243176 161492 243228 161498
rect 243176 161434 243228 161440
rect 243188 157486 243216 161434
rect 243176 157480 243228 157486
rect 244476 157434 244504 182135
rect 243176 157422 243228 157428
rect 244384 157406 244504 157434
rect 243176 157344 243228 157350
rect 243176 157286 243228 157292
rect 244384 157298 244412 157406
rect 243188 135266 243216 157286
rect 244384 157270 244504 157298
rect 244476 138038 244504 157270
rect 244464 138032 244516 138038
rect 244464 137974 244516 137980
rect 244464 137896 244516 137902
rect 244464 137838 244516 137844
rect 243096 135238 243216 135266
rect 243096 133890 243124 135238
rect 243084 133884 243136 133890
rect 243084 133826 243136 133832
rect 243268 124228 243320 124234
rect 243268 124170 243320 124176
rect 243280 119218 243308 124170
rect 243096 119190 243308 119218
rect 243096 109070 243124 119190
rect 243084 109064 243136 109070
rect 243084 109006 243136 109012
rect 243176 108996 243228 109002
rect 243176 108938 243228 108944
rect 243188 106214 243216 108938
rect 243176 106208 243228 106214
rect 243176 106150 243228 106156
rect 243176 96756 243228 96762
rect 243176 96698 243228 96704
rect 243188 96626 243216 96698
rect 243084 96620 243136 96626
rect 243084 96562 243136 96568
rect 243176 96620 243228 96626
rect 243176 96562 243228 96568
rect 243096 86902 243124 96562
rect 243084 86896 243136 86902
rect 243084 86838 243136 86844
rect 243268 86896 243320 86902
rect 243268 86838 243320 86844
rect 243280 77489 243308 86838
rect 244476 80102 244504 137838
rect 244464 80096 244516 80102
rect 244464 80038 244516 80044
rect 244464 79960 244516 79966
rect 244464 79902 244516 79908
rect 243266 77480 243322 77489
rect 243266 77415 243322 77424
rect 243082 75984 243138 75993
rect 243082 75919 243138 75928
rect 243096 70446 243124 75919
rect 243084 70440 243136 70446
rect 243084 70382 243136 70388
rect 243176 70304 243228 70310
rect 243176 70246 243228 70252
rect 243188 64870 243216 70246
rect 243176 64864 243228 64870
rect 243176 64806 243228 64812
rect 244476 60738 244504 79902
rect 244384 60710 244504 60738
rect 244384 60602 244412 60710
rect 244384 60574 244504 60602
rect 244476 56574 244504 60574
rect 244464 56568 244516 56574
rect 244464 56510 244516 56516
rect 242992 55276 243044 55282
rect 242992 55218 243044 55224
rect 243004 50946 243032 55218
rect 243004 50918 243216 50946
rect 243188 46918 243216 50918
rect 244372 46980 244424 46986
rect 244372 46922 244424 46928
rect 243176 46912 243228 46918
rect 243176 46854 243228 46860
rect 243268 46912 243320 46918
rect 243268 46854 243320 46860
rect 243280 45558 243308 46854
rect 243268 45552 243320 45558
rect 243268 45494 243320 45500
rect 244384 42106 244412 46922
rect 244384 42078 244504 42106
rect 242992 35964 243044 35970
rect 242992 35906 243044 35912
rect 243004 31634 243032 35906
rect 243004 31606 243124 31634
rect 243096 15978 243124 31606
rect 244476 28966 244504 42078
rect 244464 28960 244516 28966
rect 244464 28902 244516 28908
rect 244556 28960 244608 28966
rect 244556 28902 244608 28908
rect 244186 16824 244242 16833
rect 244370 16824 244426 16833
rect 244242 16782 244370 16810
rect 244186 16759 244242 16768
rect 244370 16759 244426 16768
rect 243084 15972 243136 15978
rect 243084 15914 243136 15920
rect 244188 14476 244240 14482
rect 244188 14418 244240 14424
rect 242900 7744 242952 7750
rect 242900 7686 242952 7692
rect 241980 6996 242032 7002
rect 241980 6938 242032 6944
rect 241796 3528 241848 3534
rect 241796 3470 241848 3476
rect 241992 480 242020 6938
rect 244200 3670 244228 14418
rect 244568 9722 244596 28902
rect 244280 9716 244332 9722
rect 244280 9658 244332 9664
rect 244556 9716 244608 9722
rect 244556 9658 244608 9664
rect 244292 7818 244320 9658
rect 244280 7812 244332 7818
rect 244280 7754 244332 7760
rect 245568 7744 245620 7750
rect 245568 7686 245620 7692
rect 244372 5092 244424 5098
rect 244372 5034 244424 5040
rect 243176 3664 243228 3670
rect 243176 3606 243228 3612
rect 244188 3664 244240 3670
rect 244188 3606 244240 3612
rect 243188 480 243216 3606
rect 244384 480 244412 5034
rect 245580 480 245608 7686
rect 245672 3738 245700 335514
rect 245764 15910 245792 340054
rect 246304 337544 246356 337550
rect 246304 337486 246356 337492
rect 245752 15904 245804 15910
rect 245752 15846 245804 15852
rect 246316 14142 246344 337486
rect 246500 335578 246528 340068
rect 247158 340054 247264 340082
rect 246488 335572 246540 335578
rect 246488 335514 246540 335520
rect 246304 14136 246356 14142
rect 246304 14078 246356 14084
rect 246764 9920 246816 9926
rect 246764 9862 246816 9868
rect 245660 3732 245712 3738
rect 245660 3674 245712 3680
rect 246776 480 246804 9862
rect 247236 7886 247264 340054
rect 247696 337822 247724 340068
rect 247684 337816 247736 337822
rect 247684 337758 247736 337764
rect 248340 337618 248368 340068
rect 248524 340054 248998 340082
rect 248420 337748 248472 337754
rect 248420 337690 248472 337696
rect 248328 337612 248380 337618
rect 248328 337554 248380 337560
rect 248328 170332 248380 170338
rect 248328 170274 248380 170280
rect 248340 170105 248368 170274
rect 248326 170096 248382 170105
rect 248326 170031 248382 170040
rect 247224 7880 247276 7886
rect 247224 7822 247276 7828
rect 247960 5160 248012 5166
rect 247960 5102 248012 5108
rect 247972 480 248000 5102
rect 248432 3806 248460 337690
rect 248524 7954 248552 340054
rect 249536 337754 249564 340068
rect 249812 340054 250194 340082
rect 249524 337748 249576 337754
rect 249524 337690 249576 337696
rect 249246 307728 249302 307737
rect 249246 307663 249302 307672
rect 249260 298353 249288 307663
rect 249246 298344 249302 298353
rect 249246 298279 249302 298288
rect 249246 279848 249302 279857
rect 249246 279783 249302 279792
rect 249260 270609 249288 279783
rect 249246 270600 249302 270609
rect 249246 270535 249302 270544
rect 249246 270464 249302 270473
rect 249246 270399 249302 270408
rect 249260 260953 249288 270399
rect 249246 260944 249302 260953
rect 249246 260879 249302 260888
rect 249246 251152 249302 251161
rect 249246 251087 249302 251096
rect 249260 241777 249288 251087
rect 249246 241768 249302 241777
rect 249246 241703 249302 241712
rect 249430 222184 249486 222193
rect 249430 222119 249486 222128
rect 249444 214577 249472 222119
rect 249430 214568 249486 214577
rect 249430 214503 249486 214512
rect 249522 199880 249578 199889
rect 249522 199815 249578 199824
rect 249536 185609 249564 199815
rect 249522 185600 249578 185609
rect 249522 185535 249578 185544
rect 249614 179344 249670 179353
rect 249614 179279 249670 179288
rect 249628 169969 249656 179279
rect 249614 169960 249670 169969
rect 249614 169895 249670 169904
rect 248512 7948 248564 7954
rect 248512 7890 248564 7896
rect 249156 7812 249208 7818
rect 249156 7754 249208 7760
rect 248420 3800 248472 3806
rect 248420 3742 248472 3748
rect 249168 480 249196 7754
rect 249812 3874 249840 340054
rect 250824 337754 250852 340068
rect 251376 337890 251404 340068
rect 251364 337884 251416 337890
rect 251364 337826 251416 337832
rect 249984 337748 250036 337754
rect 249984 337690 250036 337696
rect 250812 337748 250864 337754
rect 250812 337690 250864 337696
rect 249996 321706 250024 337690
rect 252020 337346 252048 340068
rect 252008 337340 252060 337346
rect 252008 337282 252060 337288
rect 252560 336320 252612 336326
rect 252560 336262 252612 336268
rect 251824 334416 251876 334422
rect 251824 334358 251876 334364
rect 249984 321700 250036 321706
rect 249984 321642 250036 321648
rect 249984 317484 250036 317490
rect 249984 317426 250036 317432
rect 249996 311914 250024 317426
rect 249984 311908 250036 311914
rect 249984 311850 250036 311856
rect 249892 311840 249944 311846
rect 249892 311782 249944 311788
rect 249904 302410 249932 311782
rect 249904 302382 250116 302410
rect 250088 299418 250116 302382
rect 249904 299390 250116 299418
rect 249904 298110 249932 299390
rect 249892 298104 249944 298110
rect 249892 298046 249944 298052
rect 249892 288448 249944 288454
rect 249892 288390 249944 288396
rect 249904 285870 249932 288390
rect 249892 285864 249944 285870
rect 249892 285806 249944 285812
rect 250076 278792 250128 278798
rect 250076 278734 250128 278740
rect 250088 273170 250116 278734
rect 249996 273142 250116 273170
rect 249996 260846 250024 273142
rect 249984 260840 250036 260846
rect 249984 260782 250036 260788
rect 250076 260772 250128 260778
rect 250076 260714 250128 260720
rect 250088 253858 250116 260714
rect 249996 253830 250116 253858
rect 249996 196058 250024 253830
rect 249904 196030 250024 196058
rect 249904 195922 249932 196030
rect 249904 195894 250024 195922
rect 249996 186946 250024 195894
rect 249996 186918 250116 186946
rect 250088 174010 250116 186918
rect 250076 174004 250128 174010
rect 250076 173946 250128 173952
rect 249984 173868 250036 173874
rect 249984 173810 250036 173816
rect 249996 157434 250024 173810
rect 249904 157406 250024 157434
rect 249904 157298 249932 157406
rect 249904 157270 250024 157298
rect 249996 138038 250024 157270
rect 249984 138032 250036 138038
rect 249984 137974 250036 137980
rect 249984 137896 250036 137902
rect 249984 137838 250036 137844
rect 249996 60738 250024 137838
rect 249904 60710 250024 60738
rect 249904 60602 249932 60710
rect 249904 60574 250024 60602
rect 249996 56574 250024 60574
rect 249984 56568 250036 56574
rect 249984 56510 250036 56516
rect 249984 46980 250036 46986
rect 249984 46922 250036 46928
rect 249996 28914 250024 46922
rect 249996 28886 250116 28914
rect 250088 9722 250116 28886
rect 250352 9852 250404 9858
rect 250352 9794 250404 9800
rect 249984 9716 250036 9722
rect 249984 9658 250036 9664
rect 250076 9716 250128 9722
rect 250076 9658 250128 9664
rect 249996 8022 250024 9658
rect 249984 8016 250036 8022
rect 249984 7958 250036 7964
rect 249800 3868 249852 3874
rect 249800 3810 249852 3816
rect 250364 480 250392 9794
rect 251456 5228 251508 5234
rect 251456 5170 251508 5176
rect 251468 480 251496 5170
rect 251836 3942 251864 334358
rect 252572 309194 252600 336262
rect 252664 328438 252692 340068
rect 253216 334422 253244 340068
rect 253860 336326 253888 340068
rect 253952 340054 254518 340082
rect 253848 336320 253900 336326
rect 253848 336262 253900 336268
rect 253204 334416 253256 334422
rect 253204 334358 253256 334364
rect 253204 334280 253256 334286
rect 253204 334222 253256 334228
rect 252652 328432 252704 328438
rect 252652 328374 252704 328380
rect 252652 320136 252704 320142
rect 252652 320078 252704 320084
rect 252560 309188 252612 309194
rect 252560 309130 252612 309136
rect 252466 212528 252522 212537
rect 252466 212463 252522 212472
rect 252480 202910 252508 212463
rect 252468 202904 252520 202910
rect 252468 202846 252520 202852
rect 252560 202904 252612 202910
rect 252560 202846 252612 202852
rect 252572 193254 252600 202846
rect 252560 193248 252612 193254
rect 252560 193190 252612 193196
rect 252560 164212 252612 164218
rect 252560 164154 252612 164160
rect 252572 154601 252600 164154
rect 252558 154592 252614 154601
rect 252558 154527 252614 154536
rect 252560 145580 252612 145586
rect 252560 145522 252612 145528
rect 252572 135289 252600 145522
rect 252558 135280 252614 135289
rect 252558 135215 252614 135224
rect 252664 8090 252692 320078
rect 252744 309188 252796 309194
rect 252744 309130 252796 309136
rect 252756 270502 252784 309130
rect 252744 270496 252796 270502
rect 252744 270438 252796 270444
rect 252744 260908 252796 260914
rect 252744 260850 252796 260856
rect 252756 251190 252784 260850
rect 252744 251184 252796 251190
rect 252744 251126 252796 251132
rect 252756 241534 252784 241565
rect 252744 241528 252796 241534
rect 252796 241476 252876 241482
rect 252744 241470 252876 241476
rect 252756 241454 252876 241470
rect 252848 231962 252876 241454
rect 252756 231934 252876 231962
rect 252756 231849 252784 231934
rect 252742 231840 252798 231849
rect 252742 231775 252798 231784
rect 252926 231840 252982 231849
rect 252926 231775 252982 231784
rect 252756 222222 252784 222253
rect 252940 222222 252968 231775
rect 252744 222216 252796 222222
rect 252928 222216 252980 222222
rect 252796 222164 252876 222170
rect 252744 222158 252876 222164
rect 252928 222158 252980 222164
rect 252756 222142 252876 222158
rect 252848 212566 252876 222142
rect 252744 212560 252796 212566
rect 252742 212528 252744 212537
rect 252836 212560 252888 212566
rect 252796 212528 252798 212537
rect 252836 212502 252888 212508
rect 252742 212463 252798 212472
rect 252744 193248 252796 193254
rect 252744 193190 252796 193196
rect 252756 183598 252784 193190
rect 252744 183592 252796 183598
rect 252744 183534 252796 183540
rect 252836 183456 252888 183462
rect 252836 183398 252888 183404
rect 252848 182170 252876 183398
rect 252836 182164 252888 182170
rect 252836 182106 252888 182112
rect 252836 172576 252888 172582
rect 252836 172518 252888 172524
rect 252848 164218 252876 172518
rect 252836 164212 252888 164218
rect 252836 164154 252888 164160
rect 252742 154592 252798 154601
rect 252742 154527 252798 154536
rect 252756 145586 252784 154527
rect 252744 145580 252796 145586
rect 252744 145522 252796 145528
rect 252742 135280 252798 135289
rect 252742 135215 252798 135224
rect 252756 125594 252784 135215
rect 252744 125588 252796 125594
rect 252744 125530 252796 125536
rect 252928 125588 252980 125594
rect 252928 125530 252980 125536
rect 252940 115977 252968 125530
rect 252742 115968 252798 115977
rect 252742 115903 252798 115912
rect 252926 115968 252982 115977
rect 252926 115903 252982 115912
rect 252756 106214 252784 115903
rect 252744 106208 252796 106214
rect 252744 106150 252796 106156
rect 252744 96688 252796 96694
rect 252744 96630 252796 96636
rect 252756 86902 252784 96630
rect 252744 86896 252796 86902
rect 252744 86838 252796 86844
rect 252744 77308 252796 77314
rect 252744 77250 252796 77256
rect 252756 37398 252784 77250
rect 252744 37392 252796 37398
rect 252744 37334 252796 37340
rect 252836 29028 252888 29034
rect 252836 28970 252888 28976
rect 252848 27606 252876 28970
rect 252836 27600 252888 27606
rect 252836 27542 252888 27548
rect 252836 18012 252888 18018
rect 252836 17954 252888 17960
rect 252848 12458 252876 17954
rect 252756 12430 252876 12458
rect 252652 8084 252704 8090
rect 252652 8026 252704 8032
rect 252652 7880 252704 7886
rect 252652 7822 252704 7828
rect 251824 3936 251876 3942
rect 251824 3878 251876 3884
rect 252664 480 252692 7822
rect 252756 4010 252784 12430
rect 253216 4078 253244 334222
rect 253848 9784 253900 9790
rect 253848 9726 253900 9732
rect 253204 4072 253256 4078
rect 253204 4014 253256 4020
rect 252744 4004 252796 4010
rect 252744 3946 252796 3952
rect 253860 480 253888 9726
rect 253952 6225 253980 340054
rect 255056 335170 255084 340068
rect 254124 335164 254176 335170
rect 254124 335106 254176 335112
rect 255044 335164 255096 335170
rect 255044 335106 255096 335112
rect 254136 331106 254164 335106
rect 255700 334286 255728 340068
rect 255884 340054 256358 340082
rect 256804 340054 256910 340082
rect 255688 334280 255740 334286
rect 255688 334222 255740 334228
rect 255884 331242 255912 340054
rect 255964 337340 256016 337346
rect 255964 337282 256016 337288
rect 255516 331214 255912 331242
rect 254136 331078 254256 331106
rect 254228 321314 254256 331078
rect 254136 321286 254256 321314
rect 254136 318730 254164 321286
rect 254136 318702 254256 318730
rect 254228 298110 254256 318702
rect 255516 317506 255544 331214
rect 255424 317478 255544 317506
rect 255424 317422 255452 317478
rect 255412 317416 255464 317422
rect 255412 317358 255464 317364
rect 255596 317416 255648 317422
rect 255596 317358 255648 317364
rect 255608 316033 255636 317358
rect 255594 316024 255650 316033
rect 255594 315959 255650 315968
rect 255778 316024 255834 316033
rect 255778 315959 255834 315968
rect 255792 307442 255820 315959
rect 255608 307414 255820 307442
rect 255608 298194 255636 307414
rect 255516 298166 255636 298194
rect 255516 298110 255544 298166
rect 254216 298104 254268 298110
rect 254216 298046 254268 298052
rect 254492 298104 254544 298110
rect 254492 298046 254544 298052
rect 255504 298104 255556 298110
rect 255504 298046 255556 298052
rect 254504 296721 254532 298046
rect 254306 296712 254362 296721
rect 254306 296647 254362 296656
rect 254490 296712 254546 296721
rect 254490 296647 254546 296656
rect 254320 288130 254348 296647
rect 255504 288448 255556 288454
rect 255504 288390 255556 288396
rect 254320 288102 254532 288130
rect 254504 278798 254532 288102
rect 254216 278792 254268 278798
rect 254216 278734 254268 278740
rect 254492 278792 254544 278798
rect 254492 278734 254544 278740
rect 254228 273358 254256 278734
rect 254216 273352 254268 273358
rect 255516 273306 255544 288390
rect 254216 273294 254268 273300
rect 255424 273278 255544 273306
rect 254124 273216 254176 273222
rect 254124 273158 254176 273164
rect 255424 273170 255452 273278
rect 254136 265690 254164 273158
rect 255424 273142 255544 273170
rect 254136 265662 254256 265690
rect 254228 260846 254256 265662
rect 255516 260846 255544 273142
rect 254032 260840 254084 260846
rect 254032 260782 254084 260788
rect 254216 260840 254268 260846
rect 254216 260782 254268 260788
rect 255504 260840 255556 260846
rect 255504 260782 255556 260788
rect 254044 259457 254072 260782
rect 255596 260772 255648 260778
rect 255596 260714 255648 260720
rect 254030 259448 254086 259457
rect 254030 259383 254086 259392
rect 254214 259448 254270 259457
rect 254214 259383 254270 259392
rect 254228 251122 254256 259383
rect 255608 253858 255636 260714
rect 255516 253830 255636 253858
rect 254032 251116 254084 251122
rect 254032 251058 254084 251064
rect 254216 251116 254268 251122
rect 254216 251058 254268 251064
rect 254044 241534 254072 251058
rect 254032 241528 254084 241534
rect 254030 241496 254032 241505
rect 254216 241528 254268 241534
rect 254084 241496 254086 241505
rect 254030 241431 254086 241440
rect 254214 241496 254216 241505
rect 254268 241496 254270 241505
rect 254214 241431 254270 241440
rect 254044 236586 254072 241431
rect 254044 236558 254164 236586
rect 254136 225010 254164 236558
rect 254124 225004 254176 225010
rect 254124 224946 254176 224952
rect 254216 224868 254268 224874
rect 254216 224810 254268 224816
rect 254228 217462 254256 224810
rect 254216 217456 254268 217462
rect 254216 217398 254268 217404
rect 254124 217388 254176 217394
rect 254124 217330 254176 217336
rect 254136 212514 254164 217330
rect 254136 212486 254348 212514
rect 254320 205578 254348 212486
rect 254228 205550 254348 205578
rect 254228 202858 254256 205550
rect 254228 202830 254348 202858
rect 254320 193254 254348 202830
rect 254124 193248 254176 193254
rect 254122 193216 254124 193225
rect 254308 193248 254360 193254
rect 254176 193216 254178 193225
rect 254122 193151 254178 193160
rect 254306 193216 254308 193225
rect 254360 193216 254362 193225
rect 254306 193151 254362 193160
rect 254320 183598 254348 193151
rect 254308 183592 254360 183598
rect 254308 183534 254360 183540
rect 254216 183524 254268 183530
rect 254216 183466 254268 183472
rect 254228 177342 254256 183466
rect 254216 177336 254268 177342
rect 254216 177278 254268 177284
rect 255516 176746 255544 253830
rect 255424 176718 255544 176746
rect 255424 176610 255452 176718
rect 255424 176582 255544 176610
rect 254124 172576 254176 172582
rect 254124 172518 254176 172524
rect 254136 164218 254164 172518
rect 255516 164218 255544 176582
rect 254124 164212 254176 164218
rect 254124 164154 254176 164160
rect 254308 164212 254360 164218
rect 254308 164154 254360 164160
rect 255504 164212 255556 164218
rect 255504 164154 255556 164160
rect 255596 164212 255648 164218
rect 255596 164154 255648 164160
rect 254320 154601 254348 164154
rect 255608 157332 255636 164154
rect 255516 157304 255636 157332
rect 254306 154592 254362 154601
rect 254306 154527 254362 154536
rect 254306 154456 254362 154465
rect 254306 154391 254362 154400
rect 254320 147506 254348 154391
rect 254228 147478 254348 147506
rect 254228 144906 254256 147478
rect 254216 144900 254268 144906
rect 254216 144842 254268 144848
rect 254308 144900 254360 144906
rect 254308 144842 254360 144848
rect 254320 135289 254348 144842
rect 255516 138122 255544 157304
rect 255424 138094 255544 138122
rect 255424 137714 255452 138094
rect 255424 137686 255544 137714
rect 254122 135280 254178 135289
rect 254122 135215 254178 135224
rect 254306 135280 254362 135289
rect 254306 135215 254362 135224
rect 254136 130370 254164 135215
rect 254136 130342 254256 130370
rect 254228 125594 254256 130342
rect 255516 125594 255544 137686
rect 254216 125588 254268 125594
rect 254216 125530 254268 125536
rect 254308 125588 254360 125594
rect 254308 125530 254360 125536
rect 255504 125588 255556 125594
rect 255504 125530 255556 125536
rect 255596 125588 255648 125594
rect 255596 125530 255648 125536
rect 254320 115977 254348 125530
rect 255608 118674 255636 125530
rect 255516 118646 255636 118674
rect 254122 115968 254178 115977
rect 254122 115903 254124 115912
rect 254176 115903 254178 115912
rect 254306 115968 254362 115977
rect 254306 115903 254362 115912
rect 254124 115874 254176 115880
rect 254124 108996 254176 109002
rect 254124 108938 254176 108944
rect 254136 106298 254164 108938
rect 254136 106282 254256 106298
rect 254124 106276 254268 106282
rect 254176 106270 254216 106276
rect 254124 106218 254176 106224
rect 254216 106218 254268 106224
rect 254136 86902 254164 106218
rect 254124 86896 254176 86902
rect 254124 86838 254176 86844
rect 254124 77308 254176 77314
rect 254124 77250 254176 77256
rect 254136 48414 254164 77250
rect 255516 60738 255544 118646
rect 255424 60710 255544 60738
rect 255424 60602 255452 60710
rect 255424 60574 255544 60602
rect 255516 56574 255544 60574
rect 255504 56568 255556 56574
rect 255504 56510 255556 56516
rect 254124 48408 254176 48414
rect 254124 48350 254176 48356
rect 254216 48340 254268 48346
rect 254216 48282 254268 48288
rect 254228 41562 254256 48282
rect 255412 46980 255464 46986
rect 255412 46922 255464 46928
rect 255424 44878 255452 46922
rect 255412 44872 255464 44878
rect 255412 44814 255464 44820
rect 254228 41534 254348 41562
rect 254320 39386 254348 41534
rect 254228 39358 254348 39386
rect 254228 28966 254256 39358
rect 254032 28960 254084 28966
rect 254032 28902 254084 28908
rect 254216 28960 254268 28966
rect 254216 28902 254268 28908
rect 254044 19394 254072 28902
rect 255320 27600 255372 27606
rect 255320 27542 255372 27548
rect 255332 19394 255360 27542
rect 254044 19366 254164 19394
rect 255332 19366 255452 19394
rect 254136 9704 254164 19366
rect 255424 12458 255452 19366
rect 255424 12430 255544 12458
rect 255516 9704 255544 12430
rect 254044 9676 254164 9704
rect 255332 9676 255544 9704
rect 254044 8158 254072 9676
rect 254032 8152 254084 8158
rect 254032 8094 254084 8100
rect 253938 6216 253994 6225
rect 255332 6186 255360 9676
rect 253938 6151 253994 6160
rect 255320 6180 255372 6186
rect 255320 6122 255372 6128
rect 255976 4146 256004 337282
rect 256804 8226 256832 340054
rect 257540 337958 257568 340068
rect 258198 340054 258304 340082
rect 257528 337952 257580 337958
rect 257528 337894 257580 337900
rect 257344 337408 257396 337414
rect 257344 337350 257396 337356
rect 256792 8220 256844 8226
rect 256792 8162 256844 8168
rect 256240 7948 256292 7954
rect 256240 7890 256292 7896
rect 255964 4140 256016 4146
rect 255964 4082 256016 4088
rect 255044 3868 255096 3874
rect 255044 3810 255096 3816
rect 255056 480 255084 3810
rect 256252 480 256280 7890
rect 257356 3398 257384 337350
rect 257436 9716 257488 9722
rect 257436 9658 257488 9664
rect 257344 3392 257396 3398
rect 257344 3334 257396 3340
rect 257448 480 257476 9658
rect 258276 6254 258304 340054
rect 258368 340054 258750 340082
rect 258368 8294 258396 340054
rect 258724 337748 258776 337754
rect 258724 337690 258776 337696
rect 258356 8288 258408 8294
rect 258356 8230 258408 8236
rect 258264 6248 258316 6254
rect 258264 6190 258316 6196
rect 258632 3936 258684 3942
rect 258632 3878 258684 3884
rect 258644 480 258672 3878
rect 258736 3330 258764 337690
rect 259380 337346 259408 340068
rect 259472 340054 260038 340082
rect 260300 340054 260590 340082
rect 259368 337340 259420 337346
rect 259368 337282 259420 337288
rect 259366 277400 259422 277409
rect 259366 277335 259422 277344
rect 259380 267782 259408 277335
rect 259368 267776 259420 267782
rect 259368 267718 259420 267724
rect 259366 170368 259422 170377
rect 259366 170303 259422 170312
rect 259380 169969 259408 170303
rect 259366 169960 259422 169969
rect 259366 169895 259422 169904
rect 259472 6322 259500 340054
rect 260300 335646 260328 340054
rect 261220 338026 261248 340068
rect 261208 338020 261260 338026
rect 261208 337962 261260 337968
rect 259644 335640 259696 335646
rect 259644 335582 259696 335588
rect 260288 335640 260340 335646
rect 261312 335594 261340 340190
rect 262324 340054 262430 340082
rect 261484 337476 261536 337482
rect 261484 337418 261536 337424
rect 260288 335582 260340 335588
rect 259656 331106 259684 335582
rect 261036 335566 261340 335594
rect 259656 331078 259776 331106
rect 259748 321638 259776 331078
rect 261036 321706 261064 335566
rect 261024 321700 261076 321706
rect 261024 321642 261076 321648
rect 259736 321632 259788 321638
rect 259736 321574 259788 321580
rect 261024 321564 261076 321570
rect 261024 321506 261076 321512
rect 261036 319025 261064 321506
rect 261022 319016 261078 319025
rect 261022 318951 261078 318960
rect 261022 318880 261078 318889
rect 259644 318844 259696 318850
rect 261022 318815 261078 318824
rect 259644 318786 259696 318792
rect 259656 318730 259684 318786
rect 259656 318702 259776 318730
rect 259748 292618 259776 318702
rect 261036 311930 261064 318815
rect 261036 311902 261156 311930
rect 261128 307834 261156 311902
rect 261024 307828 261076 307834
rect 261024 307770 261076 307776
rect 261116 307828 261168 307834
rect 261116 307770 261168 307776
rect 261036 307737 261064 307770
rect 261022 307728 261078 307737
rect 261022 307663 261078 307672
rect 261206 307728 261262 307737
rect 261206 307663 261262 307672
rect 261220 298178 261248 307663
rect 261024 298172 261076 298178
rect 261024 298114 261076 298120
rect 261208 298172 261260 298178
rect 261208 298114 261260 298120
rect 261036 298042 261064 298114
rect 261024 298036 261076 298042
rect 261024 297978 261076 297984
rect 261116 298036 261168 298042
rect 261116 297978 261168 297984
rect 259656 292590 259776 292618
rect 259656 289814 259684 292590
rect 261128 292482 261156 297978
rect 261036 292454 261156 292482
rect 259644 289808 259696 289814
rect 259644 289750 259696 289756
rect 259736 282804 259788 282810
rect 259736 282746 259788 282752
rect 259748 277409 259776 282746
rect 261036 280140 261064 292454
rect 260852 280112 261064 280140
rect 259734 277400 259790 277409
rect 259734 277335 259790 277344
rect 260852 272898 260880 280112
rect 260852 272870 261064 272898
rect 259552 267776 259604 267782
rect 259552 267718 259604 267724
rect 259564 259457 259592 267718
rect 259550 259448 259606 259457
rect 259550 259383 259606 259392
rect 259734 259448 259790 259457
rect 259734 259383 259790 259392
rect 259748 249830 259776 259383
rect 261036 253994 261064 272870
rect 260944 253966 261064 253994
rect 260944 253858 260972 253966
rect 260944 253830 261064 253858
rect 259552 249824 259604 249830
rect 259552 249766 259604 249772
rect 259736 249824 259788 249830
rect 259736 249766 259788 249772
rect 259564 241534 259592 249766
rect 259552 241528 259604 241534
rect 259550 241496 259552 241505
rect 259736 241528 259788 241534
rect 259604 241496 259606 241505
rect 259550 241431 259606 241440
rect 259734 241496 259736 241505
rect 259788 241496 259790 241505
rect 261036 241482 261064 253830
rect 261036 241454 261156 241482
rect 259734 241431 259790 241440
rect 259564 236586 259592 241431
rect 259564 236558 259684 236586
rect 259656 231810 259684 236558
rect 261128 234666 261156 241454
rect 261116 234660 261168 234666
rect 261116 234602 261168 234608
rect 261024 234592 261076 234598
rect 261024 234534 261076 234540
rect 259644 231804 259696 231810
rect 259644 231746 259696 231752
rect 259736 222216 259788 222222
rect 259736 222158 259788 222164
rect 259748 217462 259776 222158
rect 259736 217456 259788 217462
rect 259736 217398 259788 217404
rect 259644 217388 259696 217394
rect 259644 217330 259696 217336
rect 259656 205698 259684 217330
rect 261036 215370 261064 234534
rect 260944 215342 261064 215370
rect 260944 215234 260972 215342
rect 260944 215206 261064 215234
rect 259644 205692 259696 205698
rect 259644 205634 259696 205640
rect 259736 205556 259788 205562
rect 259736 205498 259788 205504
rect 259748 193254 259776 205498
rect 261036 202858 261064 215206
rect 261036 202830 261156 202858
rect 261128 196042 261156 202830
rect 261116 196036 261168 196042
rect 261116 195978 261168 195984
rect 261024 195968 261076 195974
rect 261024 195910 261076 195916
rect 259736 193248 259788 193254
rect 259736 193190 259788 193196
rect 259644 193180 259696 193186
rect 259644 193122 259696 193128
rect 259656 182345 259684 193122
rect 261036 183546 261064 195910
rect 260852 183518 261064 183546
rect 259642 182336 259698 182345
rect 259642 182271 259698 182280
rect 259734 182200 259790 182209
rect 259734 182135 259736 182144
rect 259788 182135 259790 182144
rect 259920 182164 259972 182170
rect 259736 182106 259788 182112
rect 259920 182106 259972 182112
rect 259932 172553 259960 182106
rect 260852 176338 260880 183518
rect 260852 176310 261064 176338
rect 259642 172544 259698 172553
rect 259642 172479 259698 172488
rect 259918 172544 259974 172553
rect 259918 172479 259974 172488
rect 259656 164218 259684 172479
rect 259644 164212 259696 164218
rect 259644 164154 259696 164160
rect 261036 157434 261064 176310
rect 260944 157406 261064 157434
rect 260944 157298 260972 157406
rect 260944 157270 261064 157298
rect 259644 154624 259696 154630
rect 259644 154566 259696 154572
rect 259656 147694 259684 154566
rect 259644 147688 259696 147694
rect 259644 147630 259696 147636
rect 259736 147620 259788 147626
rect 259736 147562 259788 147568
rect 259748 144906 259776 147562
rect 259736 144900 259788 144906
rect 259736 144842 259788 144848
rect 259828 144900 259880 144906
rect 259828 144842 259880 144848
rect 259840 135289 259868 144842
rect 259642 135280 259698 135289
rect 259642 135215 259644 135224
rect 259696 135215 259698 135224
rect 259826 135280 259882 135289
rect 259826 135215 259828 135224
rect 259644 135186 259696 135192
rect 259880 135215 259882 135224
rect 259828 135186 259880 135192
rect 259840 125610 259868 135186
rect 259748 125594 259868 125610
rect 259736 125588 259880 125594
rect 259788 125582 259828 125588
rect 259736 125530 259788 125536
rect 259828 125530 259880 125536
rect 259840 115977 259868 125530
rect 261036 118794 261064 157270
rect 261024 118788 261076 118794
rect 261024 118730 261076 118736
rect 261024 118652 261076 118658
rect 261024 118594 261076 118600
rect 259642 115968 259698 115977
rect 259642 115903 259644 115912
rect 259696 115903 259698 115912
rect 259826 115968 259882 115977
rect 259826 115903 259828 115912
rect 259644 115874 259696 115880
rect 259880 115903 259882 115912
rect 259828 115874 259880 115880
rect 259840 96665 259868 115874
rect 261036 100094 261064 118594
rect 260840 100088 260892 100094
rect 260840 100030 260892 100036
rect 261024 100088 261076 100094
rect 261024 100030 261076 100036
rect 259642 96656 259698 96665
rect 259642 96591 259698 96600
rect 259826 96656 259882 96665
rect 259826 96591 259882 96600
rect 259656 86902 259684 96591
rect 260852 90522 260880 100030
rect 260760 90494 260880 90522
rect 259644 86896 259696 86902
rect 259644 86838 259696 86844
rect 260760 85678 260788 90494
rect 260748 85672 260800 85678
rect 260748 85614 260800 85620
rect 261024 85604 261076 85610
rect 261024 85546 261076 85552
rect 259644 77308 259696 77314
rect 259644 77250 259696 77256
rect 259656 59770 259684 77250
rect 261036 76022 261064 85546
rect 261024 76016 261076 76022
rect 261024 75958 261076 75964
rect 260840 75880 260892 75886
rect 260840 75822 260892 75828
rect 260852 66366 260880 75822
rect 260840 66360 260892 66366
rect 260840 66302 260892 66308
rect 261024 66360 261076 66366
rect 261024 66302 261076 66308
rect 261036 64870 261064 66302
rect 261024 64864 261076 64870
rect 261024 64806 261076 64812
rect 259644 59764 259696 59770
rect 259644 59706 259696 59712
rect 260840 55276 260892 55282
rect 260840 55218 260892 55224
rect 260852 51626 260880 55218
rect 260852 51598 261156 51626
rect 259736 48340 259788 48346
rect 259736 48282 259788 48288
rect 259748 28966 259776 48282
rect 261128 46866 261156 51598
rect 260944 46838 261156 46866
rect 260944 40610 260972 46838
rect 260944 40582 261064 40610
rect 261036 33810 261064 40582
rect 260944 33782 261064 33810
rect 259736 28960 259788 28966
rect 259736 28902 259788 28908
rect 259828 28960 259880 28966
rect 259828 28902 259880 28908
rect 259840 27606 259868 28902
rect 259828 27600 259880 27606
rect 259828 27542 259880 27548
rect 260944 19378 260972 33782
rect 260932 19372 260984 19378
rect 260932 19314 260984 19320
rect 261024 19372 261076 19378
rect 261024 19314 261076 19320
rect 259828 18012 259880 18018
rect 259828 17954 259880 17960
rect 259840 10305 259868 17954
rect 261036 12578 261064 19314
rect 261024 12572 261076 12578
rect 261024 12514 261076 12520
rect 260932 11756 260984 11762
rect 260932 11698 260984 11704
rect 259826 10296 259882 10305
rect 259826 10231 259882 10240
rect 259828 8016 259880 8022
rect 259828 7958 259880 7964
rect 259460 6316 259512 6322
rect 259460 6258 259512 6264
rect 258724 3324 258776 3330
rect 258724 3266 258776 3272
rect 259840 480 259868 7958
rect 260944 6458 260972 11698
rect 260932 6452 260984 6458
rect 260932 6394 260984 6400
rect 261024 3460 261076 3466
rect 261024 3402 261076 3408
rect 261036 480 261064 3402
rect 261496 3262 261524 337418
rect 262324 10334 262352 340054
rect 262864 337544 262916 337550
rect 262864 337486 262916 337492
rect 262312 10328 262364 10334
rect 262312 10270 262364 10276
rect 262220 4072 262272 4078
rect 262220 4014 262272 4020
rect 261484 3256 261536 3262
rect 261484 3198 261536 3204
rect 262232 480 262260 4014
rect 262876 3194 262904 337486
rect 263060 337414 263088 340068
rect 263048 337408 263100 337414
rect 263048 337350 263100 337356
rect 263416 8084 263468 8090
rect 263416 8026 263468 8032
rect 262864 3188 262916 3194
rect 262864 3130 262916 3136
rect 263428 480 263456 8026
rect 263704 6390 263732 340068
rect 263796 340054 264270 340082
rect 263692 6384 263744 6390
rect 263692 6326 263744 6332
rect 263796 5302 263824 340054
rect 264900 338094 264928 340068
rect 264992 340054 265466 340082
rect 264888 338088 264940 338094
rect 264888 338030 264940 338036
rect 264336 337680 264388 337686
rect 264336 337622 264388 337628
rect 264244 337476 264296 337482
rect 264244 337418 264296 337424
rect 263784 5296 263836 5302
rect 263784 5238 263836 5244
rect 264256 3126 264284 337418
rect 264244 3120 264296 3126
rect 264244 3062 264296 3068
rect 264348 3058 264376 337622
rect 264992 6526 265020 340054
rect 265544 328506 265572 340190
rect 266740 337754 266768 340068
rect 266728 337748 266780 337754
rect 266728 337690 266780 337696
rect 266832 331242 266860 340190
rect 266556 331214 266860 331242
rect 267844 340054 267950 340082
rect 265256 328500 265308 328506
rect 265256 328442 265308 328448
rect 265532 328500 265584 328506
rect 265532 328442 265584 328448
rect 265268 311930 265296 328442
rect 266556 321586 266584 331214
rect 267096 328500 267148 328506
rect 267096 328442 267148 328448
rect 266464 321558 266584 321586
rect 266464 321450 266492 321558
rect 266464 321422 266584 321450
rect 265176 311902 265296 311930
rect 265176 299538 265204 311902
rect 265164 299532 265216 299538
rect 265164 299474 265216 299480
rect 265256 299532 265308 299538
rect 265256 299474 265308 299480
rect 265268 298110 265296 299474
rect 265256 298104 265308 298110
rect 265256 298046 265308 298052
rect 266556 292618 266584 321422
rect 267108 309194 267136 328442
rect 267096 309188 267148 309194
rect 267096 309130 267148 309136
rect 267096 307828 267148 307834
rect 267096 307770 267148 307776
rect 267108 298110 267136 307770
rect 267096 298104 267148 298110
rect 267096 298046 267148 298052
rect 266464 292590 266584 292618
rect 266464 292482 266492 292590
rect 266464 292454 266584 292482
rect 265256 288448 265308 288454
rect 265256 288390 265308 288396
rect 265268 284866 265296 288390
rect 265268 284838 265388 284866
rect 265360 282826 265388 284838
rect 265268 282798 265388 282826
rect 265268 280158 265296 282798
rect 265164 280152 265216 280158
rect 265164 280094 265216 280100
rect 265256 280152 265308 280158
rect 266556 280140 266584 292454
rect 267004 280220 267056 280226
rect 267004 280162 267056 280168
rect 265256 280094 265308 280100
rect 266372 280112 266584 280140
rect 265176 269113 265204 280094
rect 266372 272762 266400 280112
rect 266372 272734 266584 272762
rect 265162 269104 265218 269113
rect 265162 269039 265218 269048
rect 265438 269104 265494 269113
rect 265438 269039 265494 269048
rect 265452 253994 265480 269039
rect 266556 253994 266584 272734
rect 267016 270570 267044 280162
rect 267004 270564 267056 270570
rect 267004 270506 267056 270512
rect 267096 270564 267148 270570
rect 267096 270506 267148 270512
rect 267108 269090 267136 270506
rect 267016 269062 267136 269090
rect 267016 263634 267044 269062
rect 267004 263628 267056 263634
rect 267004 263570 267056 263576
rect 267004 259480 267056 259486
rect 267004 259422 267056 259428
rect 267016 254538 267044 259422
rect 265268 253966 265480 253994
rect 266464 253966 266584 253994
rect 266832 254510 267044 254538
rect 265268 230586 265296 253966
rect 266464 253858 266492 253966
rect 266464 253830 266584 253858
rect 265164 230580 265216 230586
rect 265164 230522 265216 230528
rect 265256 230580 265308 230586
rect 265256 230522 265308 230528
rect 265176 230489 265204 230522
rect 265162 230480 265218 230489
rect 265162 230415 265218 230424
rect 265346 230480 265402 230489
rect 265346 230415 265402 230424
rect 265360 224874 265388 230415
rect 265164 224868 265216 224874
rect 265164 224810 265216 224816
rect 265348 224868 265400 224874
rect 265348 224810 265400 224816
rect 265176 209778 265204 224810
rect 266556 215370 266584 253830
rect 266832 238082 266860 254510
rect 266832 238054 267136 238082
rect 267108 225010 267136 238054
rect 267096 225004 267148 225010
rect 267096 224946 267148 224952
rect 267096 220856 267148 220862
rect 267096 220798 267148 220804
rect 267108 219434 267136 220798
rect 267096 219428 267148 219434
rect 267096 219370 267148 219376
rect 266464 215342 266584 215370
rect 266464 215234 266492 215342
rect 266464 215206 266584 215234
rect 265164 209772 265216 209778
rect 265164 209714 265216 209720
rect 266556 202881 266584 215206
rect 267004 209840 267056 209846
rect 267004 209782 267056 209788
rect 266358 202872 266414 202881
rect 265256 202836 265308 202842
rect 266358 202807 266414 202816
rect 266542 202872 266598 202881
rect 267016 202858 267044 209782
rect 267016 202830 267136 202858
rect 266542 202807 266598 202816
rect 265256 202778 265308 202784
rect 265268 200138 265296 202778
rect 265268 200110 265388 200138
rect 265360 193322 265388 200110
rect 265164 193316 265216 193322
rect 265164 193258 265216 193264
rect 265348 193316 265400 193322
rect 265348 193258 265400 193264
rect 265176 193202 265204 193258
rect 266372 193254 266400 202807
rect 267108 202722 267136 202830
rect 267016 202694 267136 202722
rect 267016 193254 267044 202694
rect 266360 193248 266412 193254
rect 265176 193174 265296 193202
rect 266360 193190 266412 193196
rect 266544 193248 266596 193254
rect 266544 193190 266596 193196
rect 267004 193248 267056 193254
rect 267004 193190 267056 193196
rect 267096 193248 267148 193254
rect 267096 193190 267148 193196
rect 265268 174078 265296 193174
rect 266556 191826 266584 193190
rect 266544 191820 266596 191826
rect 266544 191762 266596 191768
rect 267108 186454 267136 193190
rect 267096 186448 267148 186454
rect 267096 186390 267148 186396
rect 267004 186312 267056 186318
rect 267004 186254 267056 186260
rect 267016 183569 267044 186254
rect 267002 183560 267058 183569
rect 267002 183495 267058 183504
rect 267186 183560 267242 183569
rect 267186 183495 267242 183504
rect 266452 183388 266504 183394
rect 266452 183330 266504 183336
rect 265256 174072 265308 174078
rect 265256 174014 265308 174020
rect 265256 173936 265308 173942
rect 265176 173896 265256 173924
rect 265176 164393 265204 173896
rect 265256 173878 265308 173884
rect 266464 171034 266492 183330
rect 267200 173924 267228 183495
rect 267108 173896 267228 173924
rect 266464 171006 266584 171034
rect 265162 164384 265218 164393
rect 265162 164319 265218 164328
rect 265254 164248 265310 164257
rect 265254 164183 265310 164192
rect 265268 161430 265296 164183
rect 265256 161424 265308 161430
rect 265256 161366 265308 161372
rect 266556 157434 266584 171006
rect 267108 164234 267136 173896
rect 267738 169960 267794 169969
rect 267738 169895 267740 169904
rect 267792 169895 267794 169904
rect 267740 169866 267792 169872
rect 267016 164206 267136 164234
rect 267016 157486 267044 164206
rect 266464 157406 266584 157434
rect 267004 157480 267056 157486
rect 267004 157422 267056 157428
rect 266464 157298 266492 157406
rect 266464 157270 266584 157298
rect 265256 151836 265308 151842
rect 265256 151778 265308 151784
rect 265268 143585 265296 151778
rect 265254 143576 265310 143585
rect 266556 143562 266584 157270
rect 267004 153196 267056 153202
rect 267004 153138 267056 153144
rect 267016 143614 267044 153138
rect 265254 143511 265310 143520
rect 266464 143534 266584 143562
rect 267004 143608 267056 143614
rect 267004 143550 267056 143556
rect 267096 143608 267148 143614
rect 267096 143550 267148 143556
rect 265438 143440 265494 143449
rect 265438 143375 265494 143384
rect 265452 132546 265480 143375
rect 266464 142118 266492 143534
rect 266452 142112 266504 142118
rect 266452 142054 266504 142060
rect 267108 133906 267136 143550
rect 265360 132518 265480 132546
rect 267016 133878 267136 133906
rect 266544 132524 266596 132530
rect 265360 132462 265388 132518
rect 266544 132466 266596 132472
rect 265348 132456 265400 132462
rect 265348 132398 265400 132404
rect 266556 125594 266584 132466
rect 267016 125594 267044 133878
rect 266544 125588 266596 125594
rect 266544 125530 266596 125536
rect 266728 125588 266780 125594
rect 266728 125530 266780 125536
rect 267004 125588 267056 125594
rect 267004 125530 267056 125536
rect 267280 125588 267332 125594
rect 267280 125530 267332 125536
rect 265348 124636 265400 124642
rect 265348 124578 265400 124584
rect 265360 115977 265388 124578
rect 266740 115977 266768 125530
rect 267292 115977 267320 125530
rect 265162 115968 265218 115977
rect 265346 115968 265402 115977
rect 265162 115903 265164 115912
rect 265216 115903 265218 115912
rect 265256 115932 265308 115938
rect 265164 115874 265216 115880
rect 265346 115903 265402 115912
rect 266726 115968 266782 115977
rect 266726 115903 266782 115912
rect 267094 115968 267150 115977
rect 267094 115903 267150 115912
rect 267278 115968 267334 115977
rect 267278 115903 267334 115912
rect 265256 115874 265308 115880
rect 265268 95282 265296 115874
rect 266542 115832 266598 115841
rect 266542 115767 266598 115776
rect 266556 99498 266584 115767
rect 267108 114510 267136 115903
rect 267096 114504 267148 114510
rect 267096 114446 267148 114452
rect 267004 104984 267056 104990
rect 267004 104926 267056 104932
rect 267016 104854 267044 104926
rect 267004 104848 267056 104854
rect 267004 104790 267056 104796
rect 266556 99470 266676 99498
rect 266648 97322 266676 99470
rect 265176 95254 265296 95282
rect 266556 97294 266676 97322
rect 265176 95198 265204 95254
rect 265164 95192 265216 95198
rect 265164 95134 265216 95140
rect 265164 85604 265216 85610
rect 265164 85546 265216 85552
rect 265176 77194 265204 85546
rect 265176 77166 265296 77194
rect 265268 72978 265296 77166
rect 265268 72950 265388 72978
rect 265360 48346 265388 72950
rect 266556 70514 266584 97294
rect 267096 95260 267148 95266
rect 267096 95202 267148 95208
rect 267108 85626 267136 95202
rect 267016 85598 267136 85626
rect 267016 79370 267044 85598
rect 267016 79342 267136 79370
rect 267108 74594 267136 79342
rect 267096 74588 267148 74594
rect 267096 74530 267148 74536
rect 267280 74588 267332 74594
rect 267280 74530 267332 74536
rect 266544 70508 266596 70514
rect 266544 70450 266596 70456
rect 266452 70372 266504 70378
rect 266452 70314 266504 70320
rect 266464 58002 266492 70314
rect 267292 67726 267320 74530
rect 267280 67720 267332 67726
rect 267280 67662 267332 67668
rect 267188 67584 267240 67590
rect 267188 67526 267240 67532
rect 267200 58002 267228 67526
rect 266452 57996 266504 58002
rect 266452 57938 266504 57944
rect 266544 57996 266596 58002
rect 266544 57938 266596 57944
rect 267096 57996 267148 58002
rect 267096 57938 267148 57944
rect 267188 57996 267240 58002
rect 267188 57938 267240 57944
rect 266556 48362 266584 57938
rect 265164 48340 265216 48346
rect 265164 48282 265216 48288
rect 265348 48340 265400 48346
rect 265348 48282 265400 48288
rect 266464 48334 266584 48362
rect 265176 38434 265204 48282
rect 266464 42106 266492 48334
rect 267108 47002 267136 57938
rect 267016 46974 267136 47002
rect 267016 46918 267044 46974
rect 267004 46912 267056 46918
rect 267004 46854 267056 46860
rect 267188 46912 267240 46918
rect 267188 46854 267240 46860
rect 267200 45558 267228 46854
rect 267188 45552 267240 45558
rect 267188 45494 267240 45500
rect 266464 42078 266584 42106
rect 265176 38406 265296 38434
rect 265268 28966 265296 38406
rect 266556 28966 266584 42078
rect 267004 35964 267056 35970
rect 267004 35906 267056 35912
rect 265164 28960 265216 28966
rect 265164 28902 265216 28908
rect 265256 28960 265308 28966
rect 265256 28902 265308 28908
rect 266360 28960 266412 28966
rect 266360 28902 266412 28908
rect 266544 28960 266596 28966
rect 266544 28902 266596 28908
rect 265176 14550 265204 28902
rect 266372 19394 266400 28902
rect 267016 27606 267044 35906
rect 267004 27600 267056 27606
rect 267004 27542 267056 27548
rect 267096 27600 267148 27606
rect 267096 27542 267148 27548
rect 266372 19366 266492 19394
rect 265164 14544 265216 14550
rect 266464 14498 266492 19366
rect 265164 14486 265216 14492
rect 266280 14470 266492 14498
rect 266280 12322 266308 14470
rect 266280 12294 266400 12322
rect 266372 6594 266400 12294
rect 267108 9602 267136 27542
rect 267844 14618 267872 340054
rect 268384 337884 268436 337890
rect 268384 337826 268436 337832
rect 267832 14612 267884 14618
rect 267832 14554 267884 14560
rect 266924 9574 267136 9602
rect 266360 6588 266412 6594
rect 266360 6530 266412 6536
rect 264980 6520 265032 6526
rect 264980 6462 265032 6468
rect 264612 3732 264664 3738
rect 264612 3674 264664 3680
rect 264336 3052 264388 3058
rect 264336 2994 264388 3000
rect 264624 480 264652 3674
rect 265808 3528 265860 3534
rect 265808 3470 265860 3476
rect 265820 480 265848 3470
rect 266924 2990 266952 9574
rect 267004 8152 267056 8158
rect 267004 8094 267056 8100
rect 266912 2984 266964 2990
rect 266912 2926 266964 2932
rect 267016 480 267044 8094
rect 268108 3392 268160 3398
rect 268108 3334 268160 3340
rect 268120 480 268148 3334
rect 268396 2922 268424 337826
rect 268580 336802 268608 340068
rect 268568 336796 268620 336802
rect 268568 336738 268620 336744
rect 269026 17232 269082 17241
rect 269026 17167 269082 17176
rect 269040 16833 269068 17167
rect 269026 16824 269082 16833
rect 269026 16759 269082 16768
rect 269132 6662 269160 340068
rect 269224 340054 269790 340082
rect 269224 14686 269252 340054
rect 269764 337816 269816 337822
rect 269764 337758 269816 337764
rect 269212 14680 269264 14686
rect 269212 14622 269264 14628
rect 269120 6656 269172 6662
rect 269120 6598 269172 6604
rect 269304 3664 269356 3670
rect 269304 3606 269356 3612
rect 268384 2916 268436 2922
rect 268384 2858 268436 2864
rect 269316 480 269344 3606
rect 269776 2854 269804 337758
rect 270420 337346 270448 340068
rect 270512 340054 270986 340082
rect 270408 337340 270460 337346
rect 270408 337282 270460 337288
rect 270408 191820 270460 191826
rect 270408 191762 270460 191768
rect 270420 182209 270448 191762
rect 270406 182200 270462 182209
rect 270406 182135 270462 182144
rect 270512 9602 270540 340054
rect 271064 328506 271092 340190
rect 272260 337278 272288 340068
rect 272248 337272 272300 337278
rect 272248 337214 272300 337220
rect 272352 335594 272380 340190
rect 272076 335566 272380 335594
rect 273364 340054 273470 340082
rect 270776 328500 270828 328506
rect 270776 328442 270828 328448
rect 271052 328500 271104 328506
rect 271052 328442 271104 328448
rect 270788 311930 270816 328442
rect 272076 321586 272104 335566
rect 271984 321558 272104 321586
rect 271984 321450 272012 321558
rect 271984 321422 272104 321450
rect 270696 311902 270816 311930
rect 270696 309126 270724 311902
rect 270684 309120 270736 309126
rect 270684 309062 270736 309068
rect 270776 299532 270828 299538
rect 270776 299474 270828 299480
rect 270788 298110 270816 299474
rect 270776 298104 270828 298110
rect 270776 298046 270828 298052
rect 270868 298104 270920 298110
rect 270868 298046 270920 298052
rect 270880 280158 270908 298046
rect 272076 292618 272104 321422
rect 271984 292590 272104 292618
rect 271984 292482 272012 292590
rect 271984 292454 272104 292482
rect 270592 280152 270644 280158
rect 270592 280094 270644 280100
rect 270868 280152 270920 280158
rect 270868 280094 270920 280100
rect 270604 278730 270632 280094
rect 270592 278724 270644 278730
rect 270592 278666 270644 278672
rect 272076 273222 272104 292454
rect 272064 273216 272116 273222
rect 272064 273158 272116 273164
rect 272064 273080 272116 273086
rect 272064 273022 272116 273028
rect 270776 269136 270828 269142
rect 270776 269078 270828 269084
rect 270788 260817 270816 269078
rect 270774 260808 270830 260817
rect 270774 260743 270830 260752
rect 270590 260672 270646 260681
rect 270590 260607 270646 260616
rect 270604 251190 270632 260607
rect 272076 253910 272104 273022
rect 272064 253904 272116 253910
rect 272064 253846 272116 253852
rect 272064 253768 272116 253774
rect 272064 253710 272116 253716
rect 270592 251184 270644 251190
rect 270592 251126 270644 251132
rect 270960 251184 271012 251190
rect 270960 251126 271012 251132
rect 270972 231962 271000 251126
rect 272076 234598 272104 253710
rect 272064 234592 272116 234598
rect 272064 234534 272116 234540
rect 272064 234456 272116 234462
rect 272064 234398 272116 234404
rect 270788 231934 271000 231962
rect 270788 231826 270816 231934
rect 270788 231798 271000 231826
rect 270972 212566 271000 231798
rect 272076 215286 272104 234398
rect 272064 215280 272116 215286
rect 272064 215222 272116 215228
rect 272064 215144 272116 215150
rect 272064 215086 272116 215092
rect 270776 212560 270828 212566
rect 270776 212502 270828 212508
rect 270960 212560 271012 212566
rect 270960 212502 271012 212508
rect 270788 205714 270816 212502
rect 270604 205686 270816 205714
rect 270604 203153 270632 205686
rect 270590 203144 270646 203153
rect 270590 203079 270646 203088
rect 270774 203008 270830 203017
rect 270774 202943 270830 202952
rect 270788 196110 270816 202943
rect 270776 196104 270828 196110
rect 272076 196058 272104 215086
rect 270776 196046 270828 196052
rect 271984 196030 272104 196058
rect 271984 195922 272012 196030
rect 271984 195894 272104 195922
rect 270776 193180 270828 193186
rect 270776 193122 270828 193128
rect 270788 191826 270816 193122
rect 270776 191820 270828 191826
rect 270776 191762 270828 191768
rect 272076 188442 272104 195894
rect 271984 188414 272104 188442
rect 271984 183569 272012 188414
rect 271970 183560 272026 183569
rect 271970 183495 272026 183504
rect 272246 183424 272302 183433
rect 272246 183359 272302 183368
rect 270590 182200 270646 182209
rect 270590 182135 270592 182144
rect 270644 182135 270646 182144
rect 270868 182164 270920 182170
rect 270592 182106 270644 182112
rect 270868 182106 270920 182112
rect 270880 172553 270908 182106
rect 270682 172544 270738 172553
rect 270682 172479 270738 172488
rect 270866 172544 270922 172553
rect 270866 172479 270922 172488
rect 270696 167074 270724 172479
rect 270684 167068 270736 167074
rect 270684 167010 270736 167016
rect 270776 166932 270828 166938
rect 270776 166874 270828 166880
rect 270788 157570 270816 166874
rect 272260 164257 272288 183359
rect 272062 164248 272118 164257
rect 272062 164183 272064 164192
rect 272116 164183 272118 164192
rect 272246 164248 272302 164257
rect 272246 164183 272248 164192
rect 272064 164154 272116 164160
rect 272300 164183 272302 164192
rect 272248 164154 272300 164160
rect 270788 157542 270908 157570
rect 270880 154737 270908 157542
rect 270866 154728 270922 154737
rect 270866 154663 270922 154672
rect 272260 154601 272288 164154
rect 270682 154592 270738 154601
rect 272062 154592 272118 154601
rect 270682 154527 270684 154536
rect 270736 154527 270738 154536
rect 271788 154556 271840 154562
rect 270684 154498 270736 154504
rect 272062 154527 272064 154536
rect 271788 154498 271840 154504
rect 272116 154527 272118 154536
rect 272246 154592 272302 154601
rect 272246 154527 272302 154536
rect 272064 154498 272116 154504
rect 270684 147620 270736 147626
rect 270684 147562 270736 147568
rect 270696 144922 270724 147562
rect 271800 144945 271828 154498
rect 271786 144936 271842 144945
rect 270696 144894 270816 144922
rect 270788 138258 270816 144894
rect 271786 144871 271842 144880
rect 271970 144936 272026 144945
rect 271970 144871 271972 144880
rect 272024 144871 272026 144880
rect 272064 144900 272116 144906
rect 271972 144842 272024 144848
rect 272064 144842 272116 144848
rect 272076 139890 272104 144842
rect 271984 139862 272104 139890
rect 270788 138230 270908 138258
rect 270880 135289 270908 138230
rect 270682 135280 270738 135289
rect 270682 135215 270684 135224
rect 270736 135215 270738 135224
rect 270866 135280 270922 135289
rect 270866 135215 270922 135224
rect 270684 135186 270736 135192
rect 271984 130422 272012 139862
rect 271972 130416 272024 130422
rect 271972 130358 272024 130364
rect 272156 130416 272208 130422
rect 272156 130358 272208 130364
rect 270684 128308 270736 128314
rect 270684 128250 270736 128256
rect 270696 125610 270724 128250
rect 270696 125582 270816 125610
rect 270788 120766 270816 125582
rect 270776 120760 270828 120766
rect 270776 120702 270828 120708
rect 270776 120624 270828 120630
rect 270776 120566 270828 120572
rect 270788 111058 270816 120566
rect 272168 116006 272196 130358
rect 272064 116000 272116 116006
rect 272064 115942 272116 115948
rect 272156 116000 272208 116006
rect 272156 115942 272208 115948
rect 270788 111030 270908 111058
rect 270880 102134 270908 111030
rect 270868 102128 270920 102134
rect 270868 102070 270920 102076
rect 272076 96778 272104 115942
rect 271984 96750 272104 96778
rect 271984 96642 272012 96750
rect 271984 96614 272104 96642
rect 270960 92540 271012 92546
rect 270960 92482 271012 92488
rect 270972 82822 271000 92482
rect 272076 86970 272104 96614
rect 271972 86964 272024 86970
rect 271972 86906 272024 86912
rect 272064 86964 272116 86970
rect 272064 86906 272116 86912
rect 270960 82816 271012 82822
rect 270960 82758 271012 82764
rect 271984 73250 272012 86906
rect 271984 73222 272104 73250
rect 272076 73166 272104 73222
rect 272064 73160 272116 73166
rect 272064 73102 272116 73108
rect 270684 64932 270736 64938
rect 270684 64874 270736 64880
rect 270696 57594 270724 64874
rect 271972 63572 272024 63578
rect 271972 63514 272024 63520
rect 271984 58614 272012 63514
rect 271972 58608 272024 58614
rect 271972 58550 272024 58556
rect 270684 57588 270736 57594
rect 270684 57530 270736 57536
rect 270592 46980 270644 46986
rect 270592 46922 270644 46928
rect 270604 38706 270632 46922
rect 272064 45620 272116 45626
rect 272064 45562 272116 45568
rect 272076 38758 272104 45562
rect 273074 40352 273130 40361
rect 273258 40352 273314 40361
rect 273130 40310 273258 40338
rect 273074 40287 273130 40296
rect 273258 40287 273314 40296
rect 272064 38752 272116 38758
rect 270604 38678 270724 38706
rect 272064 38694 272116 38700
rect 270696 29102 270724 38678
rect 272064 37256 272116 37262
rect 272064 37198 272116 37204
rect 270684 29096 270736 29102
rect 270684 29038 270736 29044
rect 270776 29028 270828 29034
rect 270776 28970 270828 28976
rect 270788 22642 270816 28970
rect 272076 27606 272104 37198
rect 272064 27600 272116 27606
rect 272064 27542 272116 27548
rect 270776 22636 270828 22642
rect 270776 22578 270828 22584
rect 271972 18012 272024 18018
rect 271972 17954 272024 17960
rect 271984 14498 272012 17954
rect 273364 14822 273392 340054
rect 274100 336870 274128 340068
rect 274088 336864 274140 336870
rect 274088 336806 274140 336812
rect 273352 14816 273404 14822
rect 273352 14758 273404 14764
rect 271800 14470 272012 14498
rect 271800 12322 271828 14470
rect 271800 12294 271920 12322
rect 270512 9574 270632 9602
rect 270500 8220 270552 8226
rect 270500 8162 270552 8168
rect 269764 2848 269816 2854
rect 269764 2790 269816 2796
rect 270512 480 270540 8162
rect 270604 6730 270632 9574
rect 271892 6798 271920 12294
rect 274088 8288 274140 8294
rect 274088 8230 274140 8236
rect 271880 6792 271932 6798
rect 271880 6734 271932 6740
rect 270592 6724 270644 6730
rect 270592 6666 270644 6672
rect 271696 4004 271748 4010
rect 271696 3946 271748 3952
rect 271708 480 271736 3946
rect 272892 3800 272944 3806
rect 272892 3742 272944 3748
rect 272904 480 272932 3742
rect 274100 480 274128 8230
rect 274652 7546 274680 340068
rect 274744 340054 275310 340082
rect 274744 14890 274772 340054
rect 275940 337414 275968 340068
rect 276032 340054 276506 340082
rect 276584 340054 277150 340082
rect 275928 337408 275980 337414
rect 275928 337350 275980 337356
rect 274732 14884 274784 14890
rect 274732 14826 274784 14832
rect 274640 7540 274692 7546
rect 274640 7482 274692 7488
rect 276032 7478 276060 340054
rect 276584 335730 276612 340054
rect 276664 337408 276716 337414
rect 276664 337350 276716 337356
rect 276124 335702 276612 335730
rect 276124 14958 276152 335702
rect 276112 14952 276164 14958
rect 276112 14894 276164 14900
rect 276020 7472 276072 7478
rect 276020 7414 276072 7420
rect 276676 4146 276704 337350
rect 277780 337210 277808 340068
rect 277964 340054 278346 340082
rect 278884 340054 278990 340082
rect 277768 337204 277820 337210
rect 277768 337146 277820 337152
rect 277964 335345 277992 340054
rect 277674 335336 277730 335345
rect 277674 335271 277730 335280
rect 277950 335336 278006 335345
rect 277950 335271 278006 335280
rect 277688 325689 277716 335271
rect 277674 325680 277730 325689
rect 277674 325615 277730 325624
rect 277858 325680 277914 325689
rect 277858 325615 277914 325624
rect 277688 316062 277716 316093
rect 277872 316062 277900 325615
rect 277676 316056 277728 316062
rect 277596 316004 277676 316010
rect 277596 315998 277728 316004
rect 277860 316056 277912 316062
rect 277860 315998 277912 316004
rect 277596 315982 277716 315998
rect 277596 311914 277624 315982
rect 277584 311908 277636 311914
rect 277584 311850 277636 311856
rect 277584 306400 277636 306406
rect 277584 306342 277636 306348
rect 277596 299606 277624 306342
rect 277584 299600 277636 299606
rect 277584 299542 277636 299548
rect 277584 299464 277636 299470
rect 277584 299406 277636 299412
rect 277596 298110 277624 299406
rect 277584 298104 277636 298110
rect 277584 298046 277636 298052
rect 277676 280220 277728 280226
rect 277676 280162 277728 280168
rect 277688 275126 277716 280162
rect 277676 275120 277728 275126
rect 277676 275062 277728 275068
rect 277768 269136 277820 269142
rect 277768 269078 277820 269084
rect 277780 265554 277808 269078
rect 277596 265526 277808 265554
rect 277596 260846 277624 265526
rect 277584 260840 277636 260846
rect 277584 260782 277636 260788
rect 277676 260840 277728 260846
rect 277676 260782 277728 260788
rect 277688 244202 277716 260782
rect 277596 244174 277716 244202
rect 277596 231878 277624 244174
rect 277584 231872 277636 231878
rect 277584 231814 277636 231820
rect 277676 231872 277728 231878
rect 277676 231814 277728 231820
rect 277688 224890 277716 231814
rect 277596 224862 277716 224890
rect 277596 212566 277624 224862
rect 277584 212560 277636 212566
rect 277584 212502 277636 212508
rect 277676 212560 277728 212566
rect 277676 212502 277728 212508
rect 277688 205578 277716 212502
rect 277596 205550 277716 205578
rect 277596 196058 277624 205550
rect 277504 196030 277624 196058
rect 277504 195974 277532 196030
rect 277492 195968 277544 195974
rect 277492 195910 277544 195916
rect 277676 195968 277728 195974
rect 277676 195910 277728 195916
rect 277688 183598 277716 195910
rect 277584 183592 277636 183598
rect 277584 183534 277636 183540
rect 277676 183592 277728 183598
rect 277676 183534 277728 183540
rect 277596 176662 277624 183534
rect 277584 176656 277636 176662
rect 277584 176598 277636 176604
rect 277584 176520 277636 176526
rect 277584 176462 277636 176468
rect 277596 166954 277624 176462
rect 278688 169924 278740 169930
rect 278688 169866 278740 169872
rect 278700 169833 278728 169866
rect 278686 169824 278742 169833
rect 278686 169759 278742 169768
rect 277412 166926 277624 166954
rect 277412 154601 277440 166926
rect 277398 154592 277454 154601
rect 277398 154527 277454 154536
rect 277674 154592 277730 154601
rect 277674 154527 277730 154536
rect 277688 147642 277716 154527
rect 277596 147614 277716 147642
rect 277596 138106 277624 147614
rect 277584 138100 277636 138106
rect 277584 138042 277636 138048
rect 277584 137964 277636 137970
rect 277584 137906 277636 137912
rect 277596 118538 277624 137906
rect 277596 118510 277716 118538
rect 277688 109018 277716 118510
rect 277596 108990 277716 109018
rect 277596 99414 277624 108990
rect 277584 99408 277636 99414
rect 277584 99350 277636 99356
rect 277676 99340 277728 99346
rect 277676 99282 277728 99288
rect 277688 89706 277716 99282
rect 277504 89678 277716 89706
rect 277504 80170 277532 89678
rect 277492 80164 277544 80170
rect 277492 80106 277544 80112
rect 277400 80028 277452 80034
rect 277400 79970 277452 79976
rect 277412 77246 277440 79970
rect 277400 77240 277452 77246
rect 277400 77182 277452 77188
rect 277492 70372 277544 70378
rect 277492 70314 277544 70320
rect 277504 60602 277532 70314
rect 277504 60574 277624 60602
rect 277596 57934 277624 60574
rect 277584 57928 277636 57934
rect 277584 57870 277636 57876
rect 277676 57860 277728 57866
rect 277676 57802 277728 57808
rect 277688 56574 277716 57802
rect 277492 56568 277544 56574
rect 277492 56510 277544 56516
rect 277676 56568 277728 56574
rect 277676 56510 277728 56516
rect 277504 47002 277532 56510
rect 277504 46974 277624 47002
rect 277596 45558 277624 46974
rect 277584 45552 277636 45558
rect 277584 45494 277636 45500
rect 277584 35964 277636 35970
rect 277584 35906 277636 35912
rect 277596 28914 277624 35906
rect 277596 28886 277716 28914
rect 277688 27742 277716 28886
rect 277584 27736 277636 27742
rect 277584 27678 277636 27684
rect 277676 27736 277728 27742
rect 277676 27678 277728 27684
rect 277596 26246 277624 27678
rect 277584 26240 277636 26246
rect 277584 26182 277636 26188
rect 278778 16960 278834 16969
rect 278778 16895 278780 16904
rect 278832 16895 278834 16904
rect 278780 16866 278832 16872
rect 277492 16652 277544 16658
rect 277492 16594 277544 16600
rect 277504 8537 277532 16594
rect 278884 15026 278912 340054
rect 279620 337482 279648 340068
rect 279608 337476 279660 337482
rect 279608 337418 279660 337424
rect 280068 337476 280120 337482
rect 280068 337418 280120 337424
rect 280080 170202 280108 337418
rect 280068 170196 280120 170202
rect 280068 170138 280120 170144
rect 280068 169992 280120 169998
rect 280068 169934 280120 169940
rect 278872 15020 278924 15026
rect 278872 14962 278924 14968
rect 277490 8528 277546 8537
rect 277490 8463 277546 8472
rect 277582 8392 277638 8401
rect 277582 8327 277638 8336
rect 277596 7410 277624 8327
rect 277676 7540 277728 7546
rect 277676 7482 277728 7488
rect 277584 7404 277636 7410
rect 277584 7346 277636 7352
rect 275284 4140 275336 4146
rect 275284 4082 275336 4088
rect 276664 4140 276716 4146
rect 276664 4082 276716 4088
rect 275296 480 275324 4082
rect 276480 3324 276532 3330
rect 276480 3266 276532 3272
rect 276492 480 276520 3266
rect 277688 480 277716 7482
rect 279976 6180 280028 6186
rect 279976 6122 280028 6128
rect 278872 4140 278924 4146
rect 278872 4082 278924 4088
rect 278884 480 278912 4082
rect 279988 2802 280016 6122
rect 280080 4146 280108 169934
rect 280172 10402 280200 340068
rect 280264 340054 280830 340082
rect 280264 15094 280292 340054
rect 281460 337686 281488 340068
rect 281552 340054 282026 340082
rect 282196 340054 282670 340082
rect 281448 337680 281500 337686
rect 281448 337622 281500 337628
rect 280252 15088 280304 15094
rect 280252 15030 280304 15036
rect 281552 10470 281580 340054
rect 282196 331242 282224 340054
rect 283208 337142 283236 340068
rect 283196 337136 283248 337142
rect 283196 337078 283248 337084
rect 283300 335594 283328 340190
rect 284404 340054 284510 340082
rect 283564 337680 283616 337686
rect 283564 337622 283616 337628
rect 281644 331214 282224 331242
rect 283116 335566 283328 335594
rect 281644 321450 281672 331214
rect 281644 321422 281856 321450
rect 281828 309210 281856 321422
rect 283116 318782 283144 335566
rect 283012 318776 283064 318782
rect 283012 318718 283064 318724
rect 283104 318776 283156 318782
rect 283104 318718 283156 318724
rect 283024 317422 283052 318718
rect 283012 317416 283064 317422
rect 283012 317358 283064 317364
rect 283288 317416 283340 317422
rect 283288 317358 283340 317364
rect 281644 309182 281856 309210
rect 281644 302002 281672 309182
rect 281644 301974 281856 302002
rect 281828 299470 281856 301974
rect 281816 299464 281868 299470
rect 281816 299406 281868 299412
rect 283300 292584 283328 317358
rect 283116 292556 283328 292584
rect 281632 289876 281684 289882
rect 281632 289818 281684 289824
rect 281644 289785 281672 289818
rect 281630 289776 281686 289785
rect 281630 289711 281686 289720
rect 281906 289776 281962 289785
rect 281906 289711 281962 289720
rect 281920 280226 281948 289711
rect 281724 280220 281776 280226
rect 281724 280162 281776 280168
rect 281908 280220 281960 280226
rect 281908 280162 281960 280168
rect 281736 280129 281764 280162
rect 283116 280158 283144 292556
rect 283104 280152 283156 280158
rect 281722 280120 281778 280129
rect 283104 280094 283156 280100
rect 281722 280055 281778 280064
rect 281814 279984 281870 279993
rect 281814 279919 281870 279928
rect 281828 263514 281856 279919
rect 283104 270564 283156 270570
rect 283104 270506 283156 270512
rect 281736 263486 281856 263514
rect 281736 260794 281764 263486
rect 283116 260846 283144 270506
rect 283104 260840 283156 260846
rect 281814 260808 281870 260817
rect 281736 260766 281814 260794
rect 281814 260743 281870 260752
rect 281998 260808 282054 260817
rect 283104 260782 283156 260788
rect 281998 260743 282054 260752
rect 282012 259418 282040 260743
rect 282000 259412 282052 259418
rect 282000 259354 282052 259360
rect 283104 251252 283156 251258
rect 283104 251194 283156 251200
rect 281908 241596 281960 241602
rect 281908 241538 281960 241544
rect 281920 241466 281948 241538
rect 283116 241505 283144 251194
rect 282918 241496 282974 241505
rect 281908 241460 281960 241466
rect 282918 241431 282974 241440
rect 283102 241496 283158 241505
rect 283102 241431 283158 241440
rect 281908 241402 281960 241408
rect 281908 234592 281960 234598
rect 281908 234534 281960 234540
rect 281920 222222 281948 234534
rect 282932 231878 282960 241431
rect 282920 231872 282972 231878
rect 282920 231814 282972 231820
rect 283104 231872 283156 231878
rect 283104 231814 283156 231820
rect 281908 222216 281960 222222
rect 281908 222158 281960 222164
rect 281908 220856 281960 220862
rect 281908 220798 281960 220804
rect 281920 215422 281948 220798
rect 281908 215416 281960 215422
rect 283116 215370 283144 231814
rect 281908 215358 281960 215364
rect 283024 215342 283144 215370
rect 281908 215280 281960 215286
rect 281908 215222 281960 215228
rect 283024 215234 283052 215342
rect 281920 211177 281948 215222
rect 283024 215206 283144 215234
rect 281722 211168 281778 211177
rect 281722 211103 281724 211112
rect 281776 211103 281778 211112
rect 281906 211168 281962 211177
rect 281906 211103 281962 211112
rect 281724 211074 281776 211080
rect 281816 202836 281868 202842
rect 281816 202778 281868 202784
rect 281828 201498 281856 202778
rect 281828 201470 281948 201498
rect 281920 196110 281948 201470
rect 281908 196104 281960 196110
rect 283116 196058 283144 215206
rect 281908 196046 281960 196052
rect 283024 196030 283144 196058
rect 281816 195968 281868 195974
rect 281816 195910 281868 195916
rect 283024 195922 283052 196030
rect 281828 186266 281856 195910
rect 283024 195894 283144 195922
rect 281828 186238 281948 186266
rect 281920 183546 281948 186238
rect 283116 183569 283144 195894
rect 281736 183518 281948 183546
rect 282918 183560 282974 183569
rect 281736 167006 281764 183518
rect 282918 183495 282974 183504
rect 283102 183560 283158 183569
rect 283102 183495 283158 183504
rect 282932 173942 282960 183495
rect 282920 173936 282972 173942
rect 282920 173878 282972 173884
rect 283104 173936 283156 173942
rect 283104 173878 283156 173884
rect 281724 167000 281776 167006
rect 281724 166942 281776 166948
rect 281908 167000 281960 167006
rect 281908 166942 281960 166948
rect 281920 157418 281948 166942
rect 283116 164218 283144 173878
rect 283470 169960 283526 169969
rect 283470 169895 283526 169904
rect 283484 169561 283512 169895
rect 283470 169552 283526 169561
rect 283470 169487 283526 169496
rect 283104 164212 283156 164218
rect 283104 164154 283156 164160
rect 281908 157412 281960 157418
rect 281908 157354 281960 157360
rect 281816 157344 281868 157350
rect 281816 157286 281868 157292
rect 281828 143585 281856 157286
rect 283104 154964 283156 154970
rect 283104 154906 283156 154912
rect 281630 143576 281686 143585
rect 281630 143511 281686 143520
rect 281814 143576 281870 143585
rect 281814 143511 281870 143520
rect 281644 135250 281672 143511
rect 283116 138122 283144 154906
rect 283024 138094 283144 138122
rect 283024 137850 283052 138094
rect 283024 137822 283144 137850
rect 281632 135244 281684 135250
rect 281632 135186 281684 135192
rect 281816 129056 281868 129062
rect 281816 128998 281868 129004
rect 281828 106282 281856 128998
rect 283116 125594 283144 137822
rect 283104 125588 283156 125594
rect 283104 125530 283156 125536
rect 283104 116000 283156 116006
rect 283104 115942 283156 115948
rect 283116 106282 283144 115942
rect 281816 106276 281868 106282
rect 281816 106218 281868 106224
rect 281908 106276 281960 106282
rect 281908 106218 281960 106224
rect 283104 106276 283156 106282
rect 283104 106218 283156 106224
rect 281920 96642 281948 106218
rect 281828 96626 281948 96642
rect 283104 96688 283156 96694
rect 283104 96630 283156 96636
rect 281816 96620 281948 96626
rect 281868 96614 281948 96620
rect 282000 96620 282052 96626
rect 281816 96562 281868 96568
rect 282000 96562 282052 96568
rect 281828 96531 281856 96562
rect 282012 77382 282040 96562
rect 281816 77376 281868 77382
rect 281816 77318 281868 77324
rect 282000 77376 282052 77382
rect 282000 77318 282052 77324
rect 281828 72486 281856 77318
rect 281816 72480 281868 72486
rect 281816 72422 281868 72428
rect 282000 72480 282052 72486
rect 282000 72422 282052 72428
rect 282012 67697 282040 72422
rect 281814 67688 281870 67697
rect 281736 67646 281814 67674
rect 281736 66230 281764 67646
rect 281814 67623 281870 67632
rect 281998 67688 282054 67697
rect 281998 67623 282054 67632
rect 281724 66224 281776 66230
rect 281724 66166 281776 66172
rect 283116 60738 283144 96630
rect 283024 60710 283144 60738
rect 283024 60602 283052 60710
rect 283024 60574 283144 60602
rect 281724 56636 281776 56642
rect 281724 56578 281776 56584
rect 281736 48346 281764 56578
rect 283116 56574 283144 60574
rect 283104 56568 283156 56574
rect 283104 56510 283156 56516
rect 281724 48340 281776 48346
rect 281724 48282 281776 48288
rect 281816 48340 281868 48346
rect 281816 48282 281868 48288
rect 281828 38690 281856 48282
rect 282920 47048 282972 47054
rect 282920 46990 282972 46996
rect 282932 46918 282960 46990
rect 282920 46912 282972 46918
rect 282920 46854 282972 46860
rect 283104 46912 283156 46918
rect 283104 46854 283156 46860
rect 283116 45558 283144 46854
rect 283104 45552 283156 45558
rect 283104 45494 283156 45500
rect 281632 38684 281684 38690
rect 281632 38626 281684 38632
rect 281816 38684 281868 38690
rect 281816 38626 281868 38632
rect 281644 31754 281672 38626
rect 281632 31748 281684 31754
rect 281632 31690 281684 31696
rect 281816 31748 281868 31754
rect 281816 31690 281868 31696
rect 281828 22166 281856 31690
rect 282920 27668 282972 27674
rect 282920 27610 282972 27616
rect 281816 22160 281868 22166
rect 281816 22102 281868 22108
rect 281724 22092 281776 22098
rect 281724 22034 281776 22040
rect 281736 16046 281764 22034
rect 282932 19378 282960 27610
rect 282920 19372 282972 19378
rect 282920 19314 282972 19320
rect 283196 19372 283248 19378
rect 283196 19314 283248 19320
rect 281724 16040 281776 16046
rect 281724 15982 281776 15988
rect 283208 10538 283236 19314
rect 283196 10532 283248 10538
rect 283196 10474 283248 10480
rect 281540 10464 281592 10470
rect 281540 10406 281592 10412
rect 280160 10396 280212 10402
rect 280160 10338 280212 10344
rect 283576 8106 283604 337622
rect 283656 337272 283708 337278
rect 283656 337214 283708 337220
rect 283484 8078 283604 8106
rect 281264 7472 281316 7478
rect 281264 7414 281316 7420
rect 280068 4140 280120 4146
rect 280068 4082 280120 4088
rect 279988 2774 280108 2802
rect 280080 480 280108 2774
rect 281276 480 281304 7414
rect 283484 4010 283512 8078
rect 283668 7970 283696 337214
rect 284300 134088 284352 134094
rect 284298 134056 284300 134065
rect 284352 134056 284354 134065
rect 284298 133991 284354 134000
rect 284404 16114 284432 340054
rect 285048 337550 285076 340068
rect 285036 337544 285088 337550
rect 285036 337486 285088 337492
rect 284944 337340 284996 337346
rect 284944 337282 284996 337288
rect 284392 16108 284444 16114
rect 284392 16050 284444 16056
rect 283576 7942 283696 7970
rect 283576 4554 283604 7942
rect 284760 7404 284812 7410
rect 284760 7346 284812 7352
rect 283656 6248 283708 6254
rect 283656 6190 283708 6196
rect 283564 4548 283616 4554
rect 283564 4490 283616 4496
rect 283472 4004 283524 4010
rect 283472 3946 283524 3952
rect 282460 3392 282512 3398
rect 282460 3334 282512 3340
rect 282472 480 282500 3334
rect 283668 480 283696 6190
rect 284772 480 284800 7346
rect 284956 4486 284984 337282
rect 285692 10606 285720 340068
rect 285784 340054 286350 340082
rect 285784 16182 285812 340054
rect 286888 337074 286916 340068
rect 287072 340054 287546 340082
rect 287716 340054 288190 340082
rect 286968 337544 287020 337550
rect 286968 337486 287020 337492
rect 286876 337068 286928 337074
rect 286876 337010 286928 337016
rect 285772 16176 285824 16182
rect 285772 16118 285824 16124
rect 285680 10600 285732 10606
rect 285680 10542 285732 10548
rect 284944 4480 284996 4486
rect 284944 4422 284996 4428
rect 286980 3194 287008 337486
rect 287072 10674 287100 340054
rect 287716 337906 287744 340054
rect 287256 337878 287744 337906
rect 288728 337890 288756 340068
rect 288716 337884 288768 337890
rect 287256 323626 287284 337878
rect 288716 337826 288768 337832
rect 287704 337748 287756 337754
rect 287704 337690 287756 337696
rect 287164 323598 287284 323626
rect 287164 309194 287192 323598
rect 287152 309188 287204 309194
rect 287152 309130 287204 309136
rect 287244 309188 287296 309194
rect 287244 309130 287296 309136
rect 287256 289814 287284 309130
rect 287244 289808 287296 289814
rect 287244 289750 287296 289756
rect 287244 280220 287296 280226
rect 287244 280162 287296 280168
rect 287256 270502 287284 280162
rect 287244 270496 287296 270502
rect 287244 270438 287296 270444
rect 287244 260908 287296 260914
rect 287244 260850 287296 260856
rect 287256 251190 287284 260850
rect 287244 251184 287296 251190
rect 287244 251126 287296 251132
rect 287244 241528 287296 241534
rect 287244 241470 287296 241476
rect 287256 231849 287284 241470
rect 287242 231840 287298 231849
rect 287242 231775 287298 231784
rect 287426 231840 287482 231849
rect 287426 231775 287482 231784
rect 287440 222222 287468 231775
rect 287244 222216 287296 222222
rect 287244 222158 287296 222164
rect 287428 222216 287480 222222
rect 287428 222158 287480 222164
rect 287256 193225 287284 222158
rect 287242 193216 287298 193225
rect 287242 193151 287298 193160
rect 287426 193216 287482 193225
rect 287426 193151 287482 193160
rect 287440 183598 287468 193151
rect 287244 183592 287296 183598
rect 287244 183534 287296 183540
rect 287428 183592 287480 183598
rect 287428 183534 287480 183540
rect 287256 159390 287284 183534
rect 287244 159384 287296 159390
rect 287244 159326 287296 159332
rect 287428 159384 287480 159390
rect 287428 159326 287480 159332
rect 287440 154601 287468 159326
rect 287242 154592 287298 154601
rect 287242 154527 287298 154536
rect 287426 154592 287482 154601
rect 287426 154527 287482 154536
rect 287256 140162 287284 154527
rect 287256 140134 287376 140162
rect 287348 139890 287376 140134
rect 287256 139862 287376 139890
rect 287256 80016 287284 139862
rect 287164 79988 287284 80016
rect 287164 77314 287192 79988
rect 287152 77308 287204 77314
rect 287152 77250 287204 77256
rect 287244 77308 287296 77314
rect 287244 77250 287296 77256
rect 287256 43602 287284 77250
rect 287256 43574 287376 43602
rect 287348 43330 287376 43574
rect 287256 43302 287376 43330
rect 287256 16250 287284 43302
rect 287244 16244 287296 16250
rect 287244 16186 287296 16192
rect 287060 10668 287112 10674
rect 287060 10610 287112 10616
rect 287612 10532 287664 10538
rect 287612 10474 287664 10480
rect 287152 6316 287204 6322
rect 287152 6258 287204 6264
rect 285956 3188 286008 3194
rect 285956 3130 286008 3136
rect 286968 3188 287020 3194
rect 286968 3130 287020 3136
rect 285968 480 285996 3130
rect 287164 480 287192 6258
rect 287624 3534 287652 10474
rect 287716 3738 287744 337690
rect 288820 331242 288848 340190
rect 290016 337618 290044 340068
rect 290004 337612 290056 337618
rect 290004 337554 290056 337560
rect 290568 337006 290596 340068
rect 290556 337000 290608 337006
rect 290556 336942 290608 336948
rect 288544 331214 288848 331242
rect 288544 321314 288572 331214
rect 288544 321286 288664 321314
rect 288636 318782 288664 321286
rect 288624 318776 288676 318782
rect 288624 318718 288676 318724
rect 288624 309188 288676 309194
rect 288624 309130 288676 309136
rect 288636 292534 288664 309130
rect 288624 292528 288676 292534
rect 288624 292470 288676 292476
rect 288624 292392 288676 292398
rect 288624 292334 288676 292340
rect 288636 273222 288664 292334
rect 288624 273216 288676 273222
rect 288624 273158 288676 273164
rect 288624 273080 288676 273086
rect 288624 273022 288676 273028
rect 288636 253910 288664 273022
rect 288624 253904 288676 253910
rect 288624 253846 288676 253852
rect 288624 253768 288676 253774
rect 288624 253710 288676 253716
rect 288636 234598 288664 253710
rect 288624 234592 288676 234598
rect 288624 234534 288676 234540
rect 288624 234456 288676 234462
rect 288624 234398 288676 234404
rect 288636 215370 288664 234398
rect 288544 215342 288664 215370
rect 288544 215234 288572 215342
rect 288544 215206 288664 215234
rect 288636 196058 288664 215206
rect 288544 196030 288664 196058
rect 288544 195922 288572 196030
rect 288544 195894 288664 195922
rect 288636 176662 288664 195894
rect 288624 176656 288676 176662
rect 288624 176598 288676 176604
rect 288624 176520 288676 176526
rect 288624 176462 288676 176468
rect 288636 164218 288664 176462
rect 289636 169992 289688 169998
rect 289634 169960 289636 169969
rect 289688 169960 289690 169969
rect 289634 169895 289690 169904
rect 288624 164212 288676 164218
rect 288624 164154 288676 164160
rect 288624 154964 288676 154970
rect 288624 154906 288676 154912
rect 288636 138122 288664 154906
rect 288544 138094 288664 138122
rect 288544 137850 288572 138094
rect 288544 137822 288664 137850
rect 288636 60738 288664 137822
rect 288544 60710 288664 60738
rect 288544 60602 288572 60710
rect 288544 60574 288664 60602
rect 288636 57934 288664 60574
rect 288624 57928 288676 57934
rect 288624 57870 288676 57876
rect 288532 48340 288584 48346
rect 288532 48282 288584 48288
rect 288544 48226 288572 48282
rect 288544 48198 288664 48226
rect 288636 19378 288664 48198
rect 289818 40216 289874 40225
rect 289818 40151 289874 40160
rect 289832 40089 289860 40151
rect 289818 40080 289874 40089
rect 289818 40015 289874 40024
rect 288440 19372 288492 19378
rect 288440 19314 288492 19320
rect 288624 19372 288676 19378
rect 288624 19314 288676 19320
rect 288348 16924 288400 16930
rect 288348 16866 288400 16872
rect 288360 16697 288388 16866
rect 288346 16688 288402 16697
rect 288346 16623 288402 16632
rect 288452 12594 288480 19314
rect 288360 12566 288480 12594
rect 288360 10742 288388 12566
rect 291212 10810 291240 340068
rect 291304 340054 291870 340082
rect 291304 16318 291332 340054
rect 292408 337822 292436 340068
rect 292592 340054 293066 340082
rect 293236 340054 293710 340082
rect 292396 337816 292448 337822
rect 292396 337758 292448 337764
rect 292488 64864 292540 64870
rect 292488 64806 292540 64812
rect 292500 55321 292528 64806
rect 292486 55312 292542 55321
rect 292486 55247 292542 55256
rect 291292 16312 291344 16318
rect 291292 16254 291344 16260
rect 292592 10878 292620 340054
rect 293236 329050 293264 340054
rect 293868 337612 293920 337618
rect 293868 337554 293920 337560
rect 292764 329044 292816 329050
rect 292764 328986 292816 328992
rect 293224 329044 293276 329050
rect 293224 328986 293276 328992
rect 292776 327078 292804 328986
rect 292764 327072 292816 327078
rect 292764 327014 292816 327020
rect 292764 317484 292816 317490
rect 292764 317426 292816 317432
rect 292776 307766 292804 317426
rect 292764 307760 292816 307766
rect 292764 307702 292816 307708
rect 292764 298240 292816 298246
rect 292764 298182 292816 298188
rect 292776 298110 292804 298182
rect 292764 298104 292816 298110
rect 292764 298046 292816 298052
rect 292672 288448 292724 288454
rect 292672 288390 292724 288396
rect 292684 280226 292712 288390
rect 292672 280220 292724 280226
rect 292672 280162 292724 280168
rect 292764 280220 292816 280226
rect 292764 280162 292816 280168
rect 292776 260914 292804 280162
rect 292764 260908 292816 260914
rect 292764 260850 292816 260856
rect 292764 260772 292816 260778
rect 292764 260714 292816 260720
rect 292776 259434 292804 260714
rect 292776 259406 292896 259434
rect 292868 258058 292896 259406
rect 292856 258052 292908 258058
rect 292856 257994 292908 258000
rect 292856 249756 292908 249762
rect 292856 249698 292908 249704
rect 292868 240174 292896 249698
rect 292764 240168 292816 240174
rect 292764 240110 292816 240116
rect 292856 240168 292908 240174
rect 292856 240110 292908 240116
rect 292776 235498 292804 240110
rect 292776 235470 292896 235498
rect 292868 230586 292896 235470
rect 292764 230580 292816 230586
rect 292764 230522 292816 230528
rect 292856 230580 292908 230586
rect 292856 230522 292908 230528
rect 292776 200122 292804 230522
rect 292764 200116 292816 200122
rect 292764 200058 292816 200064
rect 292856 200116 292908 200122
rect 292856 200058 292908 200064
rect 292868 198694 292896 200058
rect 292856 198688 292908 198694
rect 292856 198630 292908 198636
rect 292764 180872 292816 180878
rect 292764 180814 292816 180820
rect 292776 171290 292804 180814
rect 292764 171284 292816 171290
rect 292764 171226 292816 171232
rect 292764 171148 292816 171154
rect 292764 171090 292816 171096
rect 292776 151774 292804 171090
rect 292946 170096 293002 170105
rect 292946 170031 293002 170040
rect 292960 169998 292988 170031
rect 292948 169992 293000 169998
rect 292948 169934 293000 169940
rect 292764 151768 292816 151774
rect 292764 151710 292816 151716
rect 292764 142180 292816 142186
rect 292764 142122 292816 142128
rect 292776 113150 292804 142122
rect 293774 134328 293830 134337
rect 293774 134263 293830 134272
rect 293788 134094 293816 134263
rect 293776 134088 293828 134094
rect 293776 134030 293828 134036
rect 292764 113144 292816 113150
rect 292764 113086 292816 113092
rect 292764 103624 292816 103630
rect 292764 103566 292816 103572
rect 292776 103494 292804 103566
rect 292764 103488 292816 103494
rect 292764 103430 292816 103436
rect 292672 93900 292724 93906
rect 292672 93842 292724 93848
rect 292684 85354 292712 93842
rect 292684 85326 292804 85354
rect 292776 69086 292804 85326
rect 292764 69080 292816 69086
rect 292764 69022 292816 69028
rect 292764 68944 292816 68950
rect 292764 68886 292816 68892
rect 292776 64870 292804 68886
rect 292764 64864 292816 64870
rect 292764 64806 292816 64812
rect 292762 55312 292818 55321
rect 292762 55247 292818 55256
rect 292776 55214 292804 55247
rect 292764 55208 292816 55214
rect 292764 55150 292816 55156
rect 292948 45620 293000 45626
rect 292948 45562 293000 45568
rect 292960 37194 292988 45562
rect 292948 37188 293000 37194
rect 292948 37130 293000 37136
rect 292764 35964 292816 35970
rect 292764 35906 292816 35912
rect 292776 33810 292804 35906
rect 292776 33782 292988 33810
rect 292960 31634 292988 33782
rect 292868 31606 292988 31634
rect 292868 28966 292896 31606
rect 292764 28960 292816 28966
rect 292764 28902 292816 28908
rect 292856 28960 292908 28966
rect 292856 28902 292908 28908
rect 292776 16386 292804 28902
rect 292764 16380 292816 16386
rect 292764 16322 292816 16328
rect 292580 10872 292632 10878
rect 292580 10814 292632 10820
rect 291200 10804 291252 10810
rect 291200 10746 291252 10752
rect 288348 10736 288400 10742
rect 288348 10678 288400 10684
rect 289820 10668 289872 10674
rect 289820 10610 289872 10616
rect 287704 3732 287756 3738
rect 287704 3674 287756 3680
rect 289832 3670 289860 10610
rect 289912 10600 289964 10606
rect 289912 10542 289964 10548
rect 289820 3664 289872 3670
rect 289820 3606 289872 3612
rect 289544 3596 289596 3602
rect 289544 3538 289596 3544
rect 287612 3528 287664 3534
rect 287612 3470 287664 3476
rect 288348 3256 288400 3262
rect 288348 3198 288400 3204
rect 288360 480 288388 3198
rect 289556 480 289584 3538
rect 289924 3534 289952 10542
rect 292948 10328 293000 10334
rect 292948 10270 293000 10276
rect 290740 6384 290792 6390
rect 290740 6326 290792 6332
rect 289912 3528 289964 3534
rect 289912 3470 289964 3476
rect 290752 480 290780 6326
rect 291936 3664 291988 3670
rect 291936 3606 291988 3612
rect 291948 480 291976 3606
rect 292960 3262 292988 10270
rect 292948 3256 293000 3262
rect 292948 3198 293000 3204
rect 293880 3194 293908 337554
rect 294248 336938 294276 340068
rect 294340 340054 294906 340082
rect 295352 340054 295550 340082
rect 295812 340054 296102 340082
rect 294236 336932 294288 336938
rect 294236 336874 294288 336880
rect 294340 335345 294368 340054
rect 294604 337816 294656 337822
rect 294604 337758 294656 337764
rect 294050 335336 294106 335345
rect 294050 335271 294106 335280
rect 294326 335336 294382 335345
rect 294326 335271 294382 335280
rect 294064 333946 294092 335271
rect 294052 333940 294104 333946
rect 294052 333882 294104 333888
rect 294144 316056 294196 316062
rect 294144 315998 294196 316004
rect 294156 311982 294184 315998
rect 294144 311976 294196 311982
rect 294144 311918 294196 311924
rect 294144 311840 294196 311846
rect 294144 311782 294196 311788
rect 294156 273222 294184 311782
rect 294144 273216 294196 273222
rect 294144 273158 294196 273164
rect 294144 273080 294196 273086
rect 294144 273022 294196 273028
rect 294156 253910 294184 273022
rect 294144 253904 294196 253910
rect 294144 253846 294196 253852
rect 294144 253768 294196 253774
rect 294144 253710 294196 253716
rect 294156 234598 294184 253710
rect 294144 234592 294196 234598
rect 294144 234534 294196 234540
rect 294144 234456 294196 234462
rect 294144 234398 294196 234404
rect 294156 215370 294184 234398
rect 294064 215342 294184 215370
rect 294064 215234 294092 215342
rect 294064 215206 294184 215234
rect 294156 201657 294184 215206
rect 294142 201648 294198 201657
rect 294142 201583 294198 201592
rect 294142 201512 294198 201521
rect 294142 201447 294198 201456
rect 294156 193254 294184 201447
rect 294144 193248 294196 193254
rect 294144 193190 294196 193196
rect 294236 193180 294288 193186
rect 294236 193122 294288 193128
rect 294248 183598 294276 193122
rect 294052 183592 294104 183598
rect 294052 183534 294104 183540
rect 294236 183592 294288 183598
rect 294236 183534 294288 183540
rect 294064 176730 294092 183534
rect 294052 176724 294104 176730
rect 294052 176666 294104 176672
rect 294144 176588 294196 176594
rect 294144 176530 294196 176536
rect 294156 159390 294184 176530
rect 294144 159384 294196 159390
rect 294144 159326 294196 159332
rect 294328 159384 294380 159390
rect 294328 159326 294380 159332
rect 294340 158710 294368 159326
rect 294328 158704 294380 158710
rect 294328 158646 294380 158652
rect 294052 149116 294104 149122
rect 294052 149058 294104 149064
rect 294064 139398 294092 149058
rect 294052 139392 294104 139398
rect 294052 139334 294104 139340
rect 294144 121508 294196 121514
rect 294144 121450 294196 121456
rect 294156 121378 294184 121450
rect 294144 121372 294196 121378
rect 294144 121314 294196 121320
rect 294144 116612 294196 116618
rect 294144 116554 294196 116560
rect 294156 80170 294184 116554
rect 294144 80164 294196 80170
rect 294144 80106 294196 80112
rect 294144 80028 294196 80034
rect 294144 79970 294196 79976
rect 294156 72434 294184 79970
rect 293972 72406 294184 72434
rect 293972 58002 294000 72406
rect 293960 57996 294012 58002
rect 293960 57938 294012 57944
rect 294144 57996 294196 58002
rect 294144 57938 294196 57944
rect 294156 38622 294184 57938
rect 294144 38616 294196 38622
rect 294144 38558 294196 38564
rect 294144 29096 294196 29102
rect 294144 29038 294196 29044
rect 294156 28966 294184 29038
rect 293960 28960 294012 28966
rect 293960 28902 294012 28908
rect 294144 28960 294196 28966
rect 294144 28902 294196 28908
rect 293972 27606 294000 28902
rect 293960 27600 294012 27606
rect 293960 27542 294012 27548
rect 293960 18012 294012 18018
rect 293960 17954 294012 17960
rect 293972 12510 294000 17954
rect 293960 12504 294012 12510
rect 293960 12446 294012 12452
rect 294328 5296 294380 5302
rect 294328 5238 294380 5244
rect 293132 3188 293184 3194
rect 293132 3130 293184 3136
rect 293868 3188 293920 3194
rect 293868 3130 293920 3136
rect 293144 480 293172 3130
rect 294340 480 294368 5238
rect 294616 3398 294644 337758
rect 295246 134328 295302 134337
rect 295246 134263 295302 134272
rect 295260 133929 295288 134263
rect 295246 133920 295302 133929
rect 295246 133855 295302 133864
rect 295352 11830 295380 340054
rect 295812 338094 295840 340054
rect 295800 338088 295852 338094
rect 295800 338030 295852 338036
rect 295616 328500 295668 328506
rect 295616 328442 295668 328448
rect 295628 311930 295656 328442
rect 295536 311902 295656 311930
rect 295536 303090 295564 311902
rect 295536 303062 295748 303090
rect 295720 298110 295748 303062
rect 295708 298104 295760 298110
rect 295708 298046 295760 298052
rect 295708 293276 295760 293282
rect 295708 293218 295760 293224
rect 295720 280158 295748 293218
rect 295432 280152 295484 280158
rect 295432 280094 295484 280100
rect 295708 280152 295760 280158
rect 295708 280094 295760 280100
rect 295444 278730 295472 280094
rect 295432 278724 295484 278730
rect 295432 278666 295484 278672
rect 295616 269136 295668 269142
rect 295616 269078 295668 269084
rect 295628 260846 295656 269078
rect 295432 260840 295484 260846
rect 295432 260782 295484 260788
rect 295616 260840 295668 260846
rect 295616 260782 295668 260788
rect 295444 259418 295472 260782
rect 295432 259412 295484 259418
rect 295432 259354 295484 259360
rect 295524 240100 295576 240106
rect 295524 240042 295576 240048
rect 295536 237386 295564 240042
rect 295524 237380 295576 237386
rect 295524 237322 295576 237328
rect 295524 227792 295576 227798
rect 295524 227734 295576 227740
rect 295536 225010 295564 227734
rect 295524 225004 295576 225010
rect 295524 224946 295576 224952
rect 295616 224868 295668 224874
rect 295616 224810 295668 224816
rect 295628 215422 295656 224810
rect 295616 215416 295668 215422
rect 295616 215358 295668 215364
rect 295432 211132 295484 211138
rect 295432 211074 295484 211080
rect 295444 206310 295472 211074
rect 295432 206304 295484 206310
rect 295432 206246 295484 206252
rect 295708 206304 295760 206310
rect 295708 206246 295760 206252
rect 295720 200122 295748 206246
rect 295432 200116 295484 200122
rect 295432 200058 295484 200064
rect 295708 200116 295760 200122
rect 295708 200058 295760 200064
rect 295444 190505 295472 200058
rect 295430 190496 295486 190505
rect 295430 190431 295486 190440
rect 295614 190496 295670 190505
rect 295614 190431 295670 190440
rect 295628 188494 295656 190431
rect 295616 188488 295668 188494
rect 295616 188430 295668 188436
rect 295616 183592 295668 183598
rect 295616 183534 295668 183540
rect 295628 175930 295656 183534
rect 295536 175902 295656 175930
rect 295536 171086 295564 175902
rect 295524 171080 295576 171086
rect 295524 171022 295576 171028
rect 295524 161492 295576 161498
rect 295524 161434 295576 161440
rect 295536 155394 295564 161434
rect 295536 155366 295656 155394
rect 295628 151842 295656 155366
rect 295616 151836 295668 151842
rect 295616 151778 295668 151784
rect 295708 151700 295760 151706
rect 295708 151642 295760 151648
rect 295720 150414 295748 151642
rect 295708 150408 295760 150414
rect 295708 150350 295760 150356
rect 295616 140820 295668 140826
rect 295616 140762 295668 140768
rect 295628 140706 295656 140762
rect 295628 140678 295748 140706
rect 295720 131345 295748 140678
rect 295706 131336 295762 131345
rect 295706 131271 295762 131280
rect 295522 131200 295578 131209
rect 295522 131135 295578 131144
rect 295536 131102 295564 131135
rect 295524 131096 295576 131102
rect 295524 131038 295576 131044
rect 295616 121508 295668 121514
rect 295616 121450 295668 121456
rect 295628 118794 295656 121450
rect 295616 118788 295668 118794
rect 295616 118730 295668 118736
rect 295616 118652 295668 118658
rect 295616 118594 295668 118600
rect 295628 111790 295656 118594
rect 295616 111784 295668 111790
rect 295616 111726 295668 111732
rect 295708 102196 295760 102202
rect 295708 102138 295760 102144
rect 295720 80170 295748 102138
rect 295524 80164 295576 80170
rect 295524 80106 295576 80112
rect 295708 80164 295760 80170
rect 295708 80106 295760 80112
rect 295536 66586 295564 80106
rect 295536 66558 295656 66586
rect 295628 66314 295656 66558
rect 295536 66286 295656 66314
rect 295536 58002 295564 66286
rect 295524 57996 295576 58002
rect 295524 57938 295576 57944
rect 295616 57860 295668 57866
rect 295616 57802 295668 57808
rect 295628 48278 295656 57802
rect 295616 48272 295668 48278
rect 295616 48214 295668 48220
rect 295708 48272 295760 48278
rect 295708 48214 295760 48220
rect 295720 38350 295748 48214
rect 295708 38344 295760 38350
rect 295708 38286 295760 38292
rect 295708 38208 295760 38214
rect 295708 38150 295760 38156
rect 295720 29050 295748 38150
rect 295628 29022 295748 29050
rect 295628 28966 295656 29022
rect 295524 28960 295576 28966
rect 295524 28902 295576 28908
rect 295616 28960 295668 28966
rect 295616 28902 295668 28908
rect 295536 15162 295564 28902
rect 295524 15156 295576 15162
rect 295524 15098 295576 15104
rect 295340 11824 295392 11830
rect 295340 11766 295392 11772
rect 296732 5370 296760 340068
rect 296916 340054 297390 340082
rect 297560 340054 297942 340082
rect 298112 340054 298586 340082
rect 298664 340054 299230 340082
rect 299584 340054 299782 340082
rect 300136 340054 300426 340082
rect 300872 340054 300978 340082
rect 301056 340054 301622 340082
rect 302266 340054 302464 340082
rect 296812 335640 296864 335646
rect 296812 335582 296864 335588
rect 296824 8974 296852 335582
rect 296916 13190 296944 340054
rect 297560 335646 297588 340054
rect 297548 335640 297600 335646
rect 297548 335582 297600 335588
rect 296904 13184 296956 13190
rect 296904 13126 296956 13132
rect 296812 8968 296864 8974
rect 296812 8910 296864 8916
rect 298112 5438 298140 340054
rect 298664 335628 298692 340054
rect 298388 335600 298692 335628
rect 299480 335640 299532 335646
rect 298388 311930 298416 335600
rect 299480 335582 299532 335588
rect 298296 311902 298416 311930
rect 298296 302326 298324 311902
rect 298284 302320 298336 302326
rect 298284 302262 298336 302268
rect 298376 302116 298428 302122
rect 298376 302058 298428 302064
rect 298388 296682 298416 302058
rect 298376 296676 298428 296682
rect 298376 296618 298428 296624
rect 298468 287088 298520 287094
rect 298468 287030 298520 287036
rect 298480 280158 298508 287030
rect 298468 280152 298520 280158
rect 298468 280094 298520 280100
rect 298284 280084 298336 280090
rect 298284 280026 298336 280032
rect 298296 278769 298324 280026
rect 298282 278760 298338 278769
rect 298282 278695 298338 278704
rect 298558 278760 298614 278769
rect 298558 278695 298614 278704
rect 298572 253722 298600 278695
rect 298296 253694 298600 253722
rect 298296 251190 298324 253694
rect 298284 251184 298336 251190
rect 298284 251126 298336 251132
rect 298192 242684 298244 242690
rect 298192 242626 298244 242632
rect 298204 240106 298232 242626
rect 298192 240100 298244 240106
rect 298192 240042 298244 240048
rect 298284 240100 298336 240106
rect 298284 240042 298336 240048
rect 298296 238746 298324 240042
rect 298284 238740 298336 238746
rect 298284 238682 298336 238688
rect 298560 238740 298612 238746
rect 298560 238682 298612 238688
rect 298572 220862 298600 238682
rect 298376 220856 298428 220862
rect 298376 220798 298428 220804
rect 298560 220856 298612 220862
rect 298560 220798 298612 220804
rect 298388 215490 298416 220798
rect 298376 215484 298428 215490
rect 298376 215426 298428 215432
rect 298284 211268 298336 211274
rect 298284 211210 298336 211216
rect 298296 211138 298324 211210
rect 298284 211132 298336 211138
rect 298284 211074 298336 211080
rect 298284 205624 298336 205630
rect 298284 205566 298336 205572
rect 298296 201498 298324 205566
rect 298296 201470 298416 201498
rect 298388 193254 298416 201470
rect 298376 193248 298428 193254
rect 298376 193190 298428 193196
rect 298284 191888 298336 191894
rect 298284 191830 298336 191836
rect 298296 186522 298324 191830
rect 298284 186516 298336 186522
rect 298284 186458 298336 186464
rect 298376 183592 298428 183598
rect 298376 183534 298428 183540
rect 298388 176798 298416 183534
rect 298376 176792 298428 176798
rect 298376 176734 298428 176740
rect 298284 176656 298336 176662
rect 298284 176598 298336 176604
rect 298296 172514 298324 176598
rect 298284 172508 298336 172514
rect 298284 172450 298336 172456
rect 298190 170096 298246 170105
rect 298190 170031 298246 170040
rect 298204 169969 298232 170031
rect 298190 169960 298246 169969
rect 298190 169895 298246 169904
rect 298284 167000 298336 167006
rect 298284 166942 298336 166948
rect 298296 162874 298324 166942
rect 298296 162846 298416 162874
rect 298388 133822 298416 162846
rect 298376 133816 298428 133822
rect 298376 133758 298428 133764
rect 298376 124228 298428 124234
rect 298376 124170 298428 124176
rect 298388 119406 298416 124170
rect 298376 119400 298428 119406
rect 298376 119342 298428 119348
rect 298192 114572 298244 114578
rect 298192 114514 298244 114520
rect 298204 114442 298232 114514
rect 298192 114436 298244 114442
rect 298192 114378 298244 114384
rect 298376 104916 298428 104922
rect 298376 104858 298428 104864
rect 298388 99482 298416 104858
rect 298376 99476 298428 99482
rect 298376 99418 298428 99424
rect 298376 95260 298428 95266
rect 298376 95202 298428 95208
rect 298388 89758 298416 95202
rect 298376 89752 298428 89758
rect 298376 89694 298428 89700
rect 298376 85604 298428 85610
rect 298376 85546 298428 85552
rect 298388 80782 298416 85546
rect 298376 80776 298428 80782
rect 298376 80718 298428 80724
rect 298376 67652 298428 67658
rect 298376 67594 298428 67600
rect 298388 57916 298416 67594
rect 298296 57888 298416 57916
rect 298296 56574 298324 57888
rect 298284 56568 298336 56574
rect 298284 56510 298336 56516
rect 298376 46980 298428 46986
rect 298376 46922 298428 46928
rect 298388 42090 298416 46922
rect 298376 42084 298428 42090
rect 298376 42026 298428 42032
rect 298192 32428 298244 32434
rect 298192 32370 298244 32376
rect 298204 19394 298232 32370
rect 298204 19366 298324 19394
rect 298296 14498 298324 19366
rect 299294 16688 299350 16697
rect 299294 16623 299350 16632
rect 299308 16561 299336 16623
rect 299294 16552 299350 16561
rect 299294 16487 299350 16496
rect 298204 14470 298324 14498
rect 298204 9602 298232 14470
rect 298204 9574 298324 9602
rect 298296 7585 298324 9574
rect 298282 7576 298338 7585
rect 298282 7511 298338 7520
rect 299492 5506 299520 335582
rect 299584 8945 299612 340054
rect 300136 335646 300164 340054
rect 300124 335640 300176 335646
rect 300124 335582 300176 335588
rect 299664 10464 299716 10470
rect 299664 10406 299716 10412
rect 299570 8936 299626 8945
rect 299570 8871 299626 8880
rect 299480 5500 299532 5506
rect 299480 5442 299532 5448
rect 298100 5432 298152 5438
rect 298100 5374 298152 5380
rect 296720 5364 296772 5370
rect 296720 5306 296772 5312
rect 297916 5364 297968 5370
rect 297916 5306 297968 5312
rect 296720 3596 296772 3602
rect 296720 3538 296772 3544
rect 294604 3392 294656 3398
rect 294604 3334 294656 3340
rect 295524 3392 295576 3398
rect 295524 3334 295576 3340
rect 295536 480 295564 3334
rect 296732 480 296760 3538
rect 297928 480 297956 5306
rect 299112 3732 299164 3738
rect 299112 3674 299164 3680
rect 299124 480 299152 3674
rect 299676 3670 299704 10406
rect 300872 7342 300900 340054
rect 301056 10946 301084 340054
rect 302332 335640 302384 335646
rect 302332 335582 302384 335588
rect 302146 40080 302202 40089
rect 302146 40015 302148 40024
rect 302200 40015 302202 40024
rect 302148 39986 302200 39992
rect 302344 11014 302372 335582
rect 302436 11966 302464 340054
rect 302528 340054 302818 340082
rect 303080 340054 303462 340082
rect 303724 340054 304106 340082
rect 304368 340054 304658 340082
rect 305012 340054 305302 340082
rect 305380 340054 305946 340082
rect 302424 11960 302476 11966
rect 302424 11902 302476 11908
rect 302332 11008 302384 11014
rect 302332 10950 302384 10956
rect 301044 10940 301096 10946
rect 301044 10882 301096 10888
rect 300952 10396 301004 10402
rect 300952 10338 301004 10344
rect 300860 7336 300912 7342
rect 300860 7278 300912 7284
rect 300308 4004 300360 4010
rect 300308 3946 300360 3952
rect 299664 3664 299716 3670
rect 299664 3606 299716 3612
rect 300320 480 300348 3946
rect 300964 3738 300992 10338
rect 302528 7274 302556 340054
rect 303080 335646 303108 340054
rect 303068 335640 303120 335646
rect 303068 335582 303120 335588
rect 303620 335640 303672 335646
rect 303620 335582 303672 335588
rect 303632 13326 303660 335582
rect 303620 13320 303672 13326
rect 303620 13262 303672 13268
rect 303724 13258 303752 340054
rect 304368 335646 304396 340054
rect 304356 335640 304408 335646
rect 304356 335582 304408 335588
rect 303712 13252 303764 13258
rect 303712 13194 303764 13200
rect 305012 10266 305040 340054
rect 305380 335594 305408 340054
rect 305196 335566 305408 335594
rect 306380 335640 306432 335646
rect 306380 335582 306432 335588
rect 305196 331226 305224 335566
rect 305184 331220 305236 331226
rect 305184 331162 305236 331168
rect 305276 331152 305328 331158
rect 305276 331094 305328 331100
rect 305288 309194 305316 331094
rect 305184 309188 305236 309194
rect 305184 309130 305236 309136
rect 305276 309188 305328 309194
rect 305276 309130 305328 309136
rect 305196 299470 305224 309130
rect 305184 299464 305236 299470
rect 305184 299406 305236 299412
rect 305184 289876 305236 289882
rect 305184 289818 305236 289824
rect 305196 280158 305224 289818
rect 305184 280152 305236 280158
rect 305184 280094 305236 280100
rect 305184 270564 305236 270570
rect 305184 270506 305236 270512
rect 305196 260846 305224 270506
rect 305184 260840 305236 260846
rect 305184 260782 305236 260788
rect 305184 251252 305236 251258
rect 305184 251194 305236 251200
rect 305196 241505 305224 251194
rect 305182 241496 305238 241505
rect 305182 241431 305238 241440
rect 305366 241496 305422 241505
rect 305366 241431 305422 241440
rect 305380 231878 305408 241431
rect 305184 231872 305236 231878
rect 305184 231814 305236 231820
rect 305368 231872 305420 231878
rect 305368 231814 305420 231820
rect 305196 222193 305224 231814
rect 305182 222184 305238 222193
rect 305182 222119 305238 222128
rect 305366 222184 305422 222193
rect 305366 222119 305422 222128
rect 305380 212566 305408 222119
rect 305184 212560 305236 212566
rect 305184 212502 305236 212508
rect 305368 212560 305420 212566
rect 305368 212502 305420 212508
rect 305196 202881 305224 212502
rect 305182 202872 305238 202881
rect 305182 202807 305238 202816
rect 305366 202872 305422 202881
rect 305366 202807 305422 202816
rect 305380 193254 305408 202807
rect 305184 193248 305236 193254
rect 305184 193190 305236 193196
rect 305368 193248 305420 193254
rect 305368 193190 305420 193196
rect 305196 183569 305224 193190
rect 305182 183560 305238 183569
rect 305182 183495 305238 183504
rect 305366 183560 305422 183569
rect 305366 183495 305422 183504
rect 305380 173942 305408 183495
rect 305184 173936 305236 173942
rect 305184 173878 305236 173884
rect 305368 173936 305420 173942
rect 305368 173878 305420 173884
rect 305196 164218 305224 173878
rect 305184 164212 305236 164218
rect 305184 164154 305236 164160
rect 305276 164212 305328 164218
rect 305276 164154 305328 164160
rect 305288 120766 305316 164154
rect 305276 120760 305328 120766
rect 305276 120702 305328 120708
rect 305184 116000 305236 116006
rect 305184 115942 305236 115948
rect 305196 106282 305224 115942
rect 305184 106276 305236 106282
rect 305184 106218 305236 106224
rect 305184 96688 305236 96694
rect 305184 96630 305236 96636
rect 305196 86970 305224 96630
rect 305184 86964 305236 86970
rect 305184 86906 305236 86912
rect 305184 77308 305236 77314
rect 305184 77250 305236 77256
rect 305196 67590 305224 77250
rect 305184 67584 305236 67590
rect 305184 67526 305236 67532
rect 305276 67584 305328 67590
rect 305276 67526 305328 67532
rect 305288 22234 305316 67526
rect 305276 22228 305328 22234
rect 305276 22170 305328 22176
rect 305092 19372 305144 19378
rect 305092 19314 305144 19320
rect 305104 13530 305132 19314
rect 305092 13524 305144 13530
rect 305092 13466 305144 13472
rect 305000 10260 305052 10266
rect 305000 10202 305052 10208
rect 306392 10198 306420 335582
rect 306484 13462 306512 340068
rect 306760 340054 307142 340082
rect 307786 340054 307984 340082
rect 306760 335646 306788 340054
rect 306748 335640 306800 335646
rect 306748 335582 306800 335588
rect 307852 335640 307904 335646
rect 307852 335582 307904 335588
rect 307298 40216 307354 40225
rect 307298 40151 307354 40160
rect 307312 40050 307340 40151
rect 307300 40044 307352 40050
rect 307300 39986 307352 39992
rect 307864 13598 307892 335582
rect 307852 13592 307904 13598
rect 307852 13534 307904 13540
rect 306472 13456 306524 13462
rect 306472 13398 306524 13404
rect 307956 13394 307984 340054
rect 308048 340054 308338 340082
rect 308508 340054 308982 340082
rect 309152 340054 309626 340082
rect 309704 340054 310178 340082
rect 310532 340054 310822 340082
rect 311176 340054 311466 340082
rect 308048 335646 308076 340054
rect 308036 335640 308088 335646
rect 308036 335582 308088 335588
rect 308508 331242 308536 340054
rect 308048 331214 308536 331242
rect 308048 183569 308076 331214
rect 308034 183560 308090 183569
rect 308034 183495 308090 183504
rect 308310 183560 308366 183569
rect 308310 183495 308366 183504
rect 308324 173942 308352 183495
rect 308128 173936 308180 173942
rect 308128 173878 308180 173884
rect 308312 173936 308364 173942
rect 308312 173878 308364 173884
rect 308140 164218 308168 173878
rect 308128 164212 308180 164218
rect 308128 164154 308180 164160
rect 308312 164212 308364 164218
rect 308312 164154 308364 164160
rect 308324 154601 308352 164154
rect 308034 154592 308090 154601
rect 308034 154527 308090 154536
rect 308310 154592 308366 154601
rect 308310 154527 308366 154536
rect 308048 147642 308076 154527
rect 308048 147614 308168 147642
rect 308140 144906 308168 147614
rect 308128 144900 308180 144906
rect 308128 144842 308180 144848
rect 308312 144900 308364 144906
rect 308312 144842 308364 144848
rect 308324 135289 308352 144842
rect 308126 135280 308182 135289
rect 308126 135215 308182 135224
rect 308310 135280 308366 135289
rect 308310 135215 308366 135224
rect 308140 125594 308168 135215
rect 308128 125588 308180 125594
rect 308128 125530 308180 125536
rect 308312 125588 308364 125594
rect 308312 125530 308364 125536
rect 308324 115977 308352 125530
rect 308034 115968 308090 115977
rect 308034 115903 308090 115912
rect 308310 115968 308366 115977
rect 308310 115903 308366 115912
rect 308048 106282 308076 115903
rect 308036 106276 308088 106282
rect 308036 106218 308088 106224
rect 308220 106276 308272 106282
rect 308220 106218 308272 106224
rect 308232 96665 308260 106218
rect 308034 96656 308090 96665
rect 308034 96591 308090 96600
rect 308218 96656 308274 96665
rect 308218 96591 308274 96600
rect 308048 86970 308076 96591
rect 308036 86964 308088 86970
rect 308036 86906 308088 86912
rect 308036 77308 308088 77314
rect 308036 77250 308088 77256
rect 308048 67590 308076 77250
rect 308036 67584 308088 67590
rect 308036 67526 308088 67532
rect 308036 57996 308088 58002
rect 308036 57938 308088 57944
rect 308048 50946 308076 57938
rect 308048 50918 308168 50946
rect 308140 48278 308168 50918
rect 308128 48272 308180 48278
rect 308128 48214 308180 48220
rect 308128 38684 308180 38690
rect 308128 38626 308180 38632
rect 308140 28966 308168 38626
rect 308128 28960 308180 28966
rect 308128 28902 308180 28908
rect 308036 19372 308088 19378
rect 308036 19314 308088 19320
rect 307944 13388 307996 13394
rect 307944 13330 307996 13336
rect 308048 12594 308076 19314
rect 309046 16824 309102 16833
rect 309046 16759 309102 16768
rect 309060 16425 309088 16759
rect 309046 16416 309102 16425
rect 309046 16351 309102 16360
rect 309152 13666 309180 340054
rect 309704 331294 309732 340054
rect 309784 337952 309836 337958
rect 309784 337894 309836 337900
rect 309692 331288 309744 331294
rect 309692 331230 309744 331236
rect 309416 328500 309468 328506
rect 309416 328442 309468 328448
rect 309428 311930 309456 328442
rect 309336 311902 309456 311930
rect 309336 309126 309364 311902
rect 309324 309120 309376 309126
rect 309324 309062 309376 309068
rect 309416 299532 309468 299538
rect 309416 299474 309468 299480
rect 309428 299441 309456 299474
rect 309414 299432 309470 299441
rect 309414 299367 309470 299376
rect 309598 299432 309654 299441
rect 309598 299367 309654 299376
rect 309612 289882 309640 299367
rect 309324 289876 309376 289882
rect 309324 289818 309376 289824
rect 309600 289876 309652 289882
rect 309600 289818 309652 289824
rect 309336 289746 309364 289818
rect 309324 289740 309376 289746
rect 309324 289682 309376 289688
rect 309416 280220 309468 280226
rect 309416 280162 309468 280168
rect 309428 280129 309456 280162
rect 309414 280120 309470 280129
rect 309414 280055 309470 280064
rect 309598 280120 309654 280129
rect 309598 280055 309654 280064
rect 309612 270570 309640 280055
rect 309324 270564 309376 270570
rect 309324 270506 309376 270512
rect 309600 270564 309652 270570
rect 309600 270506 309652 270512
rect 309336 270434 309364 270506
rect 309324 270428 309376 270434
rect 309324 270370 309376 270376
rect 309416 260908 309468 260914
rect 309416 260850 309468 260856
rect 309428 260778 309456 260850
rect 309416 260772 309468 260778
rect 309416 260714 309468 260720
rect 309324 251252 309376 251258
rect 309324 251194 309376 251200
rect 309336 251161 309364 251194
rect 309322 251152 309378 251161
rect 309322 251087 309378 251096
rect 309506 251152 309562 251161
rect 309506 251087 309562 251096
rect 309520 241534 309548 251087
rect 309508 241528 309560 241534
rect 309508 241470 309560 241476
rect 309600 241528 309652 241534
rect 309600 241470 309652 241476
rect 309612 231962 309640 241470
rect 309336 231934 309640 231962
rect 309336 225010 309364 231934
rect 309324 225004 309376 225010
rect 309324 224946 309376 224952
rect 309416 224868 309468 224874
rect 309416 224810 309468 224816
rect 309428 222170 309456 224810
rect 309336 222142 309456 222170
rect 309336 215354 309364 222142
rect 309324 215348 309376 215354
rect 309324 215290 309376 215296
rect 309416 212560 309468 212566
rect 309416 212502 309468 212508
rect 309428 205698 309456 212502
rect 309416 205692 309468 205698
rect 309416 205634 309468 205640
rect 309428 202910 309456 202941
rect 309416 202904 309468 202910
rect 309336 202852 309416 202858
rect 309336 202846 309468 202852
rect 309336 202830 309456 202846
rect 309336 196042 309364 202830
rect 309324 196036 309376 196042
rect 309324 195978 309376 195984
rect 309416 193248 309468 193254
rect 309416 193190 309468 193196
rect 309428 186402 309456 193190
rect 309244 186374 309456 186402
rect 309244 183841 309272 186374
rect 309230 183832 309286 183841
rect 309230 183767 309286 183776
rect 309414 183696 309470 183705
rect 309414 183631 309470 183640
rect 309428 176798 309456 183631
rect 309416 176792 309468 176798
rect 309416 176734 309468 176740
rect 309324 176656 309376 176662
rect 309324 176598 309376 176604
rect 309336 172514 309364 176598
rect 309324 172508 309376 172514
rect 309324 172450 309376 172456
rect 309324 164212 309376 164218
rect 309324 164154 309376 164160
rect 309336 162874 309364 164154
rect 309336 162846 309456 162874
rect 309428 153218 309456 162846
rect 309336 153202 309456 153218
rect 309324 153196 309456 153202
rect 309376 153190 309456 153196
rect 309508 153196 309560 153202
rect 309324 153138 309376 153144
rect 309508 153138 309560 153144
rect 309336 153107 309364 153138
rect 309520 143562 309548 153138
rect 309520 143534 309640 143562
rect 309612 135318 309640 143534
rect 309324 135312 309376 135318
rect 309324 135254 309376 135260
rect 309600 135312 309652 135318
rect 309600 135254 309652 135260
rect 309336 132462 309364 135254
rect 309324 132456 309376 132462
rect 309324 132398 309376 132404
rect 309508 122868 309560 122874
rect 309508 122810 309560 122816
rect 309520 113218 309548 122810
rect 309324 113212 309376 113218
rect 309324 113154 309376 113160
rect 309508 113212 309560 113218
rect 309508 113154 309560 113160
rect 309336 101402 309364 113154
rect 309244 101374 309364 101402
rect 309244 99362 309272 101374
rect 309244 99334 309364 99362
rect 309336 86970 309364 99334
rect 309324 86964 309376 86970
rect 309324 86906 309376 86912
rect 309324 77308 309376 77314
rect 309324 77250 309376 77256
rect 309336 67674 309364 77250
rect 309336 67646 309456 67674
rect 309428 66230 309456 67646
rect 309416 66224 309468 66230
rect 309416 66166 309468 66172
rect 309416 48408 309468 48414
rect 309416 48350 309468 48356
rect 309428 42090 309456 48350
rect 309416 42084 309468 42090
rect 309416 42026 309468 42032
rect 309324 29028 309376 29034
rect 309324 28970 309376 28976
rect 309336 19258 309364 28970
rect 309336 19230 309456 19258
rect 309428 14346 309456 19230
rect 309416 14340 309468 14346
rect 309416 14282 309468 14288
rect 309140 13660 309192 13666
rect 309140 13602 309192 13608
rect 307864 12566 308076 12594
rect 306380 10192 306432 10198
rect 306380 10134 306432 10140
rect 307864 10130 307892 12566
rect 307852 10124 307904 10130
rect 307852 10066 307904 10072
rect 302516 7268 302568 7274
rect 302516 7210 302568 7216
rect 308588 6520 308640 6526
rect 308588 6462 308640 6468
rect 305000 6452 305052 6458
rect 305000 6394 305052 6400
rect 301412 5432 301464 5438
rect 301412 5374 301464 5380
rect 300952 3732 301004 3738
rect 300952 3674 301004 3680
rect 301424 480 301452 5374
rect 303804 3664 303856 3670
rect 303804 3606 303856 3612
rect 302608 3256 302660 3262
rect 302608 3198 302660 3204
rect 302620 480 302648 3198
rect 303816 480 303844 3606
rect 305012 480 305040 6394
rect 307392 3732 307444 3738
rect 307392 3674 307444 3680
rect 306196 3324 306248 3330
rect 306196 3266 306248 3272
rect 306208 480 306236 3266
rect 307404 480 307432 3674
rect 308600 480 308628 6462
rect 309796 3738 309824 337894
rect 310426 28928 310482 28937
rect 310426 28863 310482 28872
rect 310440 19378 310468 28863
rect 310428 19372 310480 19378
rect 310428 19314 310480 19320
rect 310532 10062 310560 340054
rect 311176 335646 311204 340054
rect 311900 337884 311952 337890
rect 311900 337826 311952 337832
rect 310704 335640 310756 335646
rect 310704 335582 310756 335588
rect 311164 335640 311216 335646
rect 311164 335582 311216 335588
rect 310716 311930 310744 335582
rect 310624 311902 310744 311930
rect 310624 311794 310652 311902
rect 310624 311766 310744 311794
rect 310716 299470 310744 311766
rect 310704 299464 310756 299470
rect 310704 299406 310756 299412
rect 310704 289876 310756 289882
rect 310704 289818 310756 289824
rect 310716 280158 310744 289818
rect 310704 280152 310756 280158
rect 310704 280094 310756 280100
rect 310704 270564 310756 270570
rect 310704 270506 310756 270512
rect 310716 260846 310744 270506
rect 310704 260840 310756 260846
rect 310704 260782 310756 260788
rect 310704 251252 310756 251258
rect 310704 251194 310756 251200
rect 310716 241505 310744 251194
rect 310702 241496 310758 241505
rect 310702 241431 310758 241440
rect 310886 241496 310942 241505
rect 310886 241431 310942 241440
rect 310900 231878 310928 241431
rect 310704 231872 310756 231878
rect 310704 231814 310756 231820
rect 310888 231872 310940 231878
rect 310888 231814 310940 231820
rect 310716 222193 310744 231814
rect 310702 222184 310758 222193
rect 310702 222119 310758 222128
rect 310886 222184 310942 222193
rect 310886 222119 310942 222128
rect 310900 212566 310928 222119
rect 310704 212560 310756 212566
rect 310704 212502 310756 212508
rect 310888 212560 310940 212566
rect 310888 212502 310940 212508
rect 310716 202881 310744 212502
rect 310702 202872 310758 202881
rect 310702 202807 310758 202816
rect 310886 202872 310942 202881
rect 310886 202807 310942 202816
rect 310900 193254 310928 202807
rect 310704 193248 310756 193254
rect 310704 193190 310756 193196
rect 310888 193248 310940 193254
rect 310888 193190 310940 193196
rect 310716 176746 310744 193190
rect 310624 176718 310744 176746
rect 310624 176610 310652 176718
rect 310624 176582 310744 176610
rect 310716 164218 310744 176582
rect 310704 164212 310756 164218
rect 310704 164154 310756 164160
rect 310888 164212 310940 164218
rect 310888 164154 310940 164160
rect 310900 154601 310928 164154
rect 310702 154592 310758 154601
rect 310702 154527 310758 154536
rect 310886 154592 310942 154601
rect 310886 154527 310942 154536
rect 310716 144906 310744 154527
rect 310704 144900 310756 144906
rect 310704 144842 310756 144848
rect 310888 144900 310940 144906
rect 310888 144842 310940 144848
rect 310900 135289 310928 144842
rect 310702 135280 310758 135289
rect 310702 135215 310758 135224
rect 310886 135280 310942 135289
rect 310886 135215 310942 135224
rect 310716 125594 310744 135215
rect 310704 125588 310756 125594
rect 310704 125530 310756 125536
rect 310704 116000 310756 116006
rect 310704 115942 310756 115948
rect 310716 106282 310744 115942
rect 310704 106276 310756 106282
rect 310704 106218 310756 106224
rect 310704 96688 310756 96694
rect 310704 96630 310756 96636
rect 310716 86970 310744 96630
rect 310704 86964 310756 86970
rect 310704 86906 310756 86912
rect 310704 77308 310756 77314
rect 310704 77250 310756 77256
rect 310716 60636 310744 77250
rect 310624 60608 310744 60636
rect 310624 60466 310652 60608
rect 310624 60438 310744 60466
rect 310716 48521 310744 60438
rect 310702 48512 310758 48521
rect 310702 48447 310758 48456
rect 310610 48376 310666 48385
rect 310610 48311 310666 48320
rect 310624 46918 310652 48311
rect 310612 46912 310664 46918
rect 310612 46854 310664 46860
rect 310612 41404 310664 41410
rect 310612 41346 310664 41352
rect 310624 28937 310652 41346
rect 310610 28928 310666 28937
rect 310610 28863 310666 28872
rect 310704 19372 310756 19378
rect 310704 19314 310756 19320
rect 310716 13734 310744 19314
rect 310704 13728 310756 13734
rect 310704 13670 310756 13676
rect 310520 10056 310572 10062
rect 310520 9998 310572 10004
rect 311912 9994 311940 337826
rect 312004 14414 312032 340068
rect 312280 340054 312662 340082
rect 313306 340054 313412 340082
rect 312280 337890 312308 340054
rect 312268 337884 312320 337890
rect 312268 337826 312320 337832
rect 311992 14408 312044 14414
rect 311992 14350 312044 14356
rect 313384 12034 313412 340054
rect 313568 340054 313858 340082
rect 314120 340054 314502 340082
rect 314764 340054 315146 340082
rect 315408 340054 315698 340082
rect 316144 340054 316342 340082
rect 316696 340054 316986 340082
rect 317432 340054 317538 340082
rect 317708 340054 318182 340082
rect 318352 340054 318734 340082
rect 318812 340054 319378 340082
rect 319548 340054 320022 340082
rect 320284 340054 320574 340082
rect 320928 340054 321218 340082
rect 321572 340054 321862 340082
rect 322124 340054 322414 340082
rect 322952 340054 323058 340082
rect 323228 340054 323702 340082
rect 323872 340054 324254 340082
rect 324332 340054 324898 340082
rect 325068 340054 325542 340082
rect 325804 340054 326094 340082
rect 326448 340054 326738 340082
rect 327092 340054 327382 340082
rect 327460 340054 327934 340082
rect 328472 340054 328578 340082
rect 328748 340054 329222 340082
rect 329392 340054 329774 340082
rect 329852 340054 330418 340082
rect 330588 340054 331062 340082
rect 331232 340054 331614 340082
rect 313464 337884 313516 337890
rect 313464 337826 313516 337832
rect 313476 14278 313504 337826
rect 313464 14272 313516 14278
rect 313464 14214 313516 14220
rect 313372 12028 313424 12034
rect 313372 11970 313424 11976
rect 311900 9988 311952 9994
rect 311900 9930 311952 9936
rect 313568 6866 313596 340054
rect 314120 337890 314148 340054
rect 314108 337884 314160 337890
rect 314108 337826 314160 337832
rect 314660 337884 314712 337890
rect 314660 337826 314712 337832
rect 314566 134464 314622 134473
rect 314566 134399 314622 134408
rect 314580 134201 314608 134399
rect 314566 134192 314622 134201
rect 314566 134127 314622 134136
rect 313556 6860 313608 6866
rect 313556 6802 313608 6808
rect 312176 6588 312228 6594
rect 312176 6530 312228 6536
rect 309784 3732 309836 3738
rect 309784 3674 309836 3680
rect 309784 3188 309836 3194
rect 309784 3130 309836 3136
rect 309796 480 309824 3130
rect 310980 2848 311032 2854
rect 310980 2790 311032 2796
rect 310992 480 311020 2790
rect 312188 480 312216 6530
rect 314672 6202 314700 337826
rect 314764 12102 314792 340054
rect 315408 337890 315436 340054
rect 316040 337952 316092 337958
rect 316040 337894 316092 337900
rect 315396 337884 315448 337890
rect 315396 337826 315448 337832
rect 316052 12170 316080 337894
rect 316144 14210 316172 340054
rect 316696 337958 316724 340054
rect 316684 337952 316736 337958
rect 316684 337894 316736 337900
rect 316684 337204 316736 337210
rect 316684 337146 316736 337152
rect 316132 14204 316184 14210
rect 316132 14146 316184 14152
rect 316040 12164 316092 12170
rect 316040 12106 316092 12112
rect 314752 12096 314804 12102
rect 314752 12038 314804 12044
rect 314580 6174 314700 6202
rect 314580 6118 314608 6174
rect 314568 6112 314620 6118
rect 314568 6054 314620 6060
rect 314660 6112 314712 6118
rect 314660 6054 314712 6060
rect 314672 4214 314700 6054
rect 316592 5976 316644 5982
rect 316592 5918 316644 5924
rect 315764 5500 315816 5506
rect 315764 5442 315816 5448
rect 314660 4208 314712 4214
rect 314660 4150 314712 4156
rect 314568 4140 314620 4146
rect 314568 4082 314620 4088
rect 313372 3120 313424 3126
rect 313372 3062 313424 3068
rect 313384 480 313412 3062
rect 314580 480 314608 4082
rect 315776 480 315804 5442
rect 316604 3806 316632 5918
rect 316696 4146 316724 337146
rect 317432 6050 317460 340054
rect 317604 337952 317656 337958
rect 317604 337894 317656 337900
rect 317510 170096 317566 170105
rect 317510 170031 317566 170040
rect 317524 169833 317552 170031
rect 317510 169824 317566 169833
rect 317510 169759 317566 169768
rect 317616 12238 317644 337894
rect 317604 12232 317656 12238
rect 317604 12174 317656 12180
rect 317708 9042 317736 340054
rect 318352 337958 318380 340054
rect 318340 337952 318392 337958
rect 318340 337894 318392 337900
rect 317696 9036 317748 9042
rect 317696 8978 317748 8984
rect 318812 6882 318840 340054
rect 319548 337770 319576 340054
rect 320180 337952 320232 337958
rect 320180 337894 320232 337900
rect 318996 337742 319576 337770
rect 318996 326194 319024 337742
rect 318984 326188 319036 326194
rect 318984 326130 319036 326136
rect 319168 317484 319220 317490
rect 319168 317426 319220 317432
rect 319180 309262 319208 317426
rect 319168 309256 319220 309262
rect 319168 309198 319220 309204
rect 318984 309120 319036 309126
rect 318984 309062 319036 309068
rect 318996 299418 319024 309062
rect 318904 299390 319024 299418
rect 318904 294522 318932 299390
rect 318904 294494 319116 294522
rect 319088 282826 319116 294494
rect 318996 282798 319116 282826
rect 318996 280158 319024 282798
rect 318984 280152 319036 280158
rect 318984 280094 319036 280100
rect 319076 280152 319128 280158
rect 319076 280094 319128 280100
rect 319088 263514 319116 280094
rect 318996 263486 319116 263514
rect 318996 260846 319024 263486
rect 318984 260840 319036 260846
rect 318984 260782 319036 260788
rect 319076 260840 319128 260846
rect 319076 260782 319128 260788
rect 319088 244202 319116 260782
rect 318996 244174 319116 244202
rect 318996 231878 319024 244174
rect 318984 231872 319036 231878
rect 318984 231814 319036 231820
rect 319076 231872 319128 231878
rect 319076 231814 319128 231820
rect 319088 224890 319116 231814
rect 318996 224862 319116 224890
rect 318996 212566 319024 224862
rect 318984 212560 319036 212566
rect 318984 212502 319036 212508
rect 319076 212560 319128 212566
rect 319076 212502 319128 212508
rect 319088 205578 319116 212502
rect 318996 205550 319116 205578
rect 318996 196058 319024 205550
rect 318904 196030 319024 196058
rect 318904 195974 318932 196030
rect 318892 195968 318944 195974
rect 318892 195910 318944 195916
rect 319076 195968 319128 195974
rect 319076 195910 319128 195916
rect 319088 183598 319116 195910
rect 318984 183592 319036 183598
rect 318984 183534 319036 183540
rect 319076 183592 319128 183598
rect 319076 183534 319128 183540
rect 318996 182170 319024 183534
rect 318984 182164 319036 182170
rect 318984 182106 319036 182112
rect 319076 182164 319128 182170
rect 319076 182106 319128 182112
rect 319088 166954 319116 182106
rect 318996 166926 319116 166954
rect 318996 157434 319024 166926
rect 318904 157406 319024 157434
rect 318904 157350 318932 157406
rect 318892 157344 318944 157350
rect 318892 157286 318944 157292
rect 319076 157344 319128 157350
rect 319076 157286 319128 157292
rect 319088 153202 319116 157286
rect 318984 153196 319036 153202
rect 318984 153138 319036 153144
rect 319076 153196 319128 153202
rect 319076 153138 319128 153144
rect 318996 138038 319024 153138
rect 318984 138032 319036 138038
rect 318984 137974 319036 137980
rect 319076 137964 319128 137970
rect 319076 137906 319128 137912
rect 319088 128330 319116 137906
rect 318996 128302 319116 128330
rect 318996 118794 319024 128302
rect 318984 118788 319036 118794
rect 318984 118730 319036 118736
rect 318984 104916 319036 104922
rect 318984 104858 319036 104864
rect 318996 99414 319024 104858
rect 318984 99408 319036 99414
rect 318984 99350 319036 99356
rect 319076 99340 319128 99346
rect 319076 99282 319128 99288
rect 319088 89706 319116 99282
rect 318996 89678 319116 89706
rect 318996 86970 319024 89678
rect 318984 86964 319036 86970
rect 318984 86906 319036 86912
rect 319076 86896 319128 86902
rect 319076 86838 319128 86844
rect 319088 67658 319116 86838
rect 319076 67652 319128 67658
rect 319076 67594 319128 67600
rect 319076 66292 319128 66298
rect 318996 66252 319076 66280
rect 318996 60042 319024 66252
rect 319076 66234 319128 66240
rect 318984 60036 319036 60042
rect 318984 59978 319036 59984
rect 318984 46980 319036 46986
rect 318984 46922 319036 46928
rect 318996 46866 319024 46922
rect 318996 46838 319116 46866
rect 319088 31822 319116 46838
rect 319076 31816 319128 31822
rect 319076 31758 319128 31764
rect 319076 31680 319128 31686
rect 319076 31622 319128 31628
rect 319088 26058 319116 31622
rect 318996 26030 319116 26058
rect 318996 14498 319024 26030
rect 318904 14470 319024 14498
rect 318904 9110 318932 14470
rect 318892 9104 318944 9110
rect 318892 9046 318944 9052
rect 318812 6854 318932 6882
rect 318800 6724 318852 6730
rect 318800 6666 318852 6672
rect 317420 6044 317472 6050
rect 317420 5986 317472 5992
rect 316684 4140 316736 4146
rect 316684 4082 316736 4088
rect 316960 3868 317012 3874
rect 316960 3810 317012 3816
rect 316592 3800 316644 3806
rect 316592 3742 316644 3748
rect 316972 480 317000 3810
rect 318064 3800 318116 3806
rect 318064 3742 318116 3748
rect 318076 480 318104 3742
rect 318812 3398 318840 6666
rect 318904 5914 318932 6854
rect 320192 6798 320220 337894
rect 320284 12306 320312 340054
rect 320928 337958 320956 340054
rect 320916 337952 320968 337958
rect 320916 337894 320968 337900
rect 320272 12300 320324 12306
rect 320272 12242 320324 12248
rect 321572 9178 321600 340054
rect 322124 331242 322152 340054
rect 322756 338020 322808 338026
rect 322756 337962 322808 337968
rect 321756 331214 322152 331242
rect 321756 196058 321784 331214
rect 321664 196030 321784 196058
rect 321664 195922 321692 196030
rect 321664 195894 321784 195922
rect 321756 186386 321784 195894
rect 321744 186380 321796 186386
rect 321744 186322 321796 186328
rect 321652 186312 321704 186318
rect 321652 186254 321704 186260
rect 321664 176730 321692 186254
rect 321652 176724 321704 176730
rect 321652 176666 321704 176672
rect 321744 176588 321796 176594
rect 321744 176530 321796 176536
rect 321756 157434 321784 176530
rect 321664 157406 321784 157434
rect 321664 157298 321692 157406
rect 321664 157270 321784 157298
rect 321756 153202 321784 157270
rect 321744 153196 321796 153202
rect 321744 153138 321796 153144
rect 321744 143608 321796 143614
rect 321744 143550 321796 143556
rect 321756 132682 321784 143550
rect 321664 132654 321784 132682
rect 321664 132546 321692 132654
rect 321664 132518 321784 132546
rect 321756 132462 321784 132518
rect 321744 132456 321796 132462
rect 321744 132398 321796 132404
rect 321744 122868 321796 122874
rect 321744 122810 321796 122816
rect 321756 118794 321784 122810
rect 321744 118788 321796 118794
rect 321744 118730 321796 118736
rect 321744 118652 321796 118658
rect 321744 118594 321796 118600
rect 321756 99482 321784 118594
rect 321744 99476 321796 99482
rect 321744 99418 321796 99424
rect 321744 99340 321796 99346
rect 321744 99282 321796 99288
rect 321756 72434 321784 99282
rect 321664 72406 321784 72434
rect 321664 58154 321692 72406
rect 321664 58126 321784 58154
rect 321756 57882 321784 58126
rect 321664 57854 321784 57882
rect 321664 27606 321692 57854
rect 321652 27600 321704 27606
rect 321652 27542 321704 27548
rect 321744 18012 321796 18018
rect 321744 17954 321796 17960
rect 321756 12374 321784 17954
rect 321744 12368 321796 12374
rect 321744 12310 321796 12316
rect 321560 9172 321612 9178
rect 321560 9114 321612 9120
rect 322572 9172 322624 9178
rect 322572 9114 322624 9120
rect 320180 6792 320232 6798
rect 320180 6734 320232 6740
rect 320180 6656 320232 6662
rect 320180 6598 320232 6604
rect 318892 5908 318944 5914
rect 318892 5850 318944 5856
rect 319260 4548 319312 4554
rect 319260 4490 319312 4496
rect 318800 3392 318852 3398
rect 318800 3334 318852 3340
rect 319272 480 319300 4490
rect 320192 3262 320220 6598
rect 321652 4140 321704 4146
rect 321652 4082 321704 4088
rect 320180 3256 320232 3262
rect 320180 3198 320232 3204
rect 320456 3052 320508 3058
rect 320456 2994 320508 3000
rect 320468 480 320496 2994
rect 321664 480 321692 4082
rect 322584 3942 322612 9114
rect 322664 5840 322716 5846
rect 322664 5782 322716 5788
rect 322676 4078 322704 5782
rect 322768 4146 322796 337962
rect 322952 6050 322980 340054
rect 323124 335640 323176 335646
rect 323124 335582 323176 335588
rect 323136 12442 323164 335582
rect 323124 12436 323176 12442
rect 323124 12378 323176 12384
rect 323228 9246 323256 340054
rect 323872 335646 323900 340054
rect 323860 335640 323912 335646
rect 323860 335582 323912 335588
rect 324226 318744 324282 318753
rect 324226 318679 324282 318688
rect 324240 309194 324268 318679
rect 324228 309188 324280 309194
rect 324228 309130 324280 309136
rect 324228 245472 324280 245478
rect 324228 245414 324280 245420
rect 324240 236706 324268 245414
rect 324228 236700 324280 236706
rect 324228 236642 324280 236648
rect 324228 191752 324280 191758
rect 324228 191694 324280 191700
rect 324240 182209 324268 191694
rect 324226 182200 324282 182209
rect 324226 182135 324282 182144
rect 324228 175432 324280 175438
rect 324228 175374 324280 175380
rect 324240 171193 324268 175374
rect 324226 171184 324282 171193
rect 324226 171119 324282 171128
rect 324226 122768 324282 122777
rect 324226 122703 324282 122712
rect 324240 118046 324268 122703
rect 324228 118040 324280 118046
rect 324228 117982 324280 117988
rect 323582 16960 323638 16969
rect 323504 16918 323582 16946
rect 323504 16833 323532 16918
rect 323582 16895 323638 16904
rect 323490 16824 323546 16833
rect 323490 16759 323546 16768
rect 323216 9240 323268 9246
rect 323216 9182 323268 9188
rect 323584 9036 323636 9042
rect 323584 8978 323636 8984
rect 322940 6044 322992 6050
rect 322940 5986 322992 5992
rect 322848 4480 322900 4486
rect 322848 4422 322900 4428
rect 322756 4140 322808 4146
rect 322756 4082 322808 4088
rect 322664 4072 322716 4078
rect 322664 4014 322716 4020
rect 322572 3936 322624 3942
rect 322572 3878 322624 3884
rect 322860 480 322888 4422
rect 323596 3194 323624 8978
rect 324332 5778 324360 340054
rect 325068 333334 325096 340054
rect 324412 333328 324464 333334
rect 324412 333270 324464 333276
rect 325056 333328 325108 333334
rect 325056 333270 325108 333276
rect 324424 328522 324452 333270
rect 325700 332784 325752 332790
rect 325700 332726 325752 332732
rect 324424 328494 324544 328522
rect 324516 321638 324544 328494
rect 324504 321632 324556 321638
rect 324504 321574 324556 321580
rect 324412 321564 324464 321570
rect 324412 321506 324464 321512
rect 324424 318753 324452 321506
rect 324410 318744 324466 318753
rect 324410 318679 324466 318688
rect 324504 309188 324556 309194
rect 324504 309130 324556 309136
rect 324516 302410 324544 309130
rect 324516 302382 324636 302410
rect 324608 302138 324636 302382
rect 324516 302110 324636 302138
rect 324516 299402 324544 302110
rect 324504 299396 324556 299402
rect 324504 299338 324556 299344
rect 324504 289876 324556 289882
rect 324504 289818 324556 289824
rect 324516 289785 324544 289818
rect 324502 289776 324558 289785
rect 324502 289711 324558 289720
rect 324686 289776 324742 289785
rect 324686 289711 324742 289720
rect 324700 280226 324728 289711
rect 324412 280220 324464 280226
rect 324412 280162 324464 280168
rect 324688 280220 324740 280226
rect 324688 280162 324740 280168
rect 324424 280106 324452 280162
rect 324424 280078 324544 280106
rect 324516 276706 324544 280078
rect 324424 276678 324544 276706
rect 324424 263634 324452 276678
rect 324412 263628 324464 263634
rect 324412 263570 324464 263576
rect 324412 260908 324464 260914
rect 324412 260850 324464 260856
rect 324424 260794 324452 260850
rect 324424 260766 324544 260794
rect 324516 255898 324544 260766
rect 324424 255870 324544 255898
rect 324424 245478 324452 255870
rect 324412 245472 324464 245478
rect 324412 245414 324464 245420
rect 324412 236700 324464 236706
rect 324412 236642 324464 236648
rect 324424 225010 324452 236642
rect 324412 225004 324464 225010
rect 324412 224946 324464 224952
rect 324412 222284 324464 222290
rect 324412 222226 324464 222232
rect 324424 222154 324452 222226
rect 324412 222148 324464 222154
rect 324412 222090 324464 222096
rect 324412 219564 324464 219570
rect 324412 219506 324464 219512
rect 324424 205698 324452 219506
rect 324412 205692 324464 205698
rect 324412 205634 324464 205640
rect 324412 202904 324464 202910
rect 324412 202846 324464 202852
rect 324424 196110 324452 202846
rect 324412 196104 324464 196110
rect 324412 196046 324464 196052
rect 324412 191888 324464 191894
rect 324412 191830 324464 191836
rect 324424 191758 324452 191830
rect 324412 191752 324464 191758
rect 324412 191694 324464 191700
rect 324502 182200 324558 182209
rect 324502 182135 324558 182144
rect 324516 175438 324544 182135
rect 324504 175432 324556 175438
rect 324504 175374 324556 175380
rect 324410 171184 324466 171193
rect 324466 171142 324544 171170
rect 324410 171119 324466 171128
rect 324516 171086 324544 171142
rect 324504 171080 324556 171086
rect 324504 171022 324556 171028
rect 324504 161492 324556 161498
rect 324504 161434 324556 161440
rect 324516 161378 324544 161434
rect 324516 161350 324728 161378
rect 324700 151858 324728 161350
rect 324608 151830 324728 151858
rect 324608 151774 324636 151830
rect 324596 151768 324648 151774
rect 324596 151710 324648 151716
rect 324596 142180 324648 142186
rect 324596 142122 324648 142128
rect 324608 133770 324636 142122
rect 325606 133920 325662 133929
rect 325606 133855 325608 133864
rect 325660 133855 325662 133864
rect 325608 133826 325660 133832
rect 324516 133742 324636 133770
rect 324516 132462 324544 133742
rect 324504 132456 324556 132462
rect 324504 132398 324556 132404
rect 324412 122868 324464 122874
rect 324412 122810 324464 122816
rect 324424 122777 324452 122810
rect 324410 122768 324466 122777
rect 324410 122703 324466 122712
rect 324412 118040 324464 118046
rect 324412 117982 324464 117988
rect 324424 104854 324452 117982
rect 324412 104848 324464 104854
rect 324412 104790 324464 104796
rect 324688 104848 324740 104854
rect 324688 104790 324740 104796
rect 324700 95305 324728 104790
rect 324502 95296 324558 95305
rect 324502 95231 324558 95240
rect 324686 95296 324742 95305
rect 324686 95231 324742 95240
rect 324516 95198 324544 95231
rect 324504 95192 324556 95198
rect 324504 95134 324556 95140
rect 324504 85604 324556 85610
rect 324504 85546 324556 85552
rect 324516 67658 324544 85546
rect 324412 67652 324464 67658
rect 324412 67594 324464 67600
rect 324504 67652 324556 67658
rect 324504 67594 324556 67600
rect 324424 57934 324452 67594
rect 324412 57928 324464 57934
rect 324412 57870 324464 57876
rect 324504 45620 324556 45626
rect 324504 45562 324556 45568
rect 324516 26382 324544 45562
rect 324504 26376 324556 26382
rect 324504 26318 324556 26324
rect 324412 26308 324464 26314
rect 324412 26250 324464 26256
rect 324424 19378 324452 26250
rect 324412 19372 324464 19378
rect 324412 19314 324464 19320
rect 324504 19372 324556 19378
rect 324504 19314 324556 19320
rect 324516 14498 324544 19314
rect 324424 14470 324544 14498
rect 324424 9314 324452 14470
rect 324412 9308 324464 9314
rect 324412 9250 324464 9256
rect 325516 9172 325568 9178
rect 325516 9114 325568 9120
rect 325332 5908 325384 5914
rect 325332 5850 325384 5856
rect 324320 5772 324372 5778
rect 324320 5714 324372 5720
rect 325240 3936 325292 3942
rect 325240 3878 325292 3884
rect 324044 3392 324096 3398
rect 324044 3334 324096 3340
rect 323584 3188 323636 3194
rect 323584 3130 323636 3136
rect 324056 480 324084 3334
rect 325252 480 325280 3878
rect 325344 3738 325372 5850
rect 325332 3732 325384 3738
rect 325332 3674 325384 3680
rect 325528 3126 325556 9114
rect 325608 6792 325660 6798
rect 325608 6734 325660 6740
rect 325620 3330 325648 6734
rect 325712 5710 325740 332726
rect 325804 11694 325832 340054
rect 326448 332790 326476 340054
rect 326436 332784 326488 332790
rect 326436 332726 326488 332732
rect 326068 169856 326120 169862
rect 326066 169824 326068 169833
rect 326120 169824 326122 169833
rect 326066 169759 326122 169768
rect 325792 11688 325844 11694
rect 325792 11630 325844 11636
rect 327092 9382 327120 340054
rect 327460 328681 327488 340054
rect 327446 328672 327502 328681
rect 327446 328607 327502 328616
rect 327170 328536 327226 328545
rect 327170 328471 327226 328480
rect 327184 321314 327212 328471
rect 327184 321286 327304 321314
rect 327276 318782 327304 321286
rect 327264 318776 327316 318782
rect 327264 318718 327316 318724
rect 327264 309188 327316 309194
rect 327264 309130 327316 309136
rect 327276 292670 327304 309130
rect 327264 292664 327316 292670
rect 327264 292606 327316 292612
rect 327264 292528 327316 292534
rect 327264 292470 327316 292476
rect 327276 280158 327304 292470
rect 327264 280152 327316 280158
rect 327264 280094 327316 280100
rect 327264 272196 327316 272202
rect 327264 272138 327316 272144
rect 327276 260846 327304 272138
rect 327264 260840 327316 260846
rect 327264 260782 327316 260788
rect 327264 251252 327316 251258
rect 327264 251194 327316 251200
rect 327276 241482 327304 251194
rect 327276 241454 327396 241482
rect 327368 234666 327396 241454
rect 327356 234660 327408 234666
rect 327356 234602 327408 234608
rect 327264 234592 327316 234598
rect 327264 234534 327316 234540
rect 327276 222170 327304 234534
rect 327276 222142 327396 222170
rect 327368 215354 327396 222142
rect 327356 215348 327408 215354
rect 327356 215290 327408 215296
rect 327264 215280 327316 215286
rect 327264 215222 327316 215228
rect 327276 196602 327304 215222
rect 327276 196574 327396 196602
rect 327368 193322 327396 196574
rect 327356 193316 327408 193322
rect 327356 193258 327408 193264
rect 327356 193180 327408 193186
rect 327356 193122 327408 193128
rect 327368 188154 327396 193122
rect 327172 188148 327224 188154
rect 327172 188090 327224 188096
rect 327356 188148 327408 188154
rect 327356 188090 327408 188096
rect 327184 176730 327212 188090
rect 327172 176724 327224 176730
rect 327172 176666 327224 176672
rect 327264 176588 327316 176594
rect 327264 176530 327316 176536
rect 327276 157434 327304 176530
rect 327184 157406 327304 157434
rect 327184 157298 327212 157406
rect 327184 157270 327304 157298
rect 327276 147694 327304 157270
rect 327264 147688 327316 147694
rect 327264 147630 327316 147636
rect 327172 147620 327224 147626
rect 327172 147562 327224 147568
rect 327184 135318 327212 147562
rect 327172 135312 327224 135318
rect 327172 135254 327224 135260
rect 327172 132524 327224 132530
rect 327172 132466 327224 132472
rect 327184 124273 327212 132466
rect 327170 124264 327226 124273
rect 327170 124199 327226 124208
rect 327170 123992 327226 124001
rect 327170 123927 327226 123936
rect 327184 114510 327212 123927
rect 327172 114504 327224 114510
rect 327172 114446 327224 114452
rect 327264 104916 327316 104922
rect 327264 104858 327316 104864
rect 327276 99550 327304 104858
rect 327264 99544 327316 99550
rect 327264 99486 327316 99492
rect 327264 99340 327316 99346
rect 327264 99282 327316 99288
rect 327276 95198 327304 99282
rect 327264 95192 327316 95198
rect 327264 95134 327316 95140
rect 327264 85604 327316 85610
rect 327264 85546 327316 85552
rect 327276 77382 327304 85546
rect 327264 77376 327316 77382
rect 327264 77318 327316 77324
rect 327172 77240 327224 77246
rect 327172 77182 327224 77188
rect 327184 75886 327212 77182
rect 327172 75880 327224 75886
rect 327172 75822 327224 75828
rect 327264 66292 327316 66298
rect 327264 66234 327316 66240
rect 327276 48414 327304 66234
rect 327264 48408 327316 48414
rect 327264 48350 327316 48356
rect 327172 48340 327224 48346
rect 327172 48282 327224 48288
rect 327184 27674 327212 48282
rect 327172 27668 327224 27674
rect 327172 27610 327224 27616
rect 327264 27668 327316 27674
rect 327264 27610 327316 27616
rect 327276 11626 327304 27610
rect 327264 11620 327316 11626
rect 327264 11562 327316 11568
rect 327080 9376 327132 9382
rect 327080 9318 327132 9324
rect 327080 9240 327132 9246
rect 327080 9182 327132 9188
rect 325700 5704 325752 5710
rect 325700 5646 325752 5652
rect 326436 4412 326488 4418
rect 326436 4354 326488 4360
rect 325608 3324 325660 3330
rect 325608 3266 325660 3272
rect 325516 3120 325568 3126
rect 325516 3062 325568 3068
rect 326448 480 326476 4354
rect 327092 3874 327120 9182
rect 328472 5642 328500 340054
rect 328644 335640 328696 335646
rect 328644 335582 328696 335588
rect 328656 11558 328684 335582
rect 328644 11552 328696 11558
rect 328644 11494 328696 11500
rect 328748 9450 328776 340054
rect 329392 335646 329420 340054
rect 329380 335640 329432 335646
rect 329380 335582 329432 335588
rect 328736 9444 328788 9450
rect 328736 9386 328788 9392
rect 328552 9104 328604 9110
rect 328552 9046 328604 9052
rect 328460 5636 328512 5642
rect 328460 5578 328512 5584
rect 327080 3868 327132 3874
rect 327080 3810 327132 3816
rect 327632 3188 327684 3194
rect 327632 3130 327684 3136
rect 327644 480 327672 3130
rect 328564 3058 328592 9046
rect 329852 5574 329880 340054
rect 330588 328506 330616 340054
rect 330024 328500 330076 328506
rect 330024 328442 330076 328448
rect 330576 328500 330628 328506
rect 330576 328442 330628 328448
rect 330036 292670 330064 328442
rect 330024 292664 330076 292670
rect 330024 292606 330076 292612
rect 330024 292528 330076 292534
rect 330024 292470 330076 292476
rect 330036 273358 330064 292470
rect 331128 280152 331180 280158
rect 331128 280094 331180 280100
rect 330024 273352 330076 273358
rect 330024 273294 330076 273300
rect 330024 273216 330076 273222
rect 330024 273158 330076 273164
rect 330036 254046 330064 273158
rect 331140 270609 331168 280094
rect 331126 270600 331182 270609
rect 331126 270535 331182 270544
rect 331128 260840 331180 260846
rect 331128 260782 331180 260788
rect 330024 254040 330076 254046
rect 330024 253982 330076 253988
rect 330024 253904 330076 253910
rect 330024 253846 330076 253852
rect 330036 241482 330064 253846
rect 331140 251297 331168 260782
rect 331126 251288 331182 251297
rect 331126 251223 331182 251232
rect 331126 251152 331182 251161
rect 331126 251087 331182 251096
rect 331140 241534 331168 251087
rect 331128 241528 331180 241534
rect 330036 241454 330156 241482
rect 331128 241470 331180 241476
rect 330128 234666 330156 241454
rect 330116 234660 330168 234666
rect 330116 234602 330168 234608
rect 330024 234592 330076 234598
rect 330024 234534 330076 234540
rect 330036 222170 330064 234534
rect 330036 222142 330156 222170
rect 330128 215354 330156 222142
rect 331128 219428 331180 219434
rect 331128 219370 331180 219376
rect 330116 215348 330168 215354
rect 330116 215290 330168 215296
rect 330024 215280 330076 215286
rect 330024 215222 330076 215228
rect 330036 202858 330064 215222
rect 331140 209817 331168 219370
rect 331126 209808 331182 209817
rect 331126 209743 331182 209752
rect 330036 202830 330156 202858
rect 330128 196042 330156 202830
rect 331036 196648 331088 196654
rect 331036 196590 331088 196596
rect 330116 196036 330168 196042
rect 330116 195978 330168 195984
rect 330024 195968 330076 195974
rect 330024 195910 330076 195916
rect 330036 157434 330064 195910
rect 331048 193202 331076 196590
rect 331232 193322 331260 340054
rect 331692 328506 331720 340190
rect 332612 340054 332902 340082
rect 333164 340054 333454 340082
rect 332508 338088 332560 338094
rect 332508 338030 332560 338036
rect 331496 328500 331548 328506
rect 331496 328442 331548 328448
rect 331680 328500 331732 328506
rect 331680 328442 331732 328448
rect 331508 309210 331536 328442
rect 331416 309182 331536 309210
rect 331416 302002 331444 309182
rect 331416 301974 331536 302002
rect 331508 299470 331536 301974
rect 331404 299464 331456 299470
rect 331404 299406 331456 299412
rect 331496 299464 331548 299470
rect 331496 299406 331548 299412
rect 331416 298110 331444 299406
rect 331404 298104 331456 298110
rect 331404 298046 331456 298052
rect 331404 288448 331456 288454
rect 331404 288390 331456 288396
rect 331416 282946 331444 288390
rect 331404 282940 331456 282946
rect 331404 282882 331456 282888
rect 331496 282804 331548 282810
rect 331496 282746 331548 282752
rect 331508 280158 331536 282746
rect 331496 280152 331548 280158
rect 331496 280094 331548 280100
rect 331310 270464 331366 270473
rect 331310 270399 331366 270408
rect 331324 263566 331352 270399
rect 331312 263560 331364 263566
rect 331312 263502 331364 263508
rect 331496 263492 331548 263498
rect 331496 263434 331548 263440
rect 331508 260846 331536 263434
rect 331496 260840 331548 260846
rect 331496 260782 331548 260788
rect 331496 241528 331548 241534
rect 331496 241470 331548 241476
rect 331508 231878 331536 241470
rect 331496 231872 331548 231878
rect 331496 231814 331548 231820
rect 331496 231736 331548 231742
rect 331496 231678 331548 231684
rect 331508 222306 331536 231678
rect 331508 222278 331628 222306
rect 331600 220862 331628 222278
rect 331312 220856 331364 220862
rect 331312 220798 331364 220804
rect 331588 220856 331640 220862
rect 331588 220798 331640 220804
rect 331324 219434 331352 220798
rect 331312 219428 331364 219434
rect 331312 219370 331364 219376
rect 331494 209808 331550 209817
rect 331494 209743 331550 209752
rect 331508 202978 331536 209743
rect 331496 202972 331548 202978
rect 331496 202914 331548 202920
rect 331404 201544 331456 201550
rect 331404 201486 331456 201492
rect 331416 196654 331444 201486
rect 331404 196648 331456 196654
rect 331404 196590 331456 196596
rect 331220 193316 331272 193322
rect 331220 193258 331272 193264
rect 331048 193174 331168 193202
rect 331140 183598 331168 193174
rect 331220 193180 331272 193186
rect 331220 193122 331272 193128
rect 331128 183592 331180 183598
rect 331128 183534 331180 183540
rect 329944 157406 330064 157434
rect 329944 157298 329972 157406
rect 329944 157270 330064 157298
rect 330036 137306 330064 157270
rect 330036 137278 330248 137306
rect 330220 135289 330248 137278
rect 330206 135280 330262 135289
rect 330206 135215 330262 135224
rect 329930 135144 329986 135153
rect 329930 135079 329986 135088
rect 329944 125610 329972 135079
rect 329944 125582 330064 125610
rect 330036 118776 330064 125582
rect 330036 118748 330156 118776
rect 330128 118538 330156 118748
rect 330036 118510 330156 118538
rect 330036 106282 330064 118510
rect 330024 106276 330076 106282
rect 330024 106218 330076 106224
rect 330208 106276 330260 106282
rect 330208 106218 330260 106224
rect 330220 95282 330248 106218
rect 330128 95254 330248 95282
rect 330128 85610 330156 95254
rect 330024 85604 330076 85610
rect 330024 85546 330076 85552
rect 330116 85604 330168 85610
rect 330116 85546 330168 85552
rect 330036 76090 330064 85546
rect 330024 76084 330076 76090
rect 330024 76026 330076 76032
rect 330116 75948 330168 75954
rect 330116 75890 330168 75896
rect 330128 75834 330156 75890
rect 330036 75806 330156 75834
rect 330036 66298 330064 75806
rect 330024 66292 330076 66298
rect 330024 66234 330076 66240
rect 330024 65000 330076 65006
rect 330024 64942 330076 64948
rect 330036 63510 330064 64942
rect 330024 63504 330076 63510
rect 330024 63446 330076 63452
rect 329932 53848 329984 53854
rect 329932 53790 329984 53796
rect 329944 45665 329972 53790
rect 329930 45656 329986 45665
rect 329930 45591 329986 45600
rect 330114 45520 330170 45529
rect 330114 45455 330170 45464
rect 330128 14550 330156 45455
rect 329932 14544 329984 14550
rect 329932 14486 329984 14492
rect 330116 14544 330168 14550
rect 330116 14486 330168 14492
rect 329944 9602 329972 14486
rect 331232 11490 331260 193122
rect 331496 183592 331548 183598
rect 331496 183534 331548 183540
rect 331508 172689 331536 183534
rect 331494 172680 331550 172689
rect 331494 172615 331550 172624
rect 331402 172544 331458 172553
rect 331402 172479 331458 172488
rect 331310 170096 331366 170105
rect 331310 170031 331366 170040
rect 331324 169862 331352 170031
rect 331312 169856 331364 169862
rect 331312 169798 331364 169804
rect 331416 161430 331444 172479
rect 331404 161424 331456 161430
rect 331404 161366 331456 161372
rect 331404 151836 331456 151842
rect 331404 151778 331456 151784
rect 331416 147762 331444 151778
rect 331404 147756 331456 147762
rect 331404 147698 331456 147704
rect 331404 147620 331456 147626
rect 331404 147562 331456 147568
rect 331416 144922 331444 147562
rect 331416 144894 331536 144922
rect 331508 135266 331536 144894
rect 331416 135238 331536 135266
rect 331416 125610 331444 135238
rect 331416 125582 331536 125610
rect 331508 118946 331536 125582
rect 331508 118918 331628 118946
rect 331600 118674 331628 118918
rect 331508 118646 331628 118674
rect 331508 106282 331536 118646
rect 331404 106276 331456 106282
rect 331404 106218 331456 106224
rect 331496 106276 331548 106282
rect 331496 106218 331548 106224
rect 331416 86902 331444 106218
rect 331404 86896 331456 86902
rect 331404 86838 331456 86844
rect 331404 77308 331456 77314
rect 331404 77250 331456 77256
rect 331416 55690 331444 77250
rect 331404 55684 331456 55690
rect 331404 55626 331456 55632
rect 331496 48340 331548 48346
rect 331496 48282 331548 48288
rect 331508 37398 331536 48282
rect 331496 37392 331548 37398
rect 331496 37334 331548 37340
rect 331404 37324 331456 37330
rect 331404 37266 331456 37272
rect 331416 13054 331444 37266
rect 331404 13048 331456 13054
rect 331404 12990 331456 12996
rect 331220 11484 331272 11490
rect 331220 11426 331272 11432
rect 329944 9574 330064 9602
rect 330036 9518 330064 9574
rect 330024 9512 330076 9518
rect 330024 9454 330076 9460
rect 329840 5568 329892 5574
rect 329840 5510 329892 5516
rect 330024 4344 330076 4350
rect 330024 4286 330076 4292
rect 328828 3256 328880 3262
rect 328828 3198 328880 3204
rect 328552 3052 328604 3058
rect 328552 2994 328604 3000
rect 328840 480 328868 3198
rect 330036 480 330064 4286
rect 332520 4146 332548 338030
rect 332612 9586 332640 340054
rect 333164 338076 333192 340054
rect 332980 338048 333192 338076
rect 332980 328506 333008 338048
rect 334084 335442 334112 340068
rect 334268 340054 334742 340082
rect 334072 335436 334124 335442
rect 334072 335378 334124 335384
rect 334164 335232 334216 335238
rect 334164 335174 334216 335180
rect 333980 331628 334032 331634
rect 333980 331570 334032 331576
rect 332692 328500 332744 328506
rect 332692 328442 332744 328448
rect 332968 328500 333020 328506
rect 332968 328442 333020 328448
rect 332704 328409 332732 328442
rect 332690 328400 332746 328409
rect 332690 328335 332746 328344
rect 332782 318880 332838 318889
rect 332782 318815 332838 318824
rect 332796 318782 332824 318815
rect 332784 318776 332836 318782
rect 332784 318718 332836 318724
rect 332784 309188 332836 309194
rect 332784 309130 332836 309136
rect 332796 292670 332824 309130
rect 332784 292664 332836 292670
rect 332784 292606 332836 292612
rect 332784 292528 332836 292534
rect 332784 292470 332836 292476
rect 332796 273358 332824 292470
rect 332784 273352 332836 273358
rect 332784 273294 332836 273300
rect 332784 273216 332836 273222
rect 332784 273158 332836 273164
rect 332796 157434 332824 273158
rect 332704 157406 332824 157434
rect 332704 157298 332732 157406
rect 332704 157270 332824 157298
rect 332796 118810 332824 157270
rect 333886 133920 333942 133929
rect 333886 133855 333888 133864
rect 333940 133855 333942 133864
rect 333888 133826 333940 133832
rect 332704 118782 332824 118810
rect 332704 118674 332732 118782
rect 332704 118646 332824 118674
rect 332796 64870 332824 118646
rect 332784 64864 332836 64870
rect 332784 64806 332836 64812
rect 332876 64864 332928 64870
rect 332876 64806 332928 64812
rect 332888 63510 332916 64806
rect 332876 63504 332928 63510
rect 332876 63446 332928 63452
rect 332876 55208 332928 55214
rect 332876 55150 332928 55156
rect 332888 46986 332916 55150
rect 332876 46980 332928 46986
rect 332876 46922 332928 46928
rect 332876 46844 332928 46850
rect 332876 46786 332928 46792
rect 332888 45558 332916 46786
rect 332876 45552 332928 45558
rect 332876 45494 332928 45500
rect 332692 35964 332744 35970
rect 332692 35906 332744 35912
rect 332704 30138 332732 35906
rect 332704 30110 332824 30138
rect 332796 11422 332824 30110
rect 332784 11416 332836 11422
rect 332784 11358 332836 11364
rect 333992 9654 334020 331570
rect 334176 13802 334204 335174
rect 334268 331634 334296 340054
rect 334256 331628 334308 331634
rect 334256 331570 334308 331576
rect 334820 328506 334848 340190
rect 335464 340054 335938 340082
rect 336200 340054 336490 340082
rect 335360 335640 335412 335646
rect 335360 335582 335412 335588
rect 334440 328500 334492 328506
rect 334440 328442 334492 328448
rect 334808 328500 334860 328506
rect 334808 328442 334860 328448
rect 334452 309194 334480 328442
rect 334440 309188 334492 309194
rect 334440 309130 334492 309136
rect 334440 307828 334492 307834
rect 334440 307770 334492 307776
rect 334452 299470 334480 307770
rect 334256 299464 334308 299470
rect 334256 299406 334308 299412
rect 334440 299464 334492 299470
rect 334440 299406 334492 299412
rect 334268 298110 334296 299406
rect 334256 298104 334308 298110
rect 334256 298046 334308 298052
rect 334440 282804 334492 282810
rect 334440 282746 334492 282752
rect 334452 280158 334480 282746
rect 334440 280152 334492 280158
rect 334440 280094 334492 280100
rect 334348 270632 334400 270638
rect 334348 270574 334400 270580
rect 334360 263634 334388 270574
rect 334348 263628 334400 263634
rect 334348 263570 334400 263576
rect 334440 263492 334492 263498
rect 334440 263434 334492 263440
rect 334452 260846 334480 263434
rect 334440 260840 334492 260846
rect 334440 260782 334492 260788
rect 334348 251320 334400 251326
rect 334348 251262 334400 251268
rect 334360 251190 334388 251262
rect 334348 251184 334400 251190
rect 334348 251126 334400 251132
rect 334348 244180 334400 244186
rect 334348 244122 334400 244128
rect 334360 232014 334388 244122
rect 334348 232008 334400 232014
rect 334348 231950 334400 231956
rect 334440 231872 334492 231878
rect 334440 231814 334492 231820
rect 334452 226930 334480 231814
rect 334360 226902 334480 226930
rect 334360 212702 334388 226902
rect 334348 212696 334400 212702
rect 334348 212638 334400 212644
rect 334440 212560 334492 212566
rect 334440 212502 334492 212508
rect 334452 207618 334480 212502
rect 334360 207590 334480 207618
rect 334360 193390 334388 207590
rect 334348 193384 334400 193390
rect 334348 193326 334400 193332
rect 334440 193248 334492 193254
rect 334440 193190 334492 193196
rect 334452 186454 334480 193190
rect 334440 186448 334492 186454
rect 334440 186390 334492 186396
rect 334452 183598 334480 183629
rect 334440 183592 334492 183598
rect 334360 183540 334440 183546
rect 334360 183534 334492 183540
rect 334360 183518 334480 183534
rect 334360 175914 334388 183518
rect 334348 175908 334400 175914
rect 334348 175850 334400 175856
rect 334532 169788 334584 169794
rect 334532 169730 334584 169736
rect 334544 161498 334572 169730
rect 334348 161492 334400 161498
rect 334348 161434 334400 161440
rect 334532 161492 334584 161498
rect 334532 161434 334584 161440
rect 334360 161378 334388 161434
rect 334268 161350 334388 161378
rect 334268 157434 334296 161350
rect 334268 157406 334480 157434
rect 334452 156754 334480 157406
rect 334360 156726 334480 156754
rect 334360 147762 334388 156726
rect 334348 147756 334400 147762
rect 334348 147698 334400 147704
rect 334348 147620 334400 147626
rect 334348 147562 334400 147568
rect 334360 144922 334388 147562
rect 334360 144906 334480 144922
rect 334360 144900 334492 144906
rect 334360 144894 334440 144900
rect 334440 144842 334492 144848
rect 334440 135176 334492 135182
rect 334440 135118 334492 135124
rect 334452 114578 334480 135118
rect 334440 114572 334492 114578
rect 334440 114514 334492 114520
rect 334348 113212 334400 113218
rect 334348 113154 334400 113160
rect 334360 104922 334388 113154
rect 334348 104916 334400 104922
rect 334348 104858 334400 104864
rect 334440 104916 334492 104922
rect 334440 104858 334492 104864
rect 334452 103494 334480 104858
rect 334440 103488 334492 103494
rect 334440 103430 334492 103436
rect 334348 93900 334400 93906
rect 334348 93842 334400 93848
rect 334360 86902 334388 93842
rect 334348 86896 334400 86902
rect 334348 86838 334400 86844
rect 334348 77308 334400 77314
rect 334348 77250 334400 77256
rect 334360 55690 334388 77250
rect 334348 55684 334400 55690
rect 334348 55626 334400 55632
rect 334440 48340 334492 48346
rect 334440 48282 334492 48288
rect 334452 37398 334480 48282
rect 335266 40216 335322 40225
rect 335266 40151 335322 40160
rect 335280 40089 335308 40151
rect 335266 40080 335322 40089
rect 335266 40015 335322 40024
rect 334440 37392 334492 37398
rect 334440 37334 334492 37340
rect 334348 37324 334400 37330
rect 334348 37266 334400 37272
rect 334360 35902 334388 37266
rect 334348 35896 334400 35902
rect 334348 35838 334400 35844
rect 334532 26308 334584 26314
rect 334532 26250 334584 26256
rect 334544 26178 334572 26250
rect 334348 26172 334400 26178
rect 334348 26114 334400 26120
rect 334532 26172 334584 26178
rect 334532 26114 334584 26120
rect 334360 21298 334388 26114
rect 334360 21270 334480 21298
rect 334164 13796 334216 13802
rect 334164 13738 334216 13744
rect 334452 11354 334480 21270
rect 335266 17232 335322 17241
rect 335266 17167 335322 17176
rect 335280 16833 335308 17167
rect 335266 16824 335322 16833
rect 335266 16759 335322 16768
rect 334440 11348 334492 11354
rect 334440 11290 334492 11296
rect 333980 9648 334032 9654
rect 333980 9590 334032 9596
rect 332600 9580 332652 9586
rect 332600 9522 332652 9528
rect 334716 8968 334768 8974
rect 334716 8910 334768 8916
rect 333612 4276 333664 4282
rect 333612 4218 333664 4224
rect 331220 4140 331272 4146
rect 331220 4082 331272 4088
rect 332508 4140 332560 4146
rect 332508 4082 332560 4088
rect 331232 480 331260 4082
rect 332416 3868 332468 3874
rect 332416 3810 332468 3816
rect 332428 480 332456 3810
rect 333624 480 333652 4218
rect 334728 480 334756 8910
rect 335372 8838 335400 335582
rect 335464 12986 335492 340054
rect 336200 335646 336228 340054
rect 337120 337278 337148 340068
rect 337108 337272 337160 337278
rect 337108 337214 337160 337220
rect 336188 335640 336240 335646
rect 336188 335582 336240 335588
rect 337212 328506 337240 340190
rect 338224 340054 338330 340082
rect 336924 328500 336976 328506
rect 336924 328442 336976 328448
rect 337200 328500 337252 328506
rect 337200 328442 337252 328448
rect 336936 309194 336964 328442
rect 336832 309188 336884 309194
rect 336832 309130 336884 309136
rect 336924 309188 336976 309194
rect 336924 309130 336976 309136
rect 336844 302274 336872 309130
rect 336752 302246 336872 302274
rect 336752 302138 336780 302246
rect 336752 302110 336872 302138
rect 336844 282962 336872 302110
rect 336752 282934 336872 282962
rect 336752 282826 336780 282934
rect 336752 282798 336872 282826
rect 336844 263650 336872 282798
rect 336752 263622 336872 263650
rect 336752 263514 336780 263622
rect 336752 263486 336872 263514
rect 336844 244338 336872 263486
rect 336752 244310 336872 244338
rect 336752 244202 336780 244310
rect 336752 244174 336872 244202
rect 336844 225026 336872 244174
rect 336752 224998 336872 225026
rect 336752 224890 336780 224998
rect 336752 224862 336872 224890
rect 336844 205714 336872 224862
rect 336752 205686 336872 205714
rect 336752 205578 336780 205686
rect 336752 205550 336872 205578
rect 336844 186402 336872 205550
rect 336752 186374 336872 186402
rect 336752 186266 336780 186374
rect 336752 186238 336872 186266
rect 336844 167090 336872 186238
rect 338026 170096 338082 170105
rect 338026 170031 338082 170040
rect 338040 169697 338068 170031
rect 338026 169688 338082 169697
rect 338026 169623 338082 169632
rect 336752 167062 336872 167090
rect 336752 166954 336780 167062
rect 336752 166926 336872 166954
rect 336844 157350 336872 166926
rect 336832 157344 336884 157350
rect 336832 157286 336884 157292
rect 336924 157276 336976 157282
rect 336924 157218 336976 157224
rect 336936 138122 336964 157218
rect 336936 138094 337056 138122
rect 337028 137714 337056 138094
rect 336936 137686 337056 137714
rect 336936 118794 336964 137686
rect 336924 118788 336976 118794
rect 336924 118730 336976 118736
rect 336832 118720 336884 118726
rect 336832 118662 336884 118668
rect 336844 109154 336872 118662
rect 336752 109126 336872 109154
rect 336752 109018 336780 109126
rect 336752 108990 336872 109018
rect 336844 89842 336872 108990
rect 336752 89814 336872 89842
rect 336752 89706 336780 89814
rect 336752 89678 336872 89706
rect 336844 66230 336872 89678
rect 336832 66224 336884 66230
rect 336832 66166 336884 66172
rect 336924 66224 336976 66230
rect 336924 66166 336976 66172
rect 336936 56574 336964 66166
rect 336924 56568 336976 56574
rect 336924 56510 336976 56516
rect 336924 46980 336976 46986
rect 336924 46922 336976 46928
rect 336936 27606 336964 46922
rect 336924 27600 336976 27606
rect 336924 27542 336976 27548
rect 336832 18012 336884 18018
rect 336832 17954 336884 17960
rect 335452 12980 335504 12986
rect 335452 12922 335504 12928
rect 336844 12850 336872 17954
rect 336832 12844 336884 12850
rect 336832 12786 336884 12792
rect 338224 8906 338252 340054
rect 338960 337346 338988 340068
rect 339618 340054 339724 340082
rect 338948 337340 339000 337346
rect 338948 337282 339000 337288
rect 339408 337272 339460 337278
rect 339408 337214 339460 337220
rect 338212 8900 338264 8906
rect 338212 8842 338264 8848
rect 335360 8832 335412 8838
rect 335360 8774 335412 8780
rect 337108 4208 337160 4214
rect 337108 4150 337160 4156
rect 335912 3120 335964 3126
rect 335912 3062 335964 3068
rect 335924 480 335952 3062
rect 337120 480 337148 4150
rect 339420 3058 339448 337214
rect 339500 335640 339552 335646
rect 339500 335582 339552 335588
rect 339512 4758 339540 335582
rect 339696 12918 339724 340054
rect 339788 340054 340170 340082
rect 340432 340054 340814 340082
rect 340984 340054 341458 340082
rect 341720 340054 342010 340082
rect 342272 340054 342654 340082
rect 339684 12912 339736 12918
rect 339684 12854 339736 12860
rect 339788 8770 339816 340054
rect 340432 335646 340460 340054
rect 340420 335640 340472 335646
rect 340420 335582 340472 335588
rect 340880 334620 340932 334626
rect 340880 334562 340932 334568
rect 339776 8764 339828 8770
rect 339776 8706 339828 8712
rect 340892 8634 340920 334562
rect 340984 12782 341012 340054
rect 341720 334626 341748 340054
rect 341708 334620 341760 334626
rect 341708 334562 341760 334568
rect 340972 12776 341024 12782
rect 340972 12718 341024 12724
rect 340880 8628 340932 8634
rect 340880 8570 340932 8576
rect 342272 4865 342300 340054
rect 342732 338042 342760 340190
rect 342640 338014 342760 338042
rect 343744 340054 343850 340082
rect 344112 340054 344494 340082
rect 342640 331294 342668 338014
rect 343640 331560 343692 331566
rect 343640 331502 343692 331508
rect 342628 331288 342680 331294
rect 342628 331230 342680 331236
rect 342628 328500 342680 328506
rect 342628 328442 342680 328448
rect 342640 309262 342668 328442
rect 342628 309256 342680 309262
rect 342628 309198 342680 309204
rect 342444 309188 342496 309194
rect 342444 309130 342496 309136
rect 342456 309058 342484 309130
rect 342444 309052 342496 309058
rect 342444 308994 342496 309000
rect 342536 299600 342588 299606
rect 342536 299542 342588 299548
rect 342548 299452 342576 299542
rect 342548 299424 342760 299452
rect 342732 289898 342760 299424
rect 342548 289870 342760 289898
rect 342548 282946 342576 289870
rect 342536 282940 342588 282946
rect 342536 282882 342588 282888
rect 342536 280288 342588 280294
rect 342536 280230 342588 280236
rect 342548 280140 342576 280230
rect 342548 280112 342760 280140
rect 342732 270586 342760 280112
rect 342548 270558 342760 270586
rect 342548 263634 342576 270558
rect 342536 263628 342588 263634
rect 342536 263570 342588 263576
rect 342536 260908 342588 260914
rect 342536 260850 342588 260856
rect 342548 260778 342576 260850
rect 342536 260772 342588 260778
rect 342536 260714 342588 260720
rect 342444 251252 342496 251258
rect 342444 251194 342496 251200
rect 342456 251161 342484 251194
rect 342442 251152 342498 251161
rect 342442 251087 342498 251096
rect 342626 251152 342682 251161
rect 342626 251087 342682 251096
rect 342640 241516 342668 251087
rect 342640 241488 342760 241516
rect 342732 234546 342760 241488
rect 342456 234518 342760 234546
rect 342456 231849 342484 234518
rect 342442 231840 342498 231849
rect 342442 231775 342498 231784
rect 342718 231840 342774 231849
rect 342718 231775 342774 231784
rect 342732 212809 342760 231775
rect 342718 212800 342774 212809
rect 342718 212735 342774 212744
rect 342442 212562 342498 212571
rect 342498 212506 342668 212514
rect 342442 212497 342668 212506
rect 342456 212486 342668 212497
rect 342640 202910 342668 212486
rect 342628 202904 342680 202910
rect 342628 202846 342680 202852
rect 342720 202904 342772 202910
rect 342720 202846 342772 202852
rect 342732 196654 342760 202846
rect 342720 196648 342772 196654
rect 342720 196590 342772 196596
rect 342904 196648 342956 196654
rect 342904 196590 342956 196596
rect 342916 191865 342944 196590
rect 342718 191856 342774 191865
rect 342718 191791 342774 191800
rect 342902 191856 342958 191865
rect 342902 191791 342958 191800
rect 342732 172553 342760 191791
rect 342442 172544 342498 172553
rect 342442 172479 342498 172488
rect 342718 172544 342774 172553
rect 342718 172479 342774 172488
rect 342456 166682 342484 172479
rect 342456 166654 342576 166682
rect 342548 164200 342576 166654
rect 342456 164172 342576 164200
rect 342456 157434 342484 164172
rect 342364 157406 342484 157434
rect 342364 154737 342392 157406
rect 342350 154728 342406 154737
rect 342350 154663 342406 154672
rect 342442 154592 342498 154601
rect 342352 154556 342404 154562
rect 342498 154562 342576 154578
rect 342498 154556 342588 154562
rect 342498 154550 342536 154556
rect 342442 154527 342498 154536
rect 342352 154498 342404 154504
rect 342536 154498 342588 154504
rect 342364 144945 342392 154498
rect 342548 154467 342576 154498
rect 342350 144936 342406 144945
rect 342350 144871 342406 144880
rect 342534 144936 342590 144945
rect 342534 144871 342590 144880
rect 342548 138106 342576 144871
rect 342536 138100 342588 138106
rect 342536 138042 342588 138048
rect 342536 137964 342588 137970
rect 342536 137906 342588 137912
rect 342548 116113 342576 137906
rect 342534 116104 342590 116113
rect 342534 116039 342590 116048
rect 342442 115968 342498 115977
rect 342442 115903 342444 115912
rect 342496 115903 342498 115912
rect 342444 115874 342496 115880
rect 342444 108996 342496 109002
rect 342444 108938 342496 108944
rect 342456 101402 342484 108938
rect 342364 101374 342484 101402
rect 342364 99362 342392 101374
rect 342364 99334 342484 99362
rect 342456 86970 342484 99334
rect 342444 86964 342496 86970
rect 342444 86906 342496 86912
rect 342444 77308 342496 77314
rect 342444 77250 342496 77256
rect 342456 51134 342484 77250
rect 342444 51128 342496 51134
rect 342444 51070 342496 51076
rect 342444 50992 342496 50998
rect 342444 50934 342496 50940
rect 342456 46918 342484 50934
rect 342444 46912 342496 46918
rect 342444 46854 342496 46860
rect 342536 37324 342588 37330
rect 342536 37266 342588 37272
rect 342548 28948 342576 37266
rect 342364 28920 342576 28948
rect 342364 12714 342392 28920
rect 342352 12708 342404 12714
rect 342352 12650 342404 12656
rect 342258 4856 342314 4865
rect 342258 4791 342314 4800
rect 339500 4752 339552 4758
rect 339500 4694 339552 4700
rect 340696 4752 340748 4758
rect 340696 4694 340748 4700
rect 339500 4072 339552 4078
rect 339500 4014 339552 4020
rect 338304 3052 338356 3058
rect 338304 2994 338356 3000
rect 339408 3052 339460 3058
rect 339408 2994 339460 3000
rect 338316 480 338344 2994
rect 339512 480 339540 4014
rect 340708 480 340736 4694
rect 343652 4690 343680 331502
rect 343744 8702 343772 340054
rect 344112 331566 344140 340054
rect 345020 335640 345072 335646
rect 345020 335582 345072 335588
rect 344100 331560 344152 331566
rect 344100 331502 344152 331508
rect 344926 40352 344982 40361
rect 344926 40287 344982 40296
rect 344940 40089 344968 40287
rect 344926 40080 344982 40089
rect 344926 40015 344982 40024
rect 343732 8696 343784 8702
rect 343732 8638 343784 8644
rect 343640 4684 343692 4690
rect 343640 4626 343692 4632
rect 344284 4684 344336 4690
rect 344284 4626 344336 4632
rect 343088 3188 343140 3194
rect 343088 3130 343140 3136
rect 341892 2984 341944 2990
rect 341892 2926 341944 2932
rect 341904 480 341932 2926
rect 343100 480 343128 3130
rect 344296 480 344324 4626
rect 345032 4622 345060 335582
rect 345124 7206 345152 340068
rect 345216 340054 345690 340082
rect 345952 340054 346334 340082
rect 346412 340054 346978 340082
rect 347056 340054 347530 340082
rect 347792 340054 348174 340082
rect 345216 8566 345244 340054
rect 345952 335646 345980 340054
rect 346308 337272 346360 337278
rect 346308 337214 346360 337220
rect 345940 335640 345992 335646
rect 345940 335582 345992 335588
rect 346214 16688 346270 16697
rect 346214 16623 346270 16632
rect 346228 16561 346256 16623
rect 346214 16552 346270 16561
rect 346214 16487 346270 16496
rect 345204 8560 345256 8566
rect 345204 8502 345256 8508
rect 345112 7200 345164 7206
rect 345112 7142 345164 7148
rect 345020 4616 345072 4622
rect 345020 4558 345072 4564
rect 346320 746 346348 337214
rect 346412 7138 346440 340054
rect 347056 335730 347084 340054
rect 346596 335702 347084 335730
rect 346596 311846 346624 335702
rect 346584 311840 346636 311846
rect 346584 311782 346636 311788
rect 346584 309188 346636 309194
rect 346584 309130 346636 309136
rect 346596 299470 346624 309130
rect 346584 299464 346636 299470
rect 346584 299406 346636 299412
rect 346584 289876 346636 289882
rect 346584 289818 346636 289824
rect 346596 280158 346624 289818
rect 346584 280152 346636 280158
rect 346584 280094 346636 280100
rect 346584 270564 346636 270570
rect 346584 270506 346636 270512
rect 346596 260846 346624 270506
rect 346584 260840 346636 260846
rect 346584 260782 346636 260788
rect 346584 251252 346636 251258
rect 346584 251194 346636 251200
rect 346596 241505 346624 251194
rect 346582 241496 346638 241505
rect 346582 241431 346638 241440
rect 346766 241496 346822 241505
rect 346766 241431 346822 241440
rect 346780 231878 346808 241431
rect 346584 231872 346636 231878
rect 346584 231814 346636 231820
rect 346768 231872 346820 231878
rect 346768 231814 346820 231820
rect 346596 222193 346624 231814
rect 346582 222184 346638 222193
rect 346582 222119 346638 222128
rect 346766 222184 346822 222193
rect 346766 222119 346822 222128
rect 346780 212566 346808 222119
rect 346584 212560 346636 212566
rect 346584 212502 346636 212508
rect 346768 212560 346820 212566
rect 346768 212502 346820 212508
rect 346596 202881 346624 212502
rect 346582 202872 346638 202881
rect 346582 202807 346638 202816
rect 346766 202872 346822 202881
rect 346766 202807 346822 202816
rect 346780 193254 346808 202807
rect 346584 193248 346636 193254
rect 346584 193190 346636 193196
rect 346768 193248 346820 193254
rect 346768 193190 346820 193196
rect 346596 183569 346624 193190
rect 346582 183560 346638 183569
rect 346582 183495 346638 183504
rect 346766 183560 346822 183569
rect 346766 183495 346822 183504
rect 346780 173942 346808 183495
rect 346584 173936 346636 173942
rect 346584 173878 346636 173884
rect 346768 173936 346820 173942
rect 346768 173878 346820 173884
rect 346596 164218 346624 173878
rect 346584 164212 346636 164218
rect 346584 164154 346636 164160
rect 346768 164212 346820 164218
rect 346768 164154 346820 164160
rect 346780 154601 346808 164154
rect 346582 154592 346638 154601
rect 346582 154527 346638 154536
rect 346766 154592 346822 154601
rect 346766 154527 346822 154536
rect 346596 144906 346624 154527
rect 346584 144900 346636 144906
rect 346584 144842 346636 144848
rect 346768 144900 346820 144906
rect 346768 144842 346820 144848
rect 346780 135289 346808 144842
rect 346582 135280 346638 135289
rect 346582 135215 346638 135224
rect 346766 135280 346822 135289
rect 346766 135215 346822 135224
rect 346596 125594 346624 135215
rect 346584 125588 346636 125594
rect 346584 125530 346636 125536
rect 346584 116000 346636 116006
rect 346584 115942 346636 115948
rect 346596 106282 346624 115942
rect 346584 106276 346636 106282
rect 346584 106218 346636 106224
rect 346584 96688 346636 96694
rect 346584 96630 346636 96636
rect 346596 86970 346624 96630
rect 346584 86964 346636 86970
rect 346584 86906 346636 86912
rect 346492 80776 346544 80782
rect 346492 80718 346544 80724
rect 346504 75970 346532 80718
rect 346504 75942 346624 75970
rect 346596 75886 346624 75942
rect 346492 75880 346544 75886
rect 346492 75822 346544 75828
rect 346584 75880 346636 75886
rect 346584 75822 346636 75828
rect 346504 66314 346532 75822
rect 346504 66286 346624 66314
rect 346596 31822 346624 66286
rect 346584 31816 346636 31822
rect 346584 31758 346636 31764
rect 346492 31748 346544 31754
rect 346492 31690 346544 31696
rect 346504 27606 346532 31690
rect 346492 27600 346544 27606
rect 346492 27542 346544 27548
rect 346492 22772 346544 22778
rect 346492 22714 346544 22720
rect 346504 9654 346532 22714
rect 347688 16720 347740 16726
rect 347686 16688 347688 16697
rect 347740 16688 347742 16697
rect 347686 16623 347742 16632
rect 346492 9648 346544 9654
rect 346492 9590 346544 9596
rect 346492 7268 346544 7274
rect 346492 7210 346544 7216
rect 346400 7132 346452 7138
rect 346400 7074 346452 7080
rect 346504 3398 346532 7210
rect 347792 4894 347820 340054
rect 348252 335594 348280 340190
rect 347976 335566 348280 335594
rect 349264 340054 349370 340082
rect 349632 340054 350014 340082
rect 347976 323626 348004 335566
rect 349160 331832 349212 331838
rect 349160 331774 349212 331780
rect 347976 323598 348096 323626
rect 348068 318782 348096 323598
rect 347964 318776 348016 318782
rect 347964 318718 348016 318724
rect 348056 318776 348108 318782
rect 348056 318718 348108 318724
rect 347976 302326 348004 318718
rect 347964 302320 348016 302326
rect 347964 302262 348016 302268
rect 347964 302184 348016 302190
rect 347964 302126 348016 302132
rect 347976 289814 348004 302126
rect 347964 289808 348016 289814
rect 347964 289750 348016 289756
rect 348056 289740 348108 289746
rect 348056 289682 348108 289688
rect 348068 278866 348096 289682
rect 348056 278860 348108 278866
rect 347976 278798 348004 278829
rect 348056 278802 348108 278808
rect 347964 278792 348016 278798
rect 348016 278740 348096 278746
rect 347964 278734 348096 278740
rect 347976 278718 348096 278734
rect 348068 277409 348096 278718
rect 347870 277400 347926 277409
rect 347870 277335 347926 277344
rect 348054 277400 348110 277409
rect 348054 277335 348110 277344
rect 347884 268818 347912 277335
rect 347884 268790 348096 268818
rect 348068 260914 348096 268790
rect 348056 260908 348108 260914
rect 348056 260850 348108 260856
rect 348148 260840 348200 260846
rect 348148 260782 348200 260788
rect 348160 254658 348188 260782
rect 348148 254652 348200 254658
rect 348148 254594 348200 254600
rect 348056 241528 348108 241534
rect 348056 241470 348108 241476
rect 348068 238746 348096 241470
rect 348056 238740 348108 238746
rect 348056 238682 348108 238688
rect 348056 230376 348108 230382
rect 348056 230318 348108 230324
rect 348068 217410 348096 230318
rect 348068 217382 348188 217410
rect 348160 212566 348188 217382
rect 347964 212560 348016 212566
rect 347964 212502 348016 212508
rect 348148 212560 348200 212566
rect 348148 212502 348200 212508
rect 347976 205698 348004 212502
rect 347964 205692 348016 205698
rect 347964 205634 348016 205640
rect 348056 205556 348108 205562
rect 348056 205498 348108 205504
rect 348068 198098 348096 205498
rect 348068 198070 348188 198098
rect 348160 193254 348188 198070
rect 347964 193248 348016 193254
rect 347962 193216 347964 193225
rect 348148 193248 348200 193254
rect 348016 193216 348018 193225
rect 347962 193151 348018 193160
rect 348146 193216 348148 193225
rect 348200 193216 348202 193225
rect 348146 193151 348202 193160
rect 348160 186266 348188 193151
rect 348068 186238 348188 186266
rect 348068 178786 348096 186238
rect 348068 178758 348188 178786
rect 348160 173942 348188 178758
rect 347964 173936 348016 173942
rect 347964 173878 348016 173884
rect 348148 173936 348200 173942
rect 348148 173878 348200 173884
rect 347976 164218 348004 173878
rect 347964 164212 348016 164218
rect 347964 164154 348016 164160
rect 347964 155780 348016 155786
rect 347964 155722 348016 155728
rect 347976 153202 348004 155722
rect 347964 153196 348016 153202
rect 347964 153138 348016 153144
rect 347964 144832 348016 144838
rect 347964 144774 348016 144780
rect 347976 128194 348004 144774
rect 348424 133748 348476 133754
rect 348424 133690 348476 133696
rect 348436 133657 348464 133690
rect 348422 133648 348478 133657
rect 348422 133583 348478 133592
rect 347976 128166 348096 128194
rect 348068 116113 348096 128166
rect 348054 116104 348110 116113
rect 348054 116039 348110 116048
rect 347962 115968 348018 115977
rect 347962 115903 347964 115912
rect 348016 115903 348018 115912
rect 348056 115932 348108 115938
rect 347964 115874 348016 115880
rect 348056 115874 348108 115880
rect 348068 101402 348096 115874
rect 347976 101374 348096 101402
rect 347976 87145 348004 101374
rect 347962 87136 348018 87145
rect 347962 87071 348018 87080
rect 347870 87000 347926 87009
rect 347870 86935 347926 86944
rect 347884 77382 347912 86935
rect 347872 77376 347924 77382
rect 347872 77318 347924 77324
rect 347872 77240 347924 77246
rect 347872 77182 347924 77188
rect 347884 67658 347912 77182
rect 347872 67652 347924 67658
rect 347872 67594 347924 67600
rect 348056 67652 348108 67658
rect 348056 67594 348108 67600
rect 348068 58002 348096 67594
rect 347964 57996 348016 58002
rect 347964 57938 348016 57944
rect 348056 57996 348108 58002
rect 348056 57938 348108 57944
rect 347976 57882 348004 57938
rect 347976 57854 348096 57882
rect 348068 28966 348096 57854
rect 348056 28960 348108 28966
rect 348056 28902 348108 28908
rect 348148 28960 348200 28966
rect 348148 28902 348200 28908
rect 348160 22778 348188 28902
rect 348148 22772 348200 22778
rect 348148 22714 348200 22720
rect 347872 12436 347924 12442
rect 347872 12378 347924 12384
rect 347884 7614 347912 12378
rect 347872 7608 347924 7614
rect 347872 7550 347924 7556
rect 347964 7336 348016 7342
rect 347964 7278 348016 7284
rect 347780 4888 347832 4894
rect 347780 4830 347832 4836
rect 347872 4888 347924 4894
rect 347872 4830 347924 4836
rect 346676 4140 346728 4146
rect 346676 4082 346728 4088
rect 346492 3392 346544 3398
rect 346492 3334 346544 3340
rect 345480 740 345532 746
rect 345480 682 345532 688
rect 346308 740 346360 746
rect 346308 682 346360 688
rect 345492 480 345520 682
rect 346688 480 346716 4082
rect 347884 480 347912 4830
rect 347976 3330 348004 7278
rect 349068 6860 349120 6866
rect 349068 6802 349120 6808
rect 347964 3324 348016 3330
rect 347964 3266 348016 3272
rect 349080 480 349108 6802
rect 349172 4826 349200 331774
rect 349264 8430 349292 340054
rect 349632 331838 349660 340054
rect 350540 335640 350592 335646
rect 350540 335582 350592 335588
rect 349620 331832 349672 331838
rect 349620 331774 349672 331780
rect 349252 8424 349304 8430
rect 349252 8366 349304 8372
rect 350552 4962 350580 335582
rect 350644 7682 350672 340068
rect 350736 340054 351210 340082
rect 351472 340054 351854 340082
rect 351932 340054 352498 340082
rect 352668 340054 353050 340082
rect 353312 340054 353694 340082
rect 353772 340054 354246 340082
rect 354784 340054 354890 340082
rect 355152 340054 355534 340082
rect 356086 340054 356192 340082
rect 350736 8362 350764 340054
rect 351472 335646 351500 340054
rect 351460 335640 351512 335646
rect 351460 335582 351512 335588
rect 351828 149728 351880 149734
rect 351828 149670 351880 149676
rect 351840 144945 351868 149670
rect 351826 144936 351882 144945
rect 351826 144871 351882 144880
rect 350724 8356 350776 8362
rect 350724 8298 350776 8304
rect 350632 7676 350684 7682
rect 350632 7618 350684 7624
rect 351828 7608 351880 7614
rect 351828 7550 351880 7556
rect 350540 4956 350592 4962
rect 350540 4898 350592 4904
rect 349160 4820 349212 4826
rect 349160 4762 349212 4768
rect 351368 4820 351420 4826
rect 351368 4762 351420 4768
rect 350264 3052 350316 3058
rect 350264 2994 350316 3000
rect 350276 480 350304 2994
rect 351380 480 351408 4762
rect 351840 2990 351868 7550
rect 351932 7070 351960 340054
rect 352668 335628 352696 340054
rect 353208 337204 353260 337210
rect 353208 337146 353260 337152
rect 352116 335600 352696 335628
rect 352116 318866 352144 335600
rect 352024 318838 352144 318866
rect 352024 318782 352052 318838
rect 352012 318776 352064 318782
rect 352012 318718 352064 318724
rect 352104 318708 352156 318714
rect 352104 318650 352156 318656
rect 352116 298110 352144 318650
rect 352104 298104 352156 298110
rect 352104 298046 352156 298052
rect 352196 298036 352248 298042
rect 352196 297978 352248 297984
rect 352208 296698 352236 297978
rect 352116 296670 352236 296698
rect 352116 287094 352144 296670
rect 352012 287088 352064 287094
rect 352012 287030 352064 287036
rect 352104 287088 352156 287094
rect 352104 287030 352156 287036
rect 352024 280226 352052 287030
rect 352012 280220 352064 280226
rect 352012 280162 352064 280168
rect 352104 280152 352156 280158
rect 352104 280094 352156 280100
rect 352116 269113 352144 280094
rect 352102 269104 352158 269113
rect 352102 269039 352158 269048
rect 352286 269104 352342 269113
rect 352286 269039 352342 269048
rect 352300 263498 352328 269039
rect 352012 263492 352064 263498
rect 352012 263434 352064 263440
rect 352288 263492 352340 263498
rect 352288 263434 352340 263440
rect 352024 234666 352052 263434
rect 352012 234660 352064 234666
rect 352012 234602 352064 234608
rect 352196 230376 352248 230382
rect 352196 230318 352248 230324
rect 352208 220862 352236 230318
rect 352012 220856 352064 220862
rect 352012 220798 352064 220804
rect 352196 220856 352248 220862
rect 352196 220798 352248 220804
rect 352024 212566 352052 220798
rect 352012 212560 352064 212566
rect 352012 212502 352064 212508
rect 352104 212560 352156 212566
rect 352104 212502 352156 212508
rect 352116 202910 352144 212502
rect 352012 202904 352064 202910
rect 352010 202872 352012 202881
rect 352104 202904 352156 202910
rect 352064 202872 352066 202881
rect 352104 202846 352156 202852
rect 352010 202807 352066 202816
rect 352102 202736 352158 202745
rect 352102 202671 352158 202680
rect 352116 186454 352144 202671
rect 352104 186448 352156 186454
rect 352104 186390 352156 186396
rect 352012 186312 352064 186318
rect 352012 186254 352064 186260
rect 352024 173942 352052 186254
rect 352012 173936 352064 173942
rect 352012 173878 352064 173884
rect 352104 173936 352156 173942
rect 352104 173878 352156 173884
rect 352116 164257 352144 173878
rect 352102 164248 352158 164257
rect 352102 164183 352158 164192
rect 352010 164112 352066 164121
rect 352010 164047 352066 164056
rect 352024 162858 352052 164047
rect 352012 162852 352064 162858
rect 352012 162794 352064 162800
rect 352012 154556 352064 154562
rect 352012 154498 352064 154504
rect 352024 149734 352052 154498
rect 352012 149728 352064 149734
rect 352012 149670 352064 149676
rect 352010 144936 352066 144945
rect 352010 144871 352012 144880
rect 352064 144871 352066 144880
rect 352196 144900 352248 144906
rect 352012 144842 352064 144848
rect 352196 144842 352248 144848
rect 352208 137714 352236 144842
rect 352116 137686 352236 137714
rect 352116 135250 352144 137686
rect 352104 135244 352156 135250
rect 352104 135186 352156 135192
rect 352196 135244 352248 135250
rect 352196 135186 352248 135192
rect 352208 125633 352236 135186
rect 352010 125624 352066 125633
rect 352010 125559 352012 125568
rect 352064 125559 352066 125568
rect 352194 125624 352250 125633
rect 352194 125559 352196 125568
rect 352012 125530 352064 125536
rect 352248 125559 352250 125568
rect 352196 125530 352248 125536
rect 352208 118402 352236 125530
rect 352116 118374 352236 118402
rect 352116 109154 352144 118374
rect 352116 109126 352236 109154
rect 352208 108882 352236 109126
rect 352024 108854 352236 108882
rect 352024 106282 352052 108854
rect 352012 106276 352064 106282
rect 352012 106218 352064 106224
rect 352196 106276 352248 106282
rect 352196 106218 352248 106224
rect 352208 99090 352236 106218
rect 352116 99062 352236 99090
rect 352116 87145 352144 99062
rect 352102 87136 352158 87145
rect 352102 87071 352158 87080
rect 352010 87000 352066 87009
rect 352010 86935 352012 86944
rect 352064 86935 352066 86944
rect 352012 86906 352064 86912
rect 352104 86896 352156 86902
rect 352104 86838 352156 86844
rect 352116 72434 352144 86838
rect 352024 72406 352144 72434
rect 352024 58138 352052 72406
rect 352012 58132 352064 58138
rect 352012 58074 352064 58080
rect 352012 53848 352064 53854
rect 352012 53790 352064 53796
rect 352024 45558 352052 53790
rect 352012 45552 352064 45558
rect 352012 45494 352064 45500
rect 352380 45552 352432 45558
rect 352380 45494 352432 45500
rect 352392 32314 352420 45494
rect 352116 32286 352420 32314
rect 352116 24290 352144 32286
rect 352116 24262 352236 24290
rect 352208 19378 352236 24262
rect 352012 19372 352064 19378
rect 352012 19314 352064 19320
rect 352196 19372 352248 19378
rect 352196 19314 352248 19320
rect 352024 14074 352052 19314
rect 352012 14068 352064 14074
rect 352012 14010 352064 14016
rect 351920 7064 351972 7070
rect 351920 7006 351972 7012
rect 353220 3738 353248 337146
rect 353312 5030 353340 340054
rect 353772 335628 353800 340054
rect 353496 335600 353800 335628
rect 354680 335640 354732 335646
rect 353496 323626 353524 335600
rect 354680 335582 354732 335588
rect 353496 323598 353616 323626
rect 353588 318782 353616 323598
rect 353484 318776 353536 318782
rect 353484 318718 353536 318724
rect 353576 318776 353628 318782
rect 353576 318718 353628 318724
rect 353496 298110 353524 318718
rect 353484 298104 353536 298110
rect 353484 298046 353536 298052
rect 353576 288448 353628 288454
rect 353576 288390 353628 288396
rect 353588 280158 353616 288390
rect 353576 280152 353628 280158
rect 353576 280094 353628 280100
rect 353668 280152 353720 280158
rect 353668 280094 353720 280100
rect 353680 270314 353708 280094
rect 353680 270286 353800 270314
rect 353772 270042 353800 270286
rect 353680 270014 353800 270042
rect 353680 254658 353708 270014
rect 353668 254652 353720 254658
rect 353668 254594 353720 254600
rect 353576 241528 353628 241534
rect 353576 241470 353628 241476
rect 353588 234734 353616 241470
rect 353576 234728 353628 234734
rect 353576 234670 353628 234676
rect 353576 234592 353628 234598
rect 353576 234534 353628 234540
rect 353588 217410 353616 234534
rect 353588 217382 353708 217410
rect 353680 212566 353708 217382
rect 353484 212560 353536 212566
rect 353484 212502 353536 212508
rect 353668 212560 353720 212566
rect 353668 212502 353720 212508
rect 353496 205698 353524 212502
rect 353484 205692 353536 205698
rect 353484 205634 353536 205640
rect 353576 205624 353628 205630
rect 353576 205566 353628 205572
rect 353588 198098 353616 205566
rect 353588 198070 353708 198098
rect 353680 193254 353708 198070
rect 353484 193248 353536 193254
rect 353482 193216 353484 193225
rect 353668 193248 353720 193254
rect 353536 193216 353538 193225
rect 353482 193151 353538 193160
rect 353666 193216 353668 193225
rect 353720 193216 353722 193225
rect 353666 193151 353722 193160
rect 353680 186266 353708 193151
rect 353588 186238 353708 186266
rect 353588 178786 353616 186238
rect 353588 178758 353708 178786
rect 353680 173942 353708 178758
rect 353484 173936 353536 173942
rect 353482 173904 353484 173913
rect 353668 173936 353720 173942
rect 353536 173904 353538 173913
rect 353668 173878 353720 173884
rect 353482 173839 353538 173848
rect 353574 173768 353630 173777
rect 353574 173703 353630 173712
rect 353588 164218 353616 173703
rect 353484 164212 353536 164218
rect 353484 164154 353536 164160
rect 353576 164212 353628 164218
rect 353576 164154 353628 164160
rect 353496 162858 353524 164154
rect 353484 162852 353536 162858
rect 353484 162794 353536 162800
rect 353484 153264 353536 153270
rect 353484 153206 353536 153212
rect 353496 153134 353524 153206
rect 353484 153128 353536 153134
rect 353484 153070 353536 153076
rect 353484 144832 353536 144838
rect 353484 144774 353536 144780
rect 353496 130370 353524 144774
rect 354588 133748 354640 133754
rect 354588 133690 354640 133696
rect 354600 133657 354628 133690
rect 354586 133648 354642 133657
rect 354586 133583 354642 133592
rect 353496 130342 353708 130370
rect 353680 128330 353708 130342
rect 353588 128302 353708 128330
rect 353588 116006 353616 128302
rect 353576 116000 353628 116006
rect 353576 115942 353628 115948
rect 353576 114572 353628 114578
rect 353576 114514 353628 114520
rect 353588 106282 353616 114514
rect 353484 106276 353536 106282
rect 353484 106218 353536 106224
rect 353576 106276 353628 106282
rect 353576 106218 353628 106224
rect 353496 104854 353524 106218
rect 353484 104848 353536 104854
rect 353484 104790 353536 104796
rect 353484 95260 353536 95266
rect 353484 95202 353536 95208
rect 353496 91746 353524 95202
rect 353496 91718 353616 91746
rect 353588 86970 353616 91718
rect 353484 86964 353536 86970
rect 353484 86906 353536 86912
rect 353576 86964 353628 86970
rect 353576 86906 353628 86912
rect 353496 85542 353524 86906
rect 353484 85536 353536 85542
rect 353484 85478 353536 85484
rect 353576 85468 353628 85474
rect 353576 85410 353628 85416
rect 353588 75886 353616 85410
rect 353576 75880 353628 75886
rect 353576 75822 353628 75828
rect 353668 66292 353720 66298
rect 353668 66234 353720 66240
rect 353680 48362 353708 66234
rect 353588 48334 353708 48362
rect 353588 28966 353616 48334
rect 353576 28960 353628 28966
rect 353576 28902 353628 28908
rect 353668 28960 353720 28966
rect 353668 28902 353720 28908
rect 353680 27606 353708 28902
rect 353668 27600 353720 27606
rect 353668 27542 353720 27548
rect 353668 19304 353720 19310
rect 353668 19246 353720 19252
rect 353680 12186 353708 19246
rect 353404 12158 353708 12186
rect 353404 7002 353432 12158
rect 353392 6996 353444 7002
rect 353392 6938 353444 6944
rect 354692 5098 354720 335582
rect 354784 14482 354812 340054
rect 355152 335646 355180 340054
rect 355140 335640 355192 335646
rect 355140 335582 355192 335588
rect 355966 170232 356022 170241
rect 355966 170167 356022 170176
rect 355980 169561 356008 170167
rect 355966 169552 356022 169561
rect 355966 169487 356022 169496
rect 355966 16960 356022 16969
rect 355966 16895 356022 16904
rect 355980 16726 356008 16895
rect 355968 16720 356020 16726
rect 355968 16662 356020 16668
rect 354772 14476 354824 14482
rect 354772 14418 354824 14424
rect 356164 7750 356192 340054
rect 356256 340054 356730 340082
rect 356256 9926 356284 340054
rect 356808 336734 356836 340190
rect 357452 340054 357926 340082
rect 358280 340054 358570 340082
rect 358832 340054 359214 340082
rect 359292 340054 359766 340082
rect 360304 340054 360410 340082
rect 360672 340054 361054 340082
rect 357348 337136 357400 337142
rect 357348 337078 357400 337084
rect 356796 336728 356848 336734
rect 356796 336670 356848 336676
rect 356520 325712 356572 325718
rect 356520 325654 356572 325660
rect 356532 315994 356560 325654
rect 356520 315988 356572 315994
rect 356520 315930 356572 315936
rect 356612 298172 356664 298178
rect 356612 298114 356664 298120
rect 356624 289898 356652 298114
rect 356440 289870 356652 289898
rect 356440 289814 356468 289870
rect 356428 289808 356480 289814
rect 356428 289750 356480 289756
rect 356520 289740 356572 289746
rect 356520 289682 356572 289688
rect 356532 280158 356560 289682
rect 356428 280152 356480 280158
rect 356428 280094 356480 280100
rect 356520 280152 356572 280158
rect 356520 280094 356572 280100
rect 356440 273358 356468 280094
rect 356428 273352 356480 273358
rect 356428 273294 356480 273300
rect 356428 273216 356480 273222
rect 356428 273158 356480 273164
rect 356440 269090 356468 273158
rect 356440 269062 356560 269090
rect 356532 260914 356560 269062
rect 356520 260908 356572 260914
rect 356520 260850 356572 260856
rect 356428 260772 356480 260778
rect 356428 260714 356480 260720
rect 356440 254046 356468 260714
rect 356428 254040 356480 254046
rect 356428 253982 356480 253988
rect 356428 251116 356480 251122
rect 356428 251058 356480 251064
rect 356440 244322 356468 251058
rect 356428 244316 356480 244322
rect 356428 244258 356480 244264
rect 356520 244180 356572 244186
rect 356520 244122 356572 244128
rect 356532 234734 356560 244122
rect 356520 234728 356572 234734
rect 356520 234670 356572 234676
rect 356428 229220 356480 229226
rect 356428 229162 356480 229168
rect 356440 229090 356468 229162
rect 356428 229084 356480 229090
rect 356428 229026 356480 229032
rect 356428 224936 356480 224942
rect 356428 224878 356480 224884
rect 356440 219450 356468 224878
rect 356440 219422 356560 219450
rect 356532 212634 356560 219422
rect 356520 212628 356572 212634
rect 356520 212570 356572 212576
rect 356428 212560 356480 212566
rect 356428 212502 356480 212508
rect 356440 211138 356468 212502
rect 356428 211132 356480 211138
rect 356428 211074 356480 211080
rect 356428 202836 356480 202842
rect 356428 202778 356480 202784
rect 356440 201498 356468 202778
rect 356440 201470 356560 201498
rect 356532 193322 356560 201470
rect 356520 193316 356572 193322
rect 356520 193258 356572 193264
rect 356428 193248 356480 193254
rect 356480 193196 356560 193202
rect 356428 193190 356560 193196
rect 356440 193174 356560 193190
rect 356532 193066 356560 193174
rect 356532 193038 356652 193066
rect 356624 173942 356652 193038
rect 356428 173936 356480 173942
rect 356426 173904 356428 173913
rect 356612 173936 356664 173942
rect 356480 173904 356482 173913
rect 356612 173878 356664 173884
rect 356426 173839 356482 173848
rect 356518 173768 356574 173777
rect 356518 173703 356574 173712
rect 356532 164218 356560 173703
rect 356428 164212 356480 164218
rect 356428 164154 356480 164160
rect 356520 164212 356572 164218
rect 356520 164154 356572 164160
rect 356440 162858 356468 164154
rect 356428 162852 356480 162858
rect 356428 162794 356480 162800
rect 356428 153264 356480 153270
rect 356428 153206 356480 153212
rect 356440 147694 356468 153206
rect 356428 147688 356480 147694
rect 356428 147630 356480 147636
rect 356520 147484 356572 147490
rect 356520 147426 356572 147432
rect 356532 144906 356560 147426
rect 356520 144900 356572 144906
rect 356520 144842 356572 144848
rect 356612 144900 356664 144906
rect 356612 144842 356664 144848
rect 356624 135289 356652 144842
rect 356426 135280 356482 135289
rect 356426 135215 356428 135224
rect 356480 135215 356482 135224
rect 356610 135280 356666 135289
rect 356610 135215 356666 135224
rect 356428 135186 356480 135192
rect 356520 135176 356572 135182
rect 356520 135118 356572 135124
rect 356532 124234 356560 135118
rect 356428 124228 356480 124234
rect 356428 124170 356480 124176
rect 356520 124228 356572 124234
rect 356520 124170 356572 124176
rect 356440 115938 356468 124170
rect 356428 115932 356480 115938
rect 356428 115874 356480 115880
rect 356612 115932 356664 115938
rect 356612 115874 356664 115880
rect 356624 114510 356652 115874
rect 356612 114504 356664 114510
rect 356612 114446 356664 114452
rect 356428 104984 356480 104990
rect 356428 104926 356480 104932
rect 356440 104854 356468 104926
rect 356428 104848 356480 104854
rect 356428 104790 356480 104796
rect 356612 95260 356664 95266
rect 356612 95202 356664 95208
rect 356624 85610 356652 95202
rect 356428 85604 356480 85610
rect 356428 85546 356480 85552
rect 356612 85604 356664 85610
rect 356612 85546 356664 85552
rect 356440 72570 356468 85546
rect 356440 72542 356652 72570
rect 356624 70258 356652 72542
rect 356532 70230 356652 70258
rect 356532 67590 356560 70230
rect 356520 67584 356572 67590
rect 356520 67526 356572 67532
rect 356428 57996 356480 58002
rect 356428 57938 356480 57944
rect 356440 57882 356468 57938
rect 356440 57854 356560 57882
rect 356532 41562 356560 57854
rect 356532 41534 356652 41562
rect 356624 39386 356652 41534
rect 356532 39358 356652 39386
rect 356532 28966 356560 39358
rect 356428 28960 356480 28966
rect 356428 28902 356480 28908
rect 356520 28960 356572 28966
rect 356520 28902 356572 28908
rect 356244 9920 356296 9926
rect 356244 9862 356296 9868
rect 356152 7744 356204 7750
rect 356152 7686 356204 7692
rect 354956 6044 355008 6050
rect 354956 5986 355008 5992
rect 354680 5092 354732 5098
rect 354680 5034 354732 5040
rect 353300 5024 353352 5030
rect 353300 4966 353352 4972
rect 352564 3732 352616 3738
rect 352564 3674 352616 3680
rect 353208 3732 353260 3738
rect 353208 3674 353260 3680
rect 351828 2984 351880 2990
rect 351828 2926 351880 2932
rect 352576 480 352604 3674
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 353772 480 353800 3334
rect 354968 480 354996 5986
rect 356440 5166 356468 28902
rect 356428 5160 356480 5166
rect 356428 5102 356480 5108
rect 356060 4616 356112 4622
rect 356060 4558 356112 4564
rect 356072 3466 356100 4558
rect 356060 3460 356112 3466
rect 356060 3402 356112 3408
rect 356150 3360 356206 3369
rect 356150 3295 356206 3304
rect 356164 480 356192 3295
rect 357360 480 357388 337078
rect 357452 7818 357480 340054
rect 358280 335646 358308 340054
rect 357624 335640 357676 335646
rect 357624 335582 357676 335588
rect 358268 335640 358320 335646
rect 358268 335582 358320 335588
rect 357636 335306 357664 335582
rect 357624 335300 357676 335306
rect 357624 335242 357676 335248
rect 357624 325848 357676 325854
rect 357624 325790 357676 325796
rect 357636 325689 357664 325790
rect 357622 325680 357678 325689
rect 357622 325615 357678 325624
rect 357806 325680 357862 325689
rect 357806 325615 357862 325624
rect 357544 316062 357572 316093
rect 357820 316062 357848 325615
rect 357532 316056 357584 316062
rect 357808 316056 357860 316062
rect 357584 316004 357664 316010
rect 357532 315998 357664 316004
rect 357808 315998 357860 316004
rect 357544 315982 357664 315998
rect 357636 306406 357664 315982
rect 357532 306400 357584 306406
rect 357532 306342 357584 306348
rect 357624 306400 357676 306406
rect 357624 306342 357676 306348
rect 357544 302954 357572 306342
rect 357544 302926 357756 302954
rect 357728 298353 357756 302926
rect 357714 298344 357770 298353
rect 357714 298279 357770 298288
rect 357622 298208 357678 298217
rect 357622 298143 357678 298152
rect 357636 296721 357664 298143
rect 357622 296712 357678 296721
rect 357622 296647 357678 296656
rect 357806 296712 357862 296721
rect 357806 296647 357862 296656
rect 357820 291922 357848 296647
rect 357624 291916 357676 291922
rect 357624 291858 357676 291864
rect 357808 291916 357860 291922
rect 357808 291858 357860 291864
rect 357636 273358 357664 291858
rect 357624 273352 357676 273358
rect 357624 273294 357676 273300
rect 357624 273216 357676 273222
rect 357624 273158 357676 273164
rect 357636 254046 357664 273158
rect 357624 254040 357676 254046
rect 357624 253982 357676 253988
rect 357624 253904 357676 253910
rect 357624 253846 357676 253852
rect 357636 241482 357664 253846
rect 357636 241454 357756 241482
rect 357728 234666 357756 241454
rect 357716 234660 357768 234666
rect 357716 234602 357768 234608
rect 357624 234592 357676 234598
rect 357624 234534 357676 234540
rect 357636 222170 357664 234534
rect 357636 222142 357756 222170
rect 357728 215354 357756 222142
rect 357716 215348 357768 215354
rect 357716 215290 357768 215296
rect 357624 215280 357676 215286
rect 357624 215222 357676 215228
rect 357636 196058 357664 215222
rect 357544 196030 357664 196058
rect 357544 195922 357572 196030
rect 357544 195894 357664 195922
rect 357636 186454 357664 195894
rect 357624 186448 357676 186454
rect 357624 186390 357676 186396
rect 357544 183598 357572 183629
rect 357532 183592 357584 183598
rect 357584 183540 357664 183546
rect 357532 183534 357664 183540
rect 357544 183518 357664 183534
rect 357636 164218 357664 183518
rect 357624 164212 357676 164218
rect 357624 164154 357676 164160
rect 357624 154624 357676 154630
rect 357624 154566 357676 154572
rect 357636 147642 357664 154566
rect 357636 147614 357756 147642
rect 357728 144974 357756 147614
rect 357624 144968 357676 144974
rect 357544 144916 357624 144922
rect 357544 144910 357676 144916
rect 357716 144968 357768 144974
rect 357716 144910 357768 144916
rect 357544 144894 357664 144910
rect 357544 143546 357572 144894
rect 357532 143540 357584 143546
rect 357532 143482 357584 143488
rect 357624 143540 357676 143546
rect 357624 143482 357676 143488
rect 357636 125594 357664 143482
rect 357624 125588 357676 125594
rect 357624 125530 357676 125536
rect 357716 125588 357768 125594
rect 357716 125530 357768 125536
rect 357728 115977 357756 125530
rect 357714 115968 357770 115977
rect 357714 115903 357770 115912
rect 357806 115832 357862 115841
rect 357806 115767 357862 115776
rect 357820 106321 357848 115767
rect 357622 106312 357678 106321
rect 357622 106247 357678 106256
rect 357806 106312 357862 106321
rect 357806 106247 357862 106256
rect 357636 86970 357664 106247
rect 357624 86964 357676 86970
rect 357624 86906 357676 86912
rect 357808 86964 357860 86970
rect 357808 86906 357860 86912
rect 357820 77353 357848 86906
rect 357622 77344 357678 77353
rect 357622 77279 357678 77288
rect 357806 77344 357862 77353
rect 357806 77279 357862 77288
rect 357636 74526 357664 77279
rect 357624 74520 357676 74526
rect 357624 74462 357676 74468
rect 357532 64932 357584 64938
rect 357532 64874 357584 64880
rect 357544 46866 357572 64874
rect 357544 46838 357664 46866
rect 357636 33810 357664 46838
rect 357544 33782 357664 33810
rect 357544 19378 357572 33782
rect 357532 19372 357584 19378
rect 357532 19314 357584 19320
rect 357624 19372 357676 19378
rect 357624 19314 357676 19320
rect 357636 9858 357664 19314
rect 357624 9852 357676 9858
rect 357624 9794 357676 9800
rect 357440 7812 357492 7818
rect 357440 7754 357492 7760
rect 358832 5234 358860 340054
rect 359292 331906 359320 340054
rect 360108 337068 360160 337074
rect 360108 337010 360160 337016
rect 359096 331900 359148 331906
rect 359096 331842 359148 331848
rect 359280 331900 359332 331906
rect 359280 331842 359332 331848
rect 359108 321638 359136 331842
rect 359096 321632 359148 321638
rect 359096 321574 359148 321580
rect 359004 318844 359056 318850
rect 359004 318786 359056 318792
rect 359016 318730 359044 318786
rect 359016 318702 359136 318730
rect 359108 292618 359136 318702
rect 359016 292590 359136 292618
rect 359016 285002 359044 292590
rect 358924 284974 359044 285002
rect 358924 282826 358952 284974
rect 358924 282798 359136 282826
rect 359108 280158 359136 282798
rect 359004 280152 359056 280158
rect 359004 280094 359056 280100
rect 359096 280152 359148 280158
rect 359096 280094 359148 280100
rect 359016 270745 359044 280094
rect 359002 270736 359058 270745
rect 359002 270671 359058 270680
rect 358910 270464 358966 270473
rect 358910 270399 358966 270408
rect 358924 263566 358952 270399
rect 358912 263560 358964 263566
rect 358912 263502 358964 263508
rect 359096 263492 359148 263498
rect 359096 263434 359148 263440
rect 359108 260846 359136 263434
rect 359096 260840 359148 260846
rect 359096 260782 359148 260788
rect 359004 251320 359056 251326
rect 359004 251262 359056 251268
rect 359016 251190 359044 251262
rect 359004 251184 359056 251190
rect 359004 251126 359056 251132
rect 359004 244180 359056 244186
rect 359004 244122 359056 244128
rect 359016 232014 359044 244122
rect 359004 232008 359056 232014
rect 359004 231950 359056 231956
rect 359096 231872 359148 231878
rect 359096 231814 359148 231820
rect 359108 226930 359136 231814
rect 359016 226902 359136 226930
rect 359016 212634 359044 226902
rect 359004 212628 359056 212634
rect 359004 212570 359056 212576
rect 358912 208412 358964 208418
rect 358912 208354 358964 208360
rect 358924 200161 358952 208354
rect 358910 200152 358966 200161
rect 358910 200087 358966 200096
rect 359094 200152 359150 200161
rect 359094 200087 359150 200096
rect 359108 196042 359136 200087
rect 358912 196036 358964 196042
rect 358912 195978 358964 195984
rect 359096 196036 359148 196042
rect 359096 195978 359148 195984
rect 358924 190505 358952 195978
rect 358910 190496 358966 190505
rect 358910 190431 358966 190440
rect 359186 190496 359242 190505
rect 359186 190431 359242 190440
rect 359200 189802 359228 190431
rect 359108 189774 359228 189802
rect 359108 178838 359136 189774
rect 359096 178832 359148 178838
rect 359096 178774 359148 178780
rect 359004 178764 359056 178770
rect 359004 178706 359056 178712
rect 359016 167074 359044 178706
rect 359004 167068 359056 167074
rect 359004 167010 359056 167016
rect 359096 166932 359148 166938
rect 359096 166874 359148 166880
rect 359108 157350 359136 166874
rect 359096 157344 359148 157350
rect 359096 157286 359148 157292
rect 359004 154624 359056 154630
rect 359004 154566 359056 154572
rect 359016 147762 359044 154566
rect 359004 147756 359056 147762
rect 359004 147698 359056 147704
rect 359004 147620 359056 147626
rect 359004 147562 359056 147568
rect 359016 135386 359044 147562
rect 359004 135380 359056 135386
rect 359004 135322 359056 135328
rect 359004 135244 359056 135250
rect 359004 135186 359056 135192
rect 359016 133906 359044 135186
rect 359016 133878 359136 133906
rect 359108 115954 359136 133878
rect 359016 115926 359136 115954
rect 359016 106298 359044 115926
rect 359016 106270 359136 106298
rect 359108 96642 359136 106270
rect 359016 96614 359136 96642
rect 359016 84402 359044 96614
rect 359016 84374 359136 84402
rect 359108 84266 359136 84374
rect 359016 84238 359136 84266
rect 359016 82822 359044 84238
rect 359004 82816 359056 82822
rect 359004 82758 359056 82764
rect 359004 73228 359056 73234
rect 359004 73170 359056 73176
rect 359016 70394 359044 73170
rect 358924 70366 359044 70394
rect 358924 64954 358952 70366
rect 358924 64926 359136 64954
rect 359108 63510 359136 64926
rect 359096 63504 359148 63510
rect 359096 63446 359148 63452
rect 359188 53848 359240 53854
rect 359188 53790 359240 53796
rect 359200 46918 359228 53790
rect 359004 46912 359056 46918
rect 359004 46854 359056 46860
rect 359188 46912 359240 46918
rect 359188 46854 359240 46860
rect 359016 45558 359044 46854
rect 359004 45552 359056 45558
rect 359004 45494 359056 45500
rect 359004 35964 359056 35970
rect 359004 35906 359056 35912
rect 359016 27606 359044 35906
rect 359004 27600 359056 27606
rect 359004 27542 359056 27548
rect 359004 18012 359056 18018
rect 359004 17954 359056 17960
rect 359016 12458 359044 17954
rect 359016 12430 359136 12458
rect 359108 12322 359136 12430
rect 358924 12294 359136 12322
rect 358924 9602 358952 12294
rect 358924 9574 359044 9602
rect 359016 7886 359044 9574
rect 359004 7880 359056 7886
rect 359004 7822 359056 7828
rect 358820 5228 358872 5234
rect 358820 5170 358872 5176
rect 358544 4956 358596 4962
rect 358544 4898 358596 4904
rect 358556 480 358584 4898
rect 360120 626 360148 337010
rect 360200 335640 360252 335646
rect 360200 335582 360252 335588
rect 360212 5914 360240 335582
rect 360304 9790 360332 340054
rect 360672 335646 360700 340054
rect 360660 335640 360712 335646
rect 360660 335582 360712 335588
rect 360292 9784 360344 9790
rect 360292 9726 360344 9732
rect 361592 7954 361620 340068
rect 361776 340054 362250 340082
rect 362512 340054 362894 340082
rect 363064 340054 363446 340082
rect 363800 340054 364090 340082
rect 364352 340054 364734 340082
rect 364996 340054 365286 340082
rect 361672 335640 361724 335646
rect 361672 335582 361724 335588
rect 361684 9314 361712 335582
rect 361776 9722 361804 340054
rect 362512 335646 362540 340054
rect 362500 335640 362552 335646
rect 362500 335582 362552 335588
rect 362960 334416 363012 334422
rect 362960 334358 363012 334364
rect 361764 9716 361816 9722
rect 361764 9658 361816 9664
rect 361672 9308 361724 9314
rect 361672 9250 361724 9256
rect 361580 7948 361632 7954
rect 361580 7890 361632 7896
rect 360200 5908 360252 5914
rect 360200 5850 360252 5856
rect 362132 5908 362184 5914
rect 362132 5850 362184 5856
rect 360936 2984 360988 2990
rect 360936 2926 360988 2932
rect 359752 598 360148 626
rect 359752 480 359780 598
rect 360948 480 360976 2926
rect 362144 480 362172 5850
rect 362972 4622 363000 334358
rect 363064 8022 363092 340054
rect 363696 336932 363748 336938
rect 363696 336874 363748 336880
rect 363604 336796 363656 336802
rect 363604 336738 363656 336744
rect 363052 8016 363104 8022
rect 363052 7958 363104 7964
rect 362960 4616 363012 4622
rect 362960 4558 363012 4564
rect 363616 4010 363644 336738
rect 363604 4004 363656 4010
rect 363604 3946 363656 3952
rect 363708 3262 363736 336874
rect 363800 334422 363828 340054
rect 363788 334416 363840 334422
rect 363788 334358 363840 334364
rect 364248 260840 364300 260846
rect 364248 260782 364300 260788
rect 364260 251297 364288 260782
rect 364246 251288 364302 251297
rect 364246 251223 364302 251232
rect 364246 251152 364302 251161
rect 364246 251087 364302 251096
rect 364260 242214 364288 251087
rect 364248 242208 364300 242214
rect 364248 242150 364300 242156
rect 364246 40488 364302 40497
rect 364246 40423 364302 40432
rect 364260 40225 364288 40423
rect 364246 40216 364302 40225
rect 364246 40151 364302 40160
rect 364352 5846 364380 340054
rect 364996 331430 365024 340054
rect 365916 337686 365944 340068
rect 365904 337680 365956 337686
rect 365904 337622 365956 337628
rect 365810 337512 365866 337521
rect 365810 337447 365866 337456
rect 365720 337340 365772 337346
rect 365720 337282 365772 337288
rect 365732 337226 365760 337282
rect 365824 337226 365852 337447
rect 365732 337198 365852 337226
rect 364524 331424 364576 331430
rect 364524 331366 364576 331372
rect 364984 331424 365036 331430
rect 364984 331366 365036 331372
rect 364536 331106 364564 331366
rect 366008 331242 366036 340190
rect 366916 337680 366968 337686
rect 366916 337622 366968 337628
rect 366364 337000 366416 337006
rect 366364 336942 366416 336948
rect 365916 331214 366036 331242
rect 364536 331078 364656 331106
rect 364628 321314 364656 331078
rect 364536 321286 364656 321314
rect 364536 318730 364564 321286
rect 364536 318702 364656 318730
rect 364628 292618 364656 318702
rect 365916 317506 365944 331214
rect 365824 317478 365944 317506
rect 365824 316033 365852 317478
rect 365810 316024 365866 316033
rect 365810 315959 365866 315968
rect 365994 316024 366050 316033
rect 365994 315959 366050 315968
rect 366008 306406 366036 315959
rect 365812 306400 365864 306406
rect 365812 306342 365864 306348
rect 365996 306400 366048 306406
rect 365996 306342 366048 306348
rect 365824 299418 365852 306342
rect 365824 299390 365944 299418
rect 365916 298110 365944 299390
rect 365904 298104 365956 298110
rect 365904 298046 365956 298052
rect 365904 297968 365956 297974
rect 365904 297910 365956 297916
rect 364536 292590 364656 292618
rect 364536 282946 364564 292590
rect 364524 282940 364576 282946
rect 364524 282882 364576 282888
rect 364616 282804 364668 282810
rect 364616 282746 364668 282752
rect 364628 280158 364656 282746
rect 364616 280152 364668 280158
rect 364616 280094 364668 280100
rect 364524 273216 364576 273222
rect 364524 273158 364576 273164
rect 364536 263634 364564 273158
rect 364524 263628 364576 263634
rect 364524 263570 364576 263576
rect 364616 263492 364668 263498
rect 364616 263434 364668 263440
rect 364628 260846 364656 263434
rect 364616 260840 364668 260846
rect 364616 260782 364668 260788
rect 364616 242208 364668 242214
rect 364616 242150 364668 242156
rect 364628 235958 364656 242150
rect 364616 235952 364668 235958
rect 364616 235894 364668 235900
rect 364432 218068 364484 218074
rect 364432 218010 364484 218016
rect 364444 217977 364472 218010
rect 364430 217968 364486 217977
rect 364430 217903 364486 217912
rect 364614 217968 364670 217977
rect 364614 217903 364670 217912
rect 364628 212378 364656 217903
rect 364444 212350 364656 212378
rect 364444 200161 364472 212350
rect 364430 200152 364486 200161
rect 364430 200087 364486 200096
rect 364614 200152 364670 200161
rect 364614 200087 364670 200096
rect 364628 196110 364656 200087
rect 364616 196104 364668 196110
rect 365916 196058 365944 297910
rect 364616 196046 364668 196052
rect 365824 196030 365944 196058
rect 364616 195968 364668 195974
rect 364616 195910 364668 195916
rect 365824 195922 365852 196030
rect 364628 190505 364656 195910
rect 365824 195894 365944 195922
rect 364614 190496 364670 190505
rect 364614 190431 364670 190440
rect 364798 190496 364854 190505
rect 364798 190431 364854 190440
rect 364812 183410 364840 190431
rect 364720 183382 364840 183410
rect 364720 172553 364748 183382
rect 364522 172544 364578 172553
rect 364522 172479 364578 172488
rect 364706 172544 364762 172553
rect 364706 172479 364762 172488
rect 364536 167686 364564 172479
rect 364524 167680 364576 167686
rect 364524 167622 364576 167628
rect 364616 154624 364668 154630
rect 364536 154572 364616 154578
rect 364536 154566 364668 154572
rect 364536 154550 364656 154566
rect 364536 151994 364564 154550
rect 364536 151966 364748 151994
rect 364720 147506 364748 151966
rect 364628 147478 364748 147506
rect 364628 144906 364656 147478
rect 364616 144900 364668 144906
rect 364616 144842 364668 144848
rect 364708 144900 364760 144906
rect 364708 144842 364760 144848
rect 364720 135289 364748 144842
rect 364522 135280 364578 135289
rect 364522 135215 364578 135224
rect 364706 135280 364762 135289
rect 364706 135215 364762 135224
rect 364536 130370 364564 135215
rect 364536 130342 364656 130370
rect 364628 125594 364656 130342
rect 364616 125588 364668 125594
rect 364616 125530 364668 125536
rect 364524 116000 364576 116006
rect 364524 115942 364576 115948
rect 364536 111058 364564 115942
rect 364444 111030 364564 111058
rect 364444 108882 364472 111030
rect 364444 108854 364656 108882
rect 364628 106282 364656 108854
rect 364524 106276 364576 106282
rect 364524 106218 364576 106224
rect 364616 106276 364668 106282
rect 364616 106218 364668 106224
rect 364536 86902 364564 106218
rect 364524 86896 364576 86902
rect 364524 86838 364576 86844
rect 364524 77308 364576 77314
rect 364524 77250 364576 77256
rect 364536 22166 364564 77250
rect 365916 60738 365944 195894
rect 365824 60710 365944 60738
rect 365824 60602 365852 60710
rect 365824 60574 365944 60602
rect 365916 41426 365944 60574
rect 365824 41398 365944 41426
rect 365824 41290 365852 41398
rect 365824 41262 365944 41290
rect 364524 22160 364576 22166
rect 364524 22102 364576 22108
rect 364524 22024 364576 22030
rect 364524 21966 364576 21972
rect 364536 8090 364564 21966
rect 365916 19394 365944 41262
rect 365824 19366 365944 19394
rect 365824 12594 365852 19366
rect 365640 12566 365852 12594
rect 365640 10538 365668 12566
rect 365628 10532 365680 10538
rect 365628 10474 365680 10480
rect 364524 8084 364576 8090
rect 364524 8026 364576 8032
rect 364340 5840 364392 5846
rect 364340 5782 364392 5788
rect 365720 5024 365772 5030
rect 365720 4966 365772 4972
rect 364524 4004 364576 4010
rect 364524 3946 364576 3952
rect 363696 3256 363748 3262
rect 363696 3198 363748 3204
rect 363328 3120 363380 3126
rect 363328 3062 363380 3068
rect 363340 480 363368 3062
rect 364536 480 364564 3946
rect 365732 480 365760 4966
rect 366376 4010 366404 336942
rect 366456 336864 366508 336870
rect 366456 336806 366508 336812
rect 366364 4004 366416 4010
rect 366364 3946 366416 3952
rect 366468 3330 366496 336806
rect 366456 3324 366508 3330
rect 366456 3266 366508 3272
rect 366928 480 366956 337622
rect 367006 170232 367062 170241
rect 367006 170167 367062 170176
rect 367020 169833 367048 170167
rect 367006 169824 367062 169833
rect 367006 169759 367062 169768
rect 367112 8158 367140 340068
rect 367296 340054 367770 340082
rect 368032 340054 368414 340082
rect 368584 340054 368966 340082
rect 367192 335640 367244 335646
rect 367192 335582 367244 335588
rect 367204 10674 367232 335582
rect 367192 10668 367244 10674
rect 367192 10610 367244 10616
rect 367296 10606 367324 340054
rect 368032 335646 368060 340054
rect 368020 335640 368072 335646
rect 368020 335582 368072 335588
rect 367284 10600 367336 10606
rect 367284 10542 367336 10548
rect 368584 8226 368612 340054
rect 369596 337482 369624 340068
rect 369872 340054 370254 340082
rect 370516 340054 370806 340082
rect 369584 337476 369636 337482
rect 369584 337418 369636 337424
rect 369768 191820 369820 191826
rect 369768 191762 369820 191768
rect 369780 182209 369808 191762
rect 369766 182200 369822 182209
rect 369766 182135 369822 182144
rect 368572 8220 368624 8226
rect 368572 8162 368624 8168
rect 367100 8152 367152 8158
rect 367100 8094 367152 8100
rect 369872 5982 369900 340054
rect 370516 336734 370544 340054
rect 371436 337414 371464 340068
rect 371620 340054 372002 340082
rect 372646 340054 372752 340082
rect 371424 337408 371476 337414
rect 371424 337350 371476 337356
rect 370504 336728 370556 336734
rect 370504 336670 370556 336676
rect 371620 331242 371648 340054
rect 372528 337408 372580 337414
rect 372528 337350 372580 337356
rect 371436 331214 371648 331242
rect 370044 327140 370096 327146
rect 370044 327082 370096 327088
rect 370056 317506 370084 327082
rect 371436 321722 371464 331214
rect 371436 321694 371556 321722
rect 371528 318866 371556 321694
rect 371436 318838 371556 318866
rect 371436 318782 371464 318838
rect 371424 318776 371476 318782
rect 371424 318718 371476 318724
rect 370056 317478 370268 317506
rect 370240 299538 370268 317478
rect 371332 309324 371384 309330
rect 371332 309266 371384 309272
rect 371344 307578 371372 309266
rect 371252 307550 371372 307578
rect 370136 299532 370188 299538
rect 370136 299474 370188 299480
rect 370228 299532 370280 299538
rect 370228 299474 370280 299480
rect 370148 298110 370176 299474
rect 371252 298178 371280 307550
rect 371240 298172 371292 298178
rect 371240 298114 371292 298120
rect 371608 298172 371660 298178
rect 371608 298114 371660 298120
rect 370136 298104 370188 298110
rect 370136 298046 370188 298052
rect 371620 292618 371648 298114
rect 371436 292590 371648 292618
rect 370228 289740 370280 289746
rect 370228 289682 370280 289688
rect 370240 280158 370268 289682
rect 371436 280158 371464 292590
rect 369952 280152 370004 280158
rect 369952 280094 370004 280100
rect 370228 280152 370280 280158
rect 370228 280094 370280 280100
rect 371424 280152 371476 280158
rect 371424 280094 371476 280100
rect 369964 278769 369992 280094
rect 369950 278760 370006 278769
rect 369950 278695 370006 278704
rect 370318 278760 370374 278769
rect 370318 278695 370374 278704
rect 370332 253858 370360 278695
rect 371424 270564 371476 270570
rect 371424 270506 371476 270512
rect 371436 260846 371464 270506
rect 371424 260840 371476 260846
rect 371424 260782 371476 260788
rect 370056 253830 370360 253858
rect 370056 251190 370084 253830
rect 371424 251252 371476 251258
rect 371424 251194 371476 251200
rect 370044 251184 370096 251190
rect 370044 251126 370096 251132
rect 369952 241528 370004 241534
rect 369952 241470 370004 241476
rect 369964 231878 369992 241470
rect 371436 234598 371464 251194
rect 371424 234592 371476 234598
rect 371424 234534 371476 234540
rect 371424 234456 371476 234462
rect 371424 234398 371476 234404
rect 369952 231872 370004 231878
rect 369952 231814 370004 231820
rect 370044 231872 370096 231878
rect 370044 231814 370096 231820
rect 370056 215422 370084 231814
rect 370044 215416 370096 215422
rect 370044 215358 370096 215364
rect 371436 215286 371464 234398
rect 370044 215280 370096 215286
rect 370044 215222 370096 215228
rect 371424 215280 371476 215286
rect 371424 215222 371476 215228
rect 370056 211138 370084 215222
rect 371424 215144 371476 215150
rect 371424 215086 371476 215092
rect 370044 211132 370096 211138
rect 370044 211074 370096 211080
rect 370228 211132 370280 211138
rect 370228 211074 370280 211080
rect 370240 201521 370268 211074
rect 370042 201512 370098 201521
rect 370042 201447 370098 201456
rect 370226 201512 370282 201521
rect 370226 201447 370282 201456
rect 370056 196110 370084 201447
rect 370044 196104 370096 196110
rect 370044 196046 370096 196052
rect 371436 195974 371464 215086
rect 370044 195968 370096 195974
rect 370044 195910 370096 195916
rect 371424 195968 371476 195974
rect 371424 195910 371476 195916
rect 370056 191826 370084 195910
rect 371424 195832 371476 195838
rect 371424 195774 371476 195780
rect 370044 191820 370096 191826
rect 370044 191762 370096 191768
rect 369950 182200 370006 182209
rect 369950 182135 369952 182144
rect 370004 182135 370006 182144
rect 370412 182164 370464 182170
rect 369952 182106 370004 182112
rect 370412 182106 370464 182112
rect 370424 172553 370452 182106
rect 371436 176662 371464 195774
rect 371424 176656 371476 176662
rect 371424 176598 371476 176604
rect 371424 176520 371476 176526
rect 371424 176462 371476 176468
rect 370226 172544 370282 172553
rect 370226 172479 370282 172488
rect 370410 172544 370466 172553
rect 370410 172479 370466 172488
rect 370240 164257 370268 172479
rect 370042 164248 370098 164257
rect 370042 164183 370098 164192
rect 370226 164248 370282 164257
rect 370226 164183 370282 164192
rect 370056 157593 370084 164183
rect 370042 157584 370098 157593
rect 370042 157519 370098 157528
rect 371436 157350 371464 176462
rect 371882 170096 371938 170105
rect 371882 170031 371938 170040
rect 371896 169833 371924 170031
rect 371882 169824 371938 169833
rect 371882 169759 371938 169768
rect 371424 157344 371476 157350
rect 371424 157286 371476 157292
rect 371424 157208 371476 157214
rect 371424 157150 371476 157156
rect 370042 154592 370098 154601
rect 370042 154527 370044 154536
rect 370096 154527 370098 154536
rect 370044 154498 370096 154504
rect 370044 147620 370096 147626
rect 370044 147562 370096 147568
rect 370056 144922 370084 147562
rect 370056 144894 370176 144922
rect 370148 138281 370176 144894
rect 370134 138272 370190 138281
rect 370134 138207 370190 138216
rect 370042 135280 370098 135289
rect 370042 135215 370044 135224
rect 370096 135215 370098 135224
rect 370044 135186 370096 135192
rect 370044 128308 370096 128314
rect 370044 128250 370096 128256
rect 370056 125610 370084 128250
rect 370056 125582 370176 125610
rect 370148 120766 370176 125582
rect 370136 120760 370188 120766
rect 370136 120702 370188 120708
rect 370136 120624 370188 120630
rect 370136 120566 370188 120572
rect 370148 109070 370176 120566
rect 370136 109064 370188 109070
rect 370136 109006 370188 109012
rect 370136 106344 370188 106350
rect 370136 106286 370188 106292
rect 370148 101402 370176 106286
rect 370148 101374 370268 101402
rect 370240 96665 370268 101374
rect 370042 96656 370098 96665
rect 370042 96591 370098 96600
rect 370226 96656 370282 96665
rect 370226 96591 370282 96600
rect 370056 86902 370084 96591
rect 370044 86896 370096 86902
rect 370044 86838 370096 86844
rect 371436 80102 371464 157150
rect 371424 80096 371476 80102
rect 371424 80038 371476 80044
rect 371424 79960 371476 79966
rect 371424 79902 371476 79908
rect 370044 77308 370096 77314
rect 370044 77250 370096 77256
rect 370056 61130 370084 77250
rect 370044 61124 370096 61130
rect 370044 61066 370096 61072
rect 371436 60654 371464 79902
rect 371424 60648 371476 60654
rect 371424 60590 371476 60596
rect 371424 56704 371476 56710
rect 371424 56646 371476 56652
rect 371436 56574 371464 56646
rect 371424 56568 371476 56574
rect 371424 56510 371476 56516
rect 370136 48340 370188 48346
rect 370136 48282 370188 48288
rect 370148 41478 370176 48282
rect 371332 47048 371384 47054
rect 371332 46990 371384 46996
rect 371344 46918 371372 46990
rect 371332 46912 371384 46918
rect 371332 46854 371384 46860
rect 371516 46844 371568 46850
rect 371516 46786 371568 46792
rect 370136 41472 370188 41478
rect 370136 41414 370188 41420
rect 369952 38616 370004 38622
rect 369952 38558 370004 38564
rect 369964 33862 369992 38558
rect 369952 33856 370004 33862
rect 369952 33798 370004 33804
rect 370228 33856 370280 33862
rect 370228 33798 370280 33804
rect 370240 19378 370268 33798
rect 371528 19378 371556 46786
rect 370044 19372 370096 19378
rect 370044 19314 370096 19320
rect 370228 19372 370280 19378
rect 370228 19314 370280 19320
rect 371332 19372 371384 19378
rect 371332 19314 371384 19320
rect 371516 19372 371568 19378
rect 371516 19314 371568 19320
rect 370056 9602 370084 19314
rect 370502 16824 370558 16833
rect 370502 16759 370558 16768
rect 370516 16425 370544 16759
rect 370502 16416 370558 16425
rect 370502 16351 370558 16360
rect 370056 9574 370176 9602
rect 370148 8294 370176 9574
rect 370136 8288 370188 8294
rect 370136 8230 370188 8236
rect 371344 6118 371372 19314
rect 371332 6112 371384 6118
rect 371332 6054 371384 6060
rect 369860 5976 369912 5982
rect 369860 5918 369912 5924
rect 369216 5840 369268 5846
rect 369216 5782 369268 5788
rect 368020 3460 368072 3466
rect 368020 3402 368072 3408
rect 368032 480 368060 3402
rect 369228 480 369256 5782
rect 372540 4010 372568 337350
rect 372724 7546 372752 340054
rect 373276 337754 373304 340068
rect 373264 337748 373316 337754
rect 373264 337690 373316 337696
rect 373368 331242 373396 340190
rect 372816 331214 373396 331242
rect 374104 340054 374486 340082
rect 372712 7540 372764 7546
rect 372712 7482 372764 7488
rect 372816 6186 372844 331214
rect 373906 40624 373962 40633
rect 373906 40559 373962 40568
rect 373920 40225 373948 40559
rect 373906 40216 373962 40225
rect 373906 40151 373962 40160
rect 374104 7478 374132 340054
rect 375116 337822 375144 340068
rect 375392 340054 375682 340082
rect 375104 337816 375156 337822
rect 375104 337758 375156 337764
rect 375288 337816 375340 337822
rect 375288 337758 375340 337764
rect 374644 336796 374696 336802
rect 374644 336738 374696 336744
rect 374092 7472 374144 7478
rect 374092 7414 374144 7420
rect 372804 6180 372856 6186
rect 372804 6122 372856 6128
rect 372896 6180 372948 6186
rect 372896 6122 372948 6128
rect 372908 4434 372936 6122
rect 372816 4406 372936 4434
rect 371608 4004 371660 4010
rect 371608 3946 371660 3952
rect 372528 4004 372580 4010
rect 372528 3946 372580 3952
rect 370412 3256 370464 3262
rect 370412 3198 370464 3204
rect 370424 480 370452 3198
rect 371620 480 371648 3946
rect 372816 480 372844 4406
rect 374656 3126 374684 336738
rect 375196 164212 375248 164218
rect 375196 164154 375248 164160
rect 375208 154601 375236 164154
rect 375194 154592 375250 154601
rect 375194 154527 375250 154536
rect 374644 3120 374696 3126
rect 374644 3062 374696 3068
rect 375196 3120 375248 3126
rect 375196 3062 375248 3068
rect 374000 3052 374052 3058
rect 374000 2994 374052 3000
rect 374012 480 374040 2994
rect 375208 480 375236 3062
rect 375300 3058 375328 337758
rect 375392 6254 375420 340054
rect 375760 336734 375788 340190
rect 376024 337748 376076 337754
rect 376024 337690 376076 337696
rect 375748 336728 375800 336734
rect 375748 336670 375800 336676
rect 375564 327140 375616 327146
rect 375564 327082 375616 327088
rect 375576 318782 375604 327082
rect 375564 318776 375616 318782
rect 375564 318718 375616 318724
rect 375748 318776 375800 318782
rect 375748 318718 375800 318724
rect 375760 317422 375788 318718
rect 375748 317416 375800 317422
rect 375748 317358 375800 317364
rect 375748 309120 375800 309126
rect 375748 309062 375800 309068
rect 375760 299538 375788 309062
rect 375656 299532 375708 299538
rect 375656 299474 375708 299480
rect 375748 299532 375800 299538
rect 375748 299474 375800 299480
rect 375668 292618 375696 299474
rect 375576 292590 375696 292618
rect 375576 289814 375604 292590
rect 375564 289808 375616 289814
rect 375564 289750 375616 289756
rect 375748 289808 375800 289814
rect 375748 289750 375800 289756
rect 375760 280158 375788 289750
rect 375472 280152 375524 280158
rect 375472 280094 375524 280100
rect 375748 280152 375800 280158
rect 375748 280094 375800 280100
rect 375484 278730 375512 280094
rect 375472 278724 375524 278730
rect 375472 278666 375524 278672
rect 375656 263492 375708 263498
rect 375656 263434 375708 263440
rect 375668 260846 375696 263434
rect 375656 260840 375708 260846
rect 375656 260782 375708 260788
rect 375564 251252 375616 251258
rect 375564 251194 375616 251200
rect 375576 251161 375604 251194
rect 375562 251152 375618 251161
rect 375562 251087 375618 251096
rect 375746 251152 375802 251161
rect 375746 251087 375802 251096
rect 375760 241534 375788 251087
rect 375748 241528 375800 241534
rect 375748 241470 375800 241476
rect 375840 241528 375892 241534
rect 375840 241470 375892 241476
rect 375852 231878 375880 241470
rect 375564 231872 375616 231878
rect 375562 231840 375564 231849
rect 375840 231872 375892 231878
rect 375616 231840 375618 231849
rect 375562 231775 375618 231784
rect 375838 231840 375840 231849
rect 375892 231840 375894 231849
rect 375838 231775 375894 231784
rect 375852 212566 375880 231775
rect 375564 212560 375616 212566
rect 375562 212528 375564 212537
rect 375840 212560 375892 212566
rect 375616 212528 375618 212537
rect 375562 212463 375618 212472
rect 375838 212528 375840 212537
rect 375892 212528 375894 212537
rect 375838 212463 375894 212472
rect 375852 201482 375880 212463
rect 375564 201476 375616 201482
rect 375564 201418 375616 201424
rect 375840 201476 375892 201482
rect 375840 201418 375892 201424
rect 375576 192001 375604 201418
rect 375562 191992 375618 192001
rect 375562 191927 375618 191936
rect 375562 191856 375618 191865
rect 375472 191820 375524 191826
rect 375562 191791 375564 191800
rect 375472 191762 375524 191768
rect 375616 191791 375618 191800
rect 375564 191762 375616 191768
rect 375484 182209 375512 191762
rect 375470 182200 375526 182209
rect 375470 182135 375526 182144
rect 375746 182200 375802 182209
rect 375746 182135 375802 182144
rect 375760 172553 375788 182135
rect 375562 172544 375618 172553
rect 375562 172479 375618 172488
rect 375746 172544 375802 172553
rect 375746 172479 375802 172488
rect 375576 164218 375604 172479
rect 375564 164212 375616 164218
rect 375564 164154 375616 164160
rect 375562 154592 375618 154601
rect 375562 154527 375564 154536
rect 375616 154527 375618 154536
rect 375748 154556 375800 154562
rect 375564 154498 375616 154504
rect 375748 154498 375800 154504
rect 375760 135425 375788 154498
rect 375746 135416 375802 135425
rect 375746 135351 375802 135360
rect 375562 135280 375618 135289
rect 375562 135215 375564 135224
rect 375616 135215 375618 135224
rect 375564 135186 375616 135192
rect 375748 135176 375800 135182
rect 375748 135118 375800 135124
rect 375760 120766 375788 135118
rect 375472 120760 375524 120766
rect 375472 120702 375524 120708
rect 375748 120760 375800 120766
rect 375748 120702 375800 120708
rect 375484 115938 375512 120702
rect 375472 115932 375524 115938
rect 375472 115874 375524 115880
rect 375748 115932 375800 115938
rect 375748 115874 375800 115880
rect 375760 96801 375788 115874
rect 375746 96792 375802 96801
rect 375746 96727 375802 96736
rect 375562 96656 375618 96665
rect 375562 96591 375618 96600
rect 375576 61130 375604 96591
rect 375564 61124 375616 61130
rect 375564 61066 375616 61072
rect 375656 48340 375708 48346
rect 375656 48282 375708 48288
rect 375668 41614 375696 48282
rect 375656 41608 375708 41614
rect 375656 41550 375708 41556
rect 375472 37324 375524 37330
rect 375472 37266 375524 37272
rect 375484 33810 375512 37266
rect 375484 33782 375788 33810
rect 375760 19378 375788 33782
rect 375564 19372 375616 19378
rect 375564 19314 375616 19320
rect 375748 19372 375800 19378
rect 375748 19314 375800 19320
rect 375576 7410 375604 19314
rect 375564 7404 375616 7410
rect 375564 7346 375616 7352
rect 375380 6248 375432 6254
rect 375380 6190 375432 6196
rect 375288 3052 375340 3058
rect 375288 2994 375340 3000
rect 376036 2922 376064 337690
rect 376956 337550 376984 340068
rect 377232 340054 377522 340082
rect 378166 340054 378364 340082
rect 376944 337544 376996 337550
rect 376944 337486 376996 337492
rect 377232 335594 377260 340054
rect 376956 335566 377260 335594
rect 378232 335640 378284 335646
rect 378232 335582 378284 335588
rect 376956 321722 376984 335566
rect 376956 321694 377076 321722
rect 377048 318866 377076 321694
rect 376956 318838 377076 318866
rect 376956 318782 376984 318838
rect 376944 318776 376996 318782
rect 376944 318718 376996 318724
rect 376852 309324 376904 309330
rect 376852 309266 376904 309272
rect 376864 309126 376892 309266
rect 376852 309120 376904 309126
rect 376852 309062 376904 309068
rect 376944 299532 376996 299538
rect 376944 299474 376996 299480
rect 376956 292618 376984 299474
rect 376864 292590 376984 292618
rect 376864 289950 376892 292590
rect 376852 289944 376904 289950
rect 376852 289886 376904 289892
rect 376944 289876 376996 289882
rect 376944 289818 376996 289824
rect 376956 280158 376984 289818
rect 376944 280152 376996 280158
rect 376944 280094 376996 280100
rect 376944 270564 376996 270570
rect 376944 270506 376996 270512
rect 376956 260846 376984 270506
rect 376944 260840 376996 260846
rect 376944 260782 376996 260788
rect 376944 251252 376996 251258
rect 376944 251194 376996 251200
rect 376956 241505 376984 251194
rect 376758 241496 376814 241505
rect 376758 241431 376814 241440
rect 376942 241496 376998 241505
rect 376942 241431 376998 241440
rect 376772 231878 376800 241431
rect 376760 231872 376812 231878
rect 376760 231814 376812 231820
rect 376944 231872 376996 231878
rect 376944 231814 376996 231820
rect 376956 222193 376984 231814
rect 376758 222184 376814 222193
rect 376758 222119 376814 222128
rect 376942 222184 376998 222193
rect 376942 222119 376998 222128
rect 376772 212566 376800 222119
rect 376760 212560 376812 212566
rect 376760 212502 376812 212508
rect 376944 212560 376996 212566
rect 376944 212502 376996 212508
rect 376956 202881 376984 212502
rect 376758 202872 376814 202881
rect 376758 202807 376814 202816
rect 376942 202872 376998 202881
rect 376942 202807 376998 202816
rect 376772 193254 376800 202807
rect 376760 193248 376812 193254
rect 376760 193190 376812 193196
rect 376944 193248 376996 193254
rect 376944 193190 376996 193196
rect 376956 183569 376984 193190
rect 376758 183560 376814 183569
rect 376758 183495 376814 183504
rect 376942 183560 376998 183569
rect 376942 183495 376998 183504
rect 376772 173942 376800 183495
rect 376760 173936 376812 173942
rect 376760 173878 376812 173884
rect 376944 173936 376996 173942
rect 376944 173878 376996 173884
rect 376956 164218 376984 173878
rect 376760 164212 376812 164218
rect 376760 164154 376812 164160
rect 376944 164212 376996 164218
rect 376944 164154 376996 164160
rect 376772 154601 376800 164154
rect 376758 154592 376814 154601
rect 376758 154527 376814 154536
rect 376942 154592 376998 154601
rect 376942 154527 376998 154536
rect 376956 144906 376984 154527
rect 376760 144900 376812 144906
rect 376760 144842 376812 144848
rect 376944 144900 376996 144906
rect 376944 144842 376996 144848
rect 376772 135289 376800 144842
rect 376758 135280 376814 135289
rect 376758 135215 376814 135224
rect 376942 135280 376998 135289
rect 376942 135215 376998 135224
rect 376956 125594 376984 135215
rect 376944 125588 376996 125594
rect 376944 125530 376996 125536
rect 376944 116000 376996 116006
rect 376944 115942 376996 115948
rect 376956 106282 376984 115942
rect 376944 106276 376996 106282
rect 376944 106218 376996 106224
rect 376944 96688 376996 96694
rect 376944 96630 376996 96636
rect 376956 80102 376984 96630
rect 376944 80096 376996 80102
rect 376944 80038 376996 80044
rect 376944 79960 376996 79966
rect 376944 79902 376996 79908
rect 376956 60738 376984 79902
rect 376864 60710 376984 60738
rect 376864 60602 376892 60710
rect 376864 60574 376984 60602
rect 376956 57934 376984 60574
rect 376944 57928 376996 57934
rect 376944 57870 376996 57876
rect 377036 57928 377088 57934
rect 377036 57870 377088 57876
rect 377048 38690 377076 57870
rect 376944 38684 376996 38690
rect 376944 38626 376996 38632
rect 377036 38684 377088 38690
rect 377036 38626 377088 38632
rect 376956 33810 376984 38626
rect 376864 33782 376984 33810
rect 376864 26194 376892 33782
rect 376864 26166 376984 26194
rect 376956 6322 376984 26166
rect 378244 6390 378272 335582
rect 378336 10334 378364 340054
rect 378428 340054 378810 340082
rect 379072 340054 379362 340082
rect 379624 340054 380006 340082
rect 378324 10328 378376 10334
rect 378324 10270 378376 10276
rect 378232 6384 378284 6390
rect 378232 6326 378284 6332
rect 376944 6316 376996 6322
rect 376944 6258 376996 6264
rect 376392 5092 376444 5098
rect 376392 5034 376444 5040
rect 376024 2916 376076 2922
rect 376024 2858 376076 2864
rect 376404 480 376432 5034
rect 378428 3534 378456 340054
rect 378506 337512 378562 337521
rect 378506 337447 378562 337456
rect 378520 337346 378548 337447
rect 378508 337340 378560 337346
rect 378508 337282 378560 337288
rect 379072 335646 379100 340054
rect 379060 335640 379112 335646
rect 379060 335582 379112 335588
rect 379624 10470 379652 340054
rect 380636 337618 380664 340068
rect 380912 340054 381202 340082
rect 381372 340054 381846 340082
rect 380624 337612 380676 337618
rect 380624 337554 380676 337560
rect 380806 183560 380862 183569
rect 380806 183495 380862 183504
rect 380820 173942 380848 183495
rect 380808 173936 380860 173942
rect 380808 173878 380860 173884
rect 379612 10464 379664 10470
rect 379612 10406 379664 10412
rect 379980 6248 380032 6254
rect 379980 6190 380032 6196
rect 378416 3528 378468 3534
rect 378416 3470 378468 3476
rect 378876 3052 378928 3058
rect 378876 2994 378928 3000
rect 377588 2984 377640 2990
rect 377588 2926 377640 2932
rect 377600 480 377628 2926
rect 378888 1578 378916 2994
rect 378796 1550 378916 1578
rect 378796 480 378824 1550
rect 379992 480 380020 6190
rect 380912 5302 380940 340054
rect 381372 336734 381400 340054
rect 382476 336802 382504 340068
rect 381544 336796 381596 336802
rect 381544 336738 381596 336744
rect 382464 336796 382516 336802
rect 382464 336738 382516 336744
rect 380992 336728 381044 336734
rect 380992 336670 381044 336676
rect 381360 336728 381412 336734
rect 381360 336670 381412 336676
rect 381004 328386 381032 336670
rect 381004 328358 381124 328386
rect 381096 318782 381124 328358
rect 381084 318776 381136 318782
rect 381084 318718 381136 318724
rect 381268 318776 381320 318782
rect 381268 318718 381320 318724
rect 381280 317422 381308 318718
rect 381268 317416 381320 317422
rect 381268 317358 381320 317364
rect 381268 307828 381320 307834
rect 381268 307770 381320 307776
rect 381280 304314 381308 307770
rect 381280 304286 381400 304314
rect 381372 289882 381400 304286
rect 381084 289876 381136 289882
rect 381084 289818 381136 289824
rect 381360 289876 381412 289882
rect 381360 289818 381412 289824
rect 381096 282946 381124 289818
rect 381084 282940 381136 282946
rect 381084 282882 381136 282888
rect 381176 282804 381228 282810
rect 381176 282746 381228 282752
rect 381188 280106 381216 282746
rect 381004 280078 381216 280106
rect 381004 270570 381032 280078
rect 380992 270564 381044 270570
rect 380992 270506 381044 270512
rect 381084 270564 381136 270570
rect 381084 270506 381136 270512
rect 381096 270434 381124 270506
rect 381084 270428 381136 270434
rect 381084 270370 381136 270376
rect 381176 260908 381228 260914
rect 381176 260850 381228 260856
rect 381188 260817 381216 260850
rect 381174 260808 381230 260817
rect 381174 260743 381230 260752
rect 381358 260808 381414 260817
rect 381358 260743 381414 260752
rect 381372 251258 381400 260743
rect 381084 251252 381136 251258
rect 381084 251194 381136 251200
rect 381360 251252 381412 251258
rect 381360 251194 381412 251200
rect 381096 251122 381124 251194
rect 381084 251116 381136 251122
rect 381084 251058 381136 251064
rect 381188 241534 381216 241565
rect 381176 241528 381228 241534
rect 381096 241476 381176 241482
rect 381096 241470 381228 241476
rect 381096 241454 381216 241470
rect 381096 234734 381124 241454
rect 381084 234728 381136 234734
rect 381084 234670 381136 234676
rect 381176 231872 381228 231878
rect 381176 231814 381228 231820
rect 381188 225010 381216 231814
rect 381176 225004 381228 225010
rect 381176 224946 381228 224952
rect 381188 222222 381216 222253
rect 381176 222216 381228 222222
rect 381096 222164 381176 222170
rect 381096 222158 381228 222164
rect 381096 222142 381216 222158
rect 381096 215422 381124 222142
rect 381084 215416 381136 215422
rect 381084 215358 381136 215364
rect 381176 212560 381228 212566
rect 381176 212502 381228 212508
rect 381188 205698 381216 212502
rect 381176 205692 381228 205698
rect 381176 205634 381228 205640
rect 381176 205556 381228 205562
rect 381176 205498 381228 205504
rect 381188 202858 381216 205498
rect 381096 202830 381216 202858
rect 381096 201482 381124 202830
rect 381084 201476 381136 201482
rect 381084 201418 381136 201424
rect 381360 201476 381412 201482
rect 381360 201418 381412 201424
rect 381188 183598 381216 183629
rect 381372 183598 381400 201418
rect 381176 183592 381228 183598
rect 381082 183560 381138 183569
rect 381138 183540 381176 183546
rect 381138 183534 381228 183540
rect 381360 183592 381412 183598
rect 381360 183534 381412 183540
rect 381138 183518 381216 183534
rect 381082 183495 381138 183504
rect 380992 173936 381044 173942
rect 380992 173878 381044 173884
rect 381004 171306 381032 173878
rect 381004 171278 381124 171306
rect 381096 164150 381124 171278
rect 380992 164144 381044 164150
rect 380992 164086 381044 164092
rect 381084 164144 381136 164150
rect 381084 164086 381136 164092
rect 381004 162858 381032 164086
rect 380992 162852 381044 162858
rect 380992 162794 381044 162800
rect 381084 147620 381136 147626
rect 381084 147562 381136 147568
rect 381096 144922 381124 147562
rect 381096 144894 381216 144922
rect 381188 144888 381216 144894
rect 381188 144860 381308 144888
rect 381280 135318 381308 144860
rect 381084 135312 381136 135318
rect 381084 135254 381136 135260
rect 381268 135312 381320 135318
rect 381268 135254 381320 135260
rect 381096 128382 381124 135254
rect 381450 134600 381506 134609
rect 381450 134535 381506 134544
rect 381464 134065 381492 134535
rect 381450 134056 381506 134065
rect 381450 133991 381506 134000
rect 381084 128376 381136 128382
rect 381084 128318 381136 128324
rect 381176 128308 381228 128314
rect 381176 128250 381228 128256
rect 381188 125576 381216 128250
rect 381188 125548 381308 125576
rect 381280 116113 381308 125548
rect 381266 116104 381322 116113
rect 381266 116039 381322 116048
rect 381082 115968 381138 115977
rect 381082 115903 381084 115912
rect 381136 115903 381138 115912
rect 381268 115932 381320 115938
rect 381084 115874 381136 115880
rect 381268 115874 381320 115880
rect 381280 96642 381308 115874
rect 381188 96614 381308 96642
rect 381188 77314 381216 96614
rect 381084 77308 381136 77314
rect 381084 77250 381136 77256
rect 381176 77308 381228 77314
rect 381176 77250 381228 77256
rect 381096 50946 381124 77250
rect 381096 50918 381216 50946
rect 381188 48278 381216 50918
rect 381176 48272 381228 48278
rect 381176 48214 381228 48220
rect 381268 48272 381320 48278
rect 381268 48214 381320 48220
rect 381280 29034 381308 48214
rect 381176 29028 381228 29034
rect 381176 28970 381228 28976
rect 381268 29028 381320 29034
rect 381268 28970 381320 28976
rect 381188 19666 381216 28970
rect 381188 19638 381308 19666
rect 381280 19378 381308 19638
rect 381084 19372 381136 19378
rect 381084 19314 381136 19320
rect 381268 19372 381320 19378
rect 381268 19314 381320 19320
rect 381096 17950 381124 19314
rect 381084 17944 381136 17950
rect 381084 17886 381136 17892
rect 380992 8356 381044 8362
rect 380992 8298 381044 8304
rect 381004 6730 381032 8298
rect 380992 6724 381044 6730
rect 380992 6666 381044 6672
rect 380900 5296 380952 5302
rect 380900 5238 380952 5244
rect 381556 3602 381584 336738
rect 382660 331242 382688 340190
rect 383686 340054 383792 340082
rect 382924 336796 382976 336802
rect 382924 336738 382976 336744
rect 382476 331214 382688 331242
rect 382476 318782 382504 331214
rect 382280 318776 382332 318782
rect 382280 318718 382332 318724
rect 382464 318776 382516 318782
rect 382464 318718 382516 318724
rect 382292 317422 382320 318718
rect 382280 317416 382332 317422
rect 382280 317358 382332 317364
rect 382464 302116 382516 302122
rect 382464 302058 382516 302064
rect 382476 299470 382504 302058
rect 382464 299464 382516 299470
rect 382464 299406 382516 299412
rect 382464 289876 382516 289882
rect 382464 289818 382516 289824
rect 382476 273222 382504 289818
rect 382464 273216 382516 273222
rect 382464 273158 382516 273164
rect 382464 273080 382516 273086
rect 382464 273022 382516 273028
rect 382476 253910 382504 273022
rect 382464 253904 382516 253910
rect 382464 253846 382516 253852
rect 382464 253768 382516 253774
rect 382464 253710 382516 253716
rect 382476 234598 382504 253710
rect 382464 234592 382516 234598
rect 382464 234534 382516 234540
rect 382464 234456 382516 234462
rect 382464 234398 382516 234404
rect 382476 215286 382504 234398
rect 382464 215280 382516 215286
rect 382464 215222 382516 215228
rect 382464 215144 382516 215150
rect 382464 215086 382516 215092
rect 382476 195974 382504 215086
rect 382464 195968 382516 195974
rect 382464 195910 382516 195916
rect 382464 195832 382516 195838
rect 382464 195774 382516 195780
rect 382476 176662 382504 195774
rect 382464 176656 382516 176662
rect 382464 176598 382516 176604
rect 382464 176520 382516 176526
rect 382464 176462 382516 176468
rect 382476 157350 382504 176462
rect 382464 157344 382516 157350
rect 382464 157286 382516 157292
rect 382464 157208 382516 157214
rect 382464 157150 382516 157156
rect 382476 80102 382504 157150
rect 382464 80096 382516 80102
rect 382464 80038 382516 80044
rect 382464 79960 382516 79966
rect 382464 79902 382516 79908
rect 382476 60738 382504 79902
rect 382384 60710 382504 60738
rect 382384 60602 382412 60710
rect 382384 60574 382504 60602
rect 382476 57934 382504 60574
rect 382464 57928 382516 57934
rect 382464 57870 382516 57876
rect 382372 48340 382424 48346
rect 382372 48282 382424 48288
rect 382384 38758 382412 48282
rect 382372 38752 382424 38758
rect 382372 38694 382424 38700
rect 382372 38616 382424 38622
rect 382372 38558 382424 38564
rect 382384 33810 382412 38558
rect 382292 33782 382412 33810
rect 382292 19378 382320 33782
rect 382280 19372 382332 19378
rect 382280 19314 382332 19320
rect 382464 19372 382516 19378
rect 382464 19314 382516 19320
rect 382476 17950 382504 19314
rect 382464 17944 382516 17950
rect 382464 17886 382516 17892
rect 382372 8356 382424 8362
rect 382372 8298 382424 8304
rect 382384 5370 382412 8298
rect 382372 5364 382424 5370
rect 382372 5306 382424 5312
rect 382936 3670 382964 336738
rect 383764 10402 383792 340054
rect 384040 340054 384330 340082
rect 384040 337550 384068 340054
rect 384028 337544 384080 337550
rect 384028 337486 384080 337492
rect 384408 331242 384436 340190
rect 383856 331214 384436 331242
rect 385144 340054 385526 340082
rect 383752 10396 383804 10402
rect 383752 10338 383804 10344
rect 383856 5438 383884 331214
rect 385144 6662 385172 340054
rect 385684 337952 385736 337958
rect 385684 337894 385736 337900
rect 385132 6656 385184 6662
rect 385132 6598 385184 6604
rect 383844 5432 383896 5438
rect 383844 5374 383896 5380
rect 383568 5160 383620 5166
rect 383568 5102 383620 5108
rect 382924 3664 382976 3670
rect 382924 3606 382976 3612
rect 381544 3596 381596 3602
rect 381544 3538 381596 3544
rect 382372 3528 382424 3534
rect 382372 3470 382424 3476
rect 381176 3188 381228 3194
rect 381176 3130 381228 3136
rect 381188 480 381216 3130
rect 382384 480 382412 3470
rect 383580 480 383608 5102
rect 384672 2916 384724 2922
rect 384672 2858 384724 2864
rect 384684 480 384712 2858
rect 385696 2854 385724 337894
rect 386156 336802 386184 340068
rect 386432 340054 386722 340082
rect 386892 340054 387366 340082
rect 386144 336796 386196 336802
rect 386144 336738 386196 336744
rect 386326 170368 386382 170377
rect 386326 170303 386382 170312
rect 386340 169969 386368 170303
rect 386326 169960 386382 169969
rect 386326 169895 386382 169904
rect 386432 6458 386460 340054
rect 386892 331242 386920 340054
rect 387996 337890 388024 340068
rect 388180 340054 388562 340082
rect 389206 340054 389312 340082
rect 387984 337884 388036 337890
rect 387984 337826 388036 337832
rect 388180 331242 388208 340054
rect 389088 337544 389140 337550
rect 389088 337486 389140 337492
rect 386616 331214 386920 331242
rect 387996 331214 388208 331242
rect 386616 331106 386644 331214
rect 386616 331078 386736 331106
rect 386708 321314 386736 331078
rect 386616 321286 386736 321314
rect 386616 318730 386644 321286
rect 387996 318782 388024 331214
rect 387892 318776 387944 318782
rect 386616 318702 386736 318730
rect 387892 318718 387944 318724
rect 387984 318776 388036 318782
rect 387984 318718 388036 318724
rect 386708 292618 386736 318702
rect 387904 317422 387932 318718
rect 387892 317416 387944 317422
rect 387892 317358 387944 317364
rect 387892 307828 387944 307834
rect 387892 307770 387944 307776
rect 387904 304910 387932 307770
rect 387892 304904 387944 304910
rect 387892 304846 387944 304852
rect 387984 298172 388036 298178
rect 387984 298114 388036 298120
rect 387996 292670 388024 298114
rect 386616 292590 386736 292618
rect 387984 292664 388036 292670
rect 387984 292606 388036 292612
rect 386616 285002 386644 292590
rect 387984 292528 388036 292534
rect 387984 292470 388036 292476
rect 386616 284974 386828 285002
rect 386800 282826 386828 284974
rect 386708 282798 386828 282826
rect 386708 280158 386736 282798
rect 387996 280158 388024 292470
rect 386696 280152 386748 280158
rect 386696 280094 386748 280100
rect 386788 280152 386840 280158
rect 386788 280094 386840 280100
rect 387984 280152 388036 280158
rect 387984 280094 388036 280100
rect 388076 280152 388128 280158
rect 388076 280094 388128 280100
rect 386800 270609 386828 280094
rect 388088 273170 388116 280094
rect 387996 273142 388116 273170
rect 386786 270600 386842 270609
rect 386786 270535 386842 270544
rect 386694 270464 386750 270473
rect 386694 270399 386750 270408
rect 386708 249898 386736 270399
rect 387996 253994 388024 273142
rect 387904 253966 388024 253994
rect 387904 253858 387932 253966
rect 387904 253830 388024 253858
rect 386604 249892 386656 249898
rect 386604 249834 386656 249840
rect 386696 249892 386748 249898
rect 386696 249834 386748 249840
rect 386616 249778 386644 249834
rect 386616 249750 386736 249778
rect 386708 244322 386736 249750
rect 386696 244316 386748 244322
rect 386696 244258 386748 244264
rect 386604 244248 386656 244254
rect 386604 244190 386656 244196
rect 386616 225010 386644 244190
rect 386604 225004 386656 225010
rect 386604 224946 386656 224952
rect 386696 224868 386748 224874
rect 386696 224810 386748 224816
rect 386708 217410 386736 224810
rect 386616 217382 386736 217410
rect 386616 212537 386644 217382
rect 386602 212528 386658 212537
rect 386602 212463 386658 212472
rect 386786 212528 386842 212537
rect 386786 212463 386842 212472
rect 386800 193322 386828 212463
rect 386604 193316 386656 193322
rect 386604 193258 386656 193264
rect 386788 193316 386840 193322
rect 386788 193258 386840 193264
rect 386616 193225 386644 193258
rect 386602 193216 386658 193225
rect 386602 193151 386658 193160
rect 386786 193216 386842 193225
rect 386786 193151 386842 193160
rect 386800 182238 386828 193151
rect 386696 182232 386748 182238
rect 386696 182174 386748 182180
rect 386788 182232 386840 182238
rect 386788 182174 386840 182180
rect 386708 180810 386736 182174
rect 386696 180804 386748 180810
rect 386696 180746 386748 180752
rect 387996 176746 388024 253830
rect 387904 176718 388024 176746
rect 387904 176610 387932 176718
rect 387904 176582 388024 176610
rect 386604 171148 386656 171154
rect 386604 171090 386656 171096
rect 386616 162858 386644 171090
rect 387996 162858 388024 176582
rect 386604 162852 386656 162858
rect 386604 162794 386656 162800
rect 386788 162852 386840 162858
rect 386788 162794 386840 162800
rect 387984 162852 388036 162858
rect 387984 162794 388036 162800
rect 386800 135289 386828 162794
rect 387984 158024 388036 158030
rect 387984 157966 388036 157972
rect 387996 138122 388024 157966
rect 387904 138094 388024 138122
rect 387904 137714 387932 138094
rect 387904 137686 388024 137714
rect 386602 135280 386658 135289
rect 386602 135215 386658 135224
rect 386786 135280 386842 135289
rect 386786 135215 386842 135224
rect 386616 130370 386644 135215
rect 386616 130342 386736 130370
rect 386708 125594 386736 130342
rect 387996 125594 388024 137686
rect 386696 125588 386748 125594
rect 386696 125530 386748 125536
rect 386788 125588 386840 125594
rect 386788 125530 386840 125536
rect 387984 125588 388036 125594
rect 387984 125530 388036 125536
rect 388076 125588 388128 125594
rect 388076 125530 388128 125536
rect 386800 115977 386828 125530
rect 388088 118658 388116 125530
rect 387984 118652 388036 118658
rect 387984 118594 388036 118600
rect 388076 118652 388128 118658
rect 388076 118594 388128 118600
rect 386602 115968 386658 115977
rect 386602 115903 386604 115912
rect 386656 115903 386658 115912
rect 386786 115968 386842 115977
rect 386786 115903 386788 115912
rect 386604 115874 386656 115880
rect 386840 115903 386842 115912
rect 386788 115874 386840 115880
rect 386800 96665 386828 115874
rect 387996 114510 388024 118594
rect 387984 114504 388036 114510
rect 387984 114446 388036 114452
rect 387984 104916 388036 104922
rect 387984 104858 388036 104864
rect 386602 96656 386658 96665
rect 386602 96591 386658 96600
rect 386786 96656 386842 96665
rect 386786 96591 386842 96600
rect 386616 86902 386644 96591
rect 387996 95198 388024 104858
rect 387984 95192 388036 95198
rect 387984 95134 388036 95140
rect 386604 86896 386656 86902
rect 386604 86838 386656 86844
rect 387984 85604 388036 85610
rect 387984 85546 388036 85552
rect 386604 77308 386656 77314
rect 386604 77250 386656 77256
rect 386616 67726 386644 77250
rect 387996 75886 388024 85546
rect 387984 75880 388036 75886
rect 387984 75822 388036 75828
rect 388168 75880 388220 75886
rect 388168 75822 388220 75828
rect 386604 67720 386656 67726
rect 386604 67662 386656 67668
rect 386696 67652 386748 67658
rect 386696 67594 386748 67600
rect 386708 58002 386736 67594
rect 388180 66337 388208 75822
rect 387982 66328 388038 66337
rect 387982 66263 388038 66272
rect 388166 66328 388222 66337
rect 388166 66263 388222 66272
rect 387996 66230 388024 66263
rect 387984 66224 388036 66230
rect 387984 66166 388036 66172
rect 386604 57996 386656 58002
rect 386604 57938 386656 57944
rect 386696 57996 386748 58002
rect 386696 57938 386748 57944
rect 386616 48346 386644 57938
rect 388076 56636 388128 56642
rect 388076 56578 388128 56584
rect 388088 48346 388116 56578
rect 386604 48340 386656 48346
rect 386604 48282 386656 48288
rect 386696 48340 386748 48346
rect 386696 48282 386748 48288
rect 387892 48340 387944 48346
rect 387892 48282 387944 48288
rect 388076 48340 388128 48346
rect 388076 48282 388128 48288
rect 386708 37398 386736 48282
rect 387904 46918 387932 48282
rect 387892 46912 387944 46918
rect 387892 46854 387944 46860
rect 386696 37392 386748 37398
rect 386696 37334 386748 37340
rect 386788 37324 386840 37330
rect 386788 37266 386840 37272
rect 387892 37324 387944 37330
rect 387892 37266 387944 37272
rect 386800 37210 386828 37266
rect 386708 37182 386828 37210
rect 386708 29034 386736 37182
rect 386696 29028 386748 29034
rect 386696 28970 386748 28976
rect 386788 28892 386840 28898
rect 386788 28834 386840 28840
rect 386800 19038 386828 28834
rect 387904 27810 387932 37266
rect 387892 27804 387944 27810
rect 387892 27746 387944 27752
rect 387800 27668 387852 27674
rect 387800 27610 387852 27616
rect 387812 19122 387840 27610
rect 387812 19094 388116 19122
rect 386788 19032 386840 19038
rect 386788 18974 386840 18980
rect 386788 18896 386840 18902
rect 386788 18838 386840 18844
rect 386510 16824 386566 16833
rect 386510 16759 386566 16768
rect 386524 16561 386552 16759
rect 386510 16552 386566 16561
rect 386510 16487 386566 16496
rect 386800 9722 386828 18838
rect 388088 9722 388116 19094
rect 386512 9716 386564 9722
rect 386512 9658 386564 9664
rect 386788 9716 386840 9722
rect 386788 9658 386840 9664
rect 387892 9716 387944 9722
rect 387892 9658 387944 9664
rect 388076 9716 388128 9722
rect 388076 9658 388128 9664
rect 386524 6798 386552 9658
rect 386512 6792 386564 6798
rect 386512 6734 386564 6740
rect 387904 6526 387932 9658
rect 387892 6520 387944 6526
rect 387892 6462 387944 6468
rect 386420 6452 386472 6458
rect 386420 6394 386472 6400
rect 387064 5228 387116 5234
rect 387064 5170 387116 5176
rect 385868 3732 385920 3738
rect 385868 3674 385920 3680
rect 385684 2848 385736 2854
rect 385684 2790 385736 2796
rect 385880 480 385908 3674
rect 387076 480 387104 5170
rect 389100 3670 389128 337486
rect 389284 9042 389312 340054
rect 389744 337958 389772 340068
rect 389836 340054 390402 340082
rect 390664 340054 391046 340082
rect 389732 337952 389784 337958
rect 389732 337894 389784 337900
rect 389836 335730 389864 340054
rect 389916 336796 389968 336802
rect 389916 336738 389968 336744
rect 389376 335702 389864 335730
rect 389272 9036 389324 9042
rect 389272 8978 389324 8984
rect 389376 6594 389404 335702
rect 389928 335594 389956 336738
rect 389836 335566 389956 335594
rect 389364 6588 389416 6594
rect 389364 6530 389416 6536
rect 389836 3806 389864 335566
rect 390664 9178 390692 340054
rect 391204 337884 391256 337890
rect 391204 337826 391256 337832
rect 390652 9172 390704 9178
rect 390652 9114 390704 9120
rect 390652 5296 390704 5302
rect 390652 5238 390704 5244
rect 389824 3800 389876 3806
rect 389824 3742 389876 3748
rect 388260 3664 388312 3670
rect 388260 3606 388312 3612
rect 389088 3664 389140 3670
rect 389088 3606 389140 3612
rect 388272 480 388300 3606
rect 389456 3596 389508 3602
rect 389456 3538 389508 3544
rect 389468 480 389496 3538
rect 390664 480 390692 5238
rect 391216 4026 391244 337826
rect 391584 337618 391612 340068
rect 391952 340054 392242 340082
rect 392412 340054 392886 340082
rect 391572 337612 391624 337618
rect 391572 337554 391624 337560
rect 391952 5506 391980 340054
rect 392412 335594 392440 340054
rect 393136 337612 393188 337618
rect 393136 337554 393188 337560
rect 392136 335566 392440 335594
rect 392136 331106 392164 335566
rect 393148 331294 393176 337554
rect 393424 336802 393452 340068
rect 393516 340054 394082 340082
rect 394726 340054 394832 340082
rect 393412 336796 393464 336802
rect 393412 336738 393464 336744
rect 393136 331288 393188 331294
rect 393136 331230 393188 331236
rect 392136 331078 392256 331106
rect 392228 321638 392256 331078
rect 393044 327140 393096 327146
rect 393044 327082 393096 327088
rect 393056 324222 393084 327082
rect 393044 324216 393096 324222
rect 393044 324158 393096 324164
rect 392216 321632 392268 321638
rect 392216 321574 392268 321580
rect 392124 318844 392176 318850
rect 392124 318786 392176 318792
rect 392136 318730 392164 318786
rect 392136 318702 392256 318730
rect 392228 292618 392256 318702
rect 393228 309188 393280 309194
rect 393228 309130 393280 309136
rect 392136 292590 392256 292618
rect 392136 289814 392164 292590
rect 392124 289808 392176 289814
rect 392124 289750 392176 289756
rect 392216 289808 392268 289814
rect 392216 289750 392268 289756
rect 392228 278798 392256 289750
rect 393240 280158 393268 309130
rect 393228 280152 393280 280158
rect 393228 280094 393280 280100
rect 392124 278792 392176 278798
rect 392124 278734 392176 278740
rect 392216 278792 392268 278798
rect 392216 278734 392268 278740
rect 392136 270502 392164 278734
rect 393228 270564 393280 270570
rect 393228 270506 393280 270512
rect 392124 270496 392176 270502
rect 392124 270438 392176 270444
rect 392216 264308 392268 264314
rect 392216 264250 392268 264256
rect 392228 249898 392256 264250
rect 392124 249892 392176 249898
rect 392124 249834 392176 249840
rect 392216 249892 392268 249898
rect 392216 249834 392268 249840
rect 392136 249801 392164 249834
rect 392122 249792 392178 249801
rect 392122 249727 392178 249736
rect 392398 249792 392454 249801
rect 392398 249727 392454 249736
rect 392412 240174 392440 249727
rect 393240 241482 393268 270506
rect 393148 241454 393268 241482
rect 392216 240168 392268 240174
rect 392216 240110 392268 240116
rect 392400 240168 392452 240174
rect 392400 240110 392452 240116
rect 392228 236774 392256 240110
rect 392216 236768 392268 236774
rect 392216 236710 392268 236716
rect 393148 231878 393176 241454
rect 393136 231872 393188 231878
rect 393228 231872 393280 231878
rect 393136 231814 393188 231820
rect 393226 231840 393228 231849
rect 393280 231840 393282 231849
rect 393226 231775 393282 231784
rect 393410 231840 393466 231849
rect 393410 231775 393466 231784
rect 393240 222222 393268 222253
rect 393424 222222 393452 231775
rect 392216 222216 392268 222222
rect 393228 222216 393280 222222
rect 392216 222158 392268 222164
rect 393148 222164 393228 222170
rect 393148 222158 393280 222164
rect 393412 222216 393464 222222
rect 393412 222158 393464 222164
rect 392228 217410 392256 222158
rect 392136 217382 392256 217410
rect 393148 222142 393268 222158
rect 392136 212537 392164 217382
rect 393148 212566 393176 222142
rect 393136 212560 393188 212566
rect 392122 212528 392178 212537
rect 392122 212463 392178 212472
rect 392306 212528 392362 212537
rect 393228 212560 393280 212566
rect 393136 212502 393188 212508
rect 393226 212528 393228 212537
rect 393280 212528 393282 212537
rect 392306 212463 392362 212472
rect 393226 212463 393282 212472
rect 393410 212528 393466 212537
rect 393410 212463 393466 212472
rect 392320 195294 392348 212463
rect 393240 202910 393268 202941
rect 393424 202910 393452 212463
rect 393228 202904 393280 202910
rect 393148 202852 393228 202858
rect 393148 202846 393280 202852
rect 393412 202904 393464 202910
rect 393412 202846 393464 202852
rect 393148 202830 393268 202846
rect 392032 195288 392084 195294
rect 392032 195230 392084 195236
rect 392308 195288 392360 195294
rect 392308 195230 392360 195236
rect 392044 190505 392072 195230
rect 393148 193254 393176 202830
rect 393136 193248 393188 193254
rect 393228 193248 393280 193254
rect 393136 193190 393188 193196
rect 393226 193216 393228 193225
rect 393280 193216 393282 193225
rect 393226 193151 393282 193160
rect 393410 193216 393466 193225
rect 393410 193151 393466 193160
rect 392030 190496 392086 190505
rect 392030 190431 392086 190440
rect 392214 190496 392270 190505
rect 392214 190431 392270 190440
rect 392228 182322 392256 190431
rect 393424 183598 393452 193151
rect 393228 183592 393280 183598
rect 393228 183534 393280 183540
rect 393412 183592 393464 183598
rect 393412 183534 393464 183540
rect 392136 182294 392256 182322
rect 392136 182186 392164 182294
rect 392136 182158 392256 182186
rect 392228 180810 392256 182158
rect 392216 180804 392268 180810
rect 392216 180746 392268 180752
rect 392124 171148 392176 171154
rect 392124 171090 392176 171096
rect 392136 162858 392164 171090
rect 392124 162852 392176 162858
rect 392124 162794 392176 162800
rect 392308 162852 392360 162858
rect 392308 162794 392360 162800
rect 392320 148374 392348 162794
rect 393240 154562 393268 183534
rect 393228 154556 393280 154562
rect 393228 154498 393280 154504
rect 393412 154556 393464 154562
rect 393412 154498 393464 154504
rect 392308 148368 392360 148374
rect 392308 148310 392360 148316
rect 393424 144945 393452 154498
rect 393226 144936 393282 144945
rect 393226 144871 393228 144880
rect 393280 144871 393282 144880
rect 393410 144936 393466 144945
rect 393410 144871 393466 144880
rect 393228 144842 393280 144848
rect 392124 135312 392176 135318
rect 392124 135254 392176 135260
rect 393228 135312 393280 135318
rect 393228 135254 393280 135260
rect 392136 130370 392164 135254
rect 392136 130342 392256 130370
rect 392228 125594 392256 130342
rect 393240 125594 393268 135254
rect 392216 125588 392268 125594
rect 392216 125530 392268 125536
rect 392308 125588 392360 125594
rect 392308 125530 392360 125536
rect 393228 125588 393280 125594
rect 393228 125530 393280 125536
rect 392320 115977 392348 125530
rect 393228 116000 393280 116006
rect 392122 115968 392178 115977
rect 392122 115903 392124 115912
rect 392176 115903 392178 115912
rect 392306 115968 392362 115977
rect 393228 115942 393280 115948
rect 392306 115903 392308 115912
rect 392124 115874 392176 115880
rect 392360 115903 392362 115912
rect 392308 115874 392360 115880
rect 392320 96665 392348 115874
rect 393240 115870 393268 115942
rect 393228 115864 393280 115870
rect 393228 115806 393280 115812
rect 393320 115864 393372 115870
rect 393320 115806 393372 115812
rect 393332 106298 393360 115806
rect 393240 106282 393360 106298
rect 393228 106276 393360 106282
rect 393280 106270 393360 106276
rect 393412 106276 393464 106282
rect 393228 106218 393280 106224
rect 393412 106218 393464 106224
rect 393424 96665 393452 106218
rect 392122 96656 392178 96665
rect 392122 96591 392178 96600
rect 392306 96656 392362 96665
rect 392306 96591 392362 96600
rect 393226 96656 393282 96665
rect 393226 96591 393282 96600
rect 393410 96656 393466 96665
rect 393410 96591 393466 96600
rect 392136 86902 392164 96591
rect 393240 95198 393268 96591
rect 393228 95192 393280 95198
rect 393228 95134 393280 95140
rect 392124 86896 392176 86902
rect 392124 86838 392176 86844
rect 393412 85604 393464 85610
rect 393412 85546 393464 85552
rect 392124 77308 392176 77314
rect 392124 77250 392176 77256
rect 392136 67726 392164 77250
rect 393424 67833 393452 85546
rect 393410 67824 393466 67833
rect 393410 67759 393466 67768
rect 392124 67720 392176 67726
rect 392124 67662 392176 67668
rect 393226 67688 393282 67697
rect 392216 67652 392268 67658
rect 393226 67623 393282 67632
rect 392216 67594 392268 67600
rect 392228 61742 392256 67594
rect 393240 67590 393268 67623
rect 393228 67584 393280 67590
rect 393228 67526 393280 67532
rect 392216 61736 392268 61742
rect 392216 61678 392268 61684
rect 392400 61736 392452 61742
rect 392400 61678 392452 61684
rect 392412 56658 392440 61678
rect 393228 57996 393280 58002
rect 393228 57938 393280 57944
rect 392320 56630 392440 56658
rect 392320 56574 392348 56630
rect 392308 56568 392360 56574
rect 392308 56510 392360 56516
rect 392124 47048 392176 47054
rect 392124 46990 392176 46996
rect 392136 46918 392164 46990
rect 392124 46912 392176 46918
rect 392124 46854 392176 46860
rect 392124 46776 392176 46782
rect 392124 46718 392176 46724
rect 392136 33810 392164 46718
rect 392044 33782 392164 33810
rect 392044 31634 392072 33782
rect 392044 31606 392256 31634
rect 392228 28966 392256 31606
rect 393240 28966 393268 57938
rect 392032 28960 392084 28966
rect 392032 28902 392084 28908
rect 392216 28960 392268 28966
rect 392216 28902 392268 28908
rect 393228 28960 393280 28966
rect 393228 28902 393280 28908
rect 392044 19394 392072 28902
rect 392044 19366 392164 19394
rect 392136 14498 392164 19366
rect 393228 19372 393280 19378
rect 393228 19314 393280 19320
rect 393240 14498 393268 19314
rect 392044 14470 392164 14498
rect 393056 14470 393268 14498
rect 392044 9246 392072 14470
rect 393056 9654 393084 14470
rect 393044 9648 393096 9654
rect 393044 9590 393096 9596
rect 392032 9240 392084 9246
rect 392032 9182 392084 9188
rect 391940 5500 391992 5506
rect 391940 5442 391992 5448
rect 393516 4554 393544 340054
rect 394804 9110 394832 340054
rect 395264 338026 395292 340068
rect 395356 340054 395922 340082
rect 396184 340054 396566 340082
rect 395252 338020 395304 338026
rect 395252 337962 395304 337968
rect 395356 335730 395384 340054
rect 395436 336932 395488 336938
rect 395436 336874 395488 336880
rect 394896 335702 395384 335730
rect 394792 9104 394844 9110
rect 394792 9046 394844 9052
rect 394240 5364 394292 5370
rect 394240 5306 394292 5312
rect 393504 4548 393556 4554
rect 393504 4490 393556 4496
rect 391124 3998 391244 4026
rect 391124 3942 391152 3998
rect 391112 3936 391164 3942
rect 391112 3878 391164 3884
rect 391848 3664 391900 3670
rect 391848 3606 391900 3612
rect 391860 480 391888 3606
rect 393044 604 393096 610
rect 393044 546 393096 552
rect 393056 480 393084 546
rect 394252 480 394280 5306
rect 394896 4486 394924 335702
rect 395448 334098 395476 336874
rect 395356 334070 395476 334098
rect 394884 4480 394936 4486
rect 394884 4422 394936 4428
rect 395356 3806 395384 334070
rect 395986 134192 396042 134201
rect 395986 134127 396042 134136
rect 396000 133793 396028 134127
rect 395986 133784 396042 133793
rect 395986 133719 396042 133728
rect 396184 7274 396212 340054
rect 397104 337890 397132 340068
rect 397472 340054 397762 340082
rect 397932 340054 398406 340082
rect 397092 337884 397144 337890
rect 397092 337826 397144 337832
rect 396724 336796 396776 336802
rect 396724 336738 396776 336744
rect 396172 7268 396224 7274
rect 396172 7210 396224 7216
rect 396736 3874 396764 336738
rect 397366 279984 397422 279993
rect 397366 279919 397422 279928
rect 397380 263498 397408 279919
rect 397368 263492 397420 263498
rect 397368 263434 397420 263440
rect 397368 260772 397420 260778
rect 397368 260714 397420 260720
rect 397380 259457 397408 260714
rect 397366 259448 397422 259457
rect 397366 259383 397422 259392
rect 397366 212528 397422 212537
rect 397366 212463 397422 212472
rect 397380 202910 397408 212463
rect 397368 202904 397420 202910
rect 397368 202846 397420 202852
rect 397368 182164 397420 182170
rect 397368 182106 397420 182112
rect 397380 172553 397408 182106
rect 397366 172544 397422 172553
rect 397366 172479 397422 172488
rect 397472 4418 397500 340054
rect 397932 328506 397960 340054
rect 398944 336870 398972 340068
rect 399036 340054 399602 340082
rect 398932 336864 398984 336870
rect 398932 336806 398984 336812
rect 397736 328500 397788 328506
rect 397736 328442 397788 328448
rect 397920 328500 397972 328506
rect 397920 328442 397972 328448
rect 397748 318782 397776 328442
rect 397736 318776 397788 318782
rect 397736 318718 397788 318724
rect 397736 312180 397788 312186
rect 397736 312122 397788 312128
rect 397748 292618 397776 312122
rect 397656 292590 397776 292618
rect 397656 282826 397684 292590
rect 397656 282798 397776 282826
rect 397748 280129 397776 282798
rect 397734 280120 397790 280129
rect 397734 280055 397790 280064
rect 397736 263492 397788 263498
rect 397736 263434 397788 263440
rect 397748 260778 397776 263434
rect 397736 260772 397788 260778
rect 397736 260714 397788 260720
rect 397918 259448 397974 259457
rect 397918 259383 397974 259392
rect 397932 231878 397960 259383
rect 397736 231872 397788 231878
rect 397736 231814 397788 231820
rect 397920 231872 397972 231878
rect 397920 231814 397972 231820
rect 397748 225010 397776 231814
rect 397736 225004 397788 225010
rect 397736 224946 397788 224952
rect 397736 224868 397788 224874
rect 397736 224810 397788 224816
rect 397748 222170 397776 224810
rect 397656 222142 397776 222170
rect 397656 215354 397684 222142
rect 397644 215348 397696 215354
rect 397644 215290 397696 215296
rect 397552 212560 397604 212566
rect 397550 212528 397552 212537
rect 397604 212528 397606 212537
rect 397550 212463 397606 212472
rect 397748 202910 397776 202941
rect 397736 202904 397788 202910
rect 397656 202852 397736 202858
rect 397656 202846 397788 202852
rect 397656 202830 397776 202846
rect 397656 196042 397684 202830
rect 397644 196036 397696 196042
rect 397644 195978 397696 195984
rect 397552 193248 397604 193254
rect 397550 193216 397552 193225
rect 397604 193216 397606 193225
rect 397550 193151 397606 193160
rect 397734 193216 397790 193225
rect 397734 193151 397790 193160
rect 397748 186386 397776 193151
rect 397736 186380 397788 186386
rect 397736 186322 397788 186328
rect 397736 186244 397788 186250
rect 397736 186186 397788 186192
rect 397748 182170 397776 186186
rect 397736 182164 397788 182170
rect 397736 182106 397788 182112
rect 397550 172544 397606 172553
rect 397550 172479 397606 172488
rect 397564 168994 397592 172479
rect 397564 168966 397684 168994
rect 397656 164234 397684 168966
rect 397656 164206 397776 164234
rect 397748 143546 397776 164206
rect 397736 143540 397788 143546
rect 397736 143482 397788 143488
rect 397736 137964 397788 137970
rect 397736 137906 397788 137912
rect 397748 118810 397776 137906
rect 397656 118782 397776 118810
rect 397656 109138 397684 118782
rect 397644 109132 397696 109138
rect 397644 109074 397696 109080
rect 397644 108996 397696 109002
rect 397644 108938 397696 108944
rect 397656 86970 397684 108938
rect 397644 86964 397696 86970
rect 397644 86906 397696 86912
rect 397644 77308 397696 77314
rect 397644 77250 397696 77256
rect 397656 67590 397684 77250
rect 397644 67584 397696 67590
rect 397644 67526 397696 67532
rect 397736 57996 397788 58002
rect 397736 57938 397788 57944
rect 397748 41426 397776 57938
rect 397656 41398 397776 41426
rect 397656 41290 397684 41398
rect 397656 41262 397776 41290
rect 397644 40384 397696 40390
rect 397642 40352 397644 40361
rect 397696 40352 397698 40361
rect 397642 40287 397698 40296
rect 397748 22114 397776 41262
rect 397656 22086 397776 22114
rect 397656 12510 397684 22086
rect 398930 16824 398986 16833
rect 398930 16759 398986 16768
rect 398944 16561 398972 16759
rect 398930 16552 398986 16561
rect 398930 16487 398986 16496
rect 397644 12504 397696 12510
rect 397644 12446 397696 12452
rect 397552 12436 397604 12442
rect 397552 12378 397604 12384
rect 397564 7342 397592 12378
rect 397552 7336 397604 7342
rect 397552 7278 397604 7284
rect 397828 5432 397880 5438
rect 397828 5374 397880 5380
rect 397460 4412 397512 4418
rect 397460 4354 397512 4360
rect 396724 3868 396776 3874
rect 396724 3810 396776 3816
rect 395344 3800 395396 3806
rect 395344 3742 395396 3748
rect 396632 3392 396684 3398
rect 396632 3334 396684 3340
rect 395436 2848 395488 2854
rect 395436 2790 395488 2796
rect 395448 480 395476 2790
rect 396644 480 396672 3334
rect 397840 480 397868 5374
rect 399036 4350 399064 340054
rect 400232 338094 400260 340068
rect 400220 338088 400272 338094
rect 400220 338030 400272 338036
rect 400784 336938 400812 340068
rect 400876 340054 401442 340082
rect 401704 340054 402086 340082
rect 400772 336932 400824 336938
rect 400772 336874 400824 336880
rect 400876 335594 400904 340054
rect 401048 336796 401100 336802
rect 401048 336738 401100 336744
rect 400600 335566 400904 335594
rect 400600 321570 400628 335566
rect 401060 335458 401088 336738
rect 400876 335430 401088 335458
rect 400404 321564 400456 321570
rect 400404 321506 400456 321512
rect 400588 321564 400640 321570
rect 400588 321506 400640 321512
rect 400416 311930 400444 321506
rect 400324 311902 400444 311930
rect 400324 309194 400352 311902
rect 400312 309188 400364 309194
rect 400312 309130 400364 309136
rect 400404 309188 400456 309194
rect 400404 309130 400456 309136
rect 400416 302326 400444 309130
rect 400404 302320 400456 302326
rect 400404 302262 400456 302268
rect 400496 302116 400548 302122
rect 400496 302058 400548 302064
rect 400508 298110 400536 302058
rect 400496 298104 400548 298110
rect 400496 298046 400548 298052
rect 400588 298104 400640 298110
rect 400588 298046 400640 298052
rect 400600 280242 400628 298046
rect 400508 280214 400628 280242
rect 400508 280158 400536 280214
rect 400496 280152 400548 280158
rect 400496 280094 400548 280100
rect 400588 270564 400640 270570
rect 400588 270506 400640 270512
rect 400600 263514 400628 270506
rect 400508 263486 400628 263514
rect 400508 260846 400536 263486
rect 400496 260840 400548 260846
rect 400496 260782 400548 260788
rect 400588 251252 400640 251258
rect 400588 251194 400640 251200
rect 400600 244202 400628 251194
rect 400508 244174 400628 244202
rect 400508 241505 400536 244174
rect 400310 241496 400366 241505
rect 400310 241431 400366 241440
rect 400494 241496 400550 241505
rect 400494 241431 400550 241440
rect 400324 231878 400352 241431
rect 400312 231872 400364 231878
rect 400312 231814 400364 231820
rect 400588 231872 400640 231878
rect 400588 231814 400640 231820
rect 400600 224890 400628 231814
rect 400508 224862 400628 224890
rect 400508 222193 400536 224862
rect 400310 222184 400366 222193
rect 400310 222119 400366 222128
rect 400494 222184 400550 222193
rect 400494 222119 400550 222128
rect 400324 212566 400352 222119
rect 400312 212560 400364 212566
rect 400312 212502 400364 212508
rect 400588 212560 400640 212566
rect 400588 212502 400640 212508
rect 400600 205578 400628 212502
rect 400508 205550 400628 205578
rect 400508 202881 400536 205550
rect 400310 202872 400366 202881
rect 400310 202807 400366 202816
rect 400494 202872 400550 202881
rect 400494 202807 400550 202816
rect 400324 193254 400352 202807
rect 400312 193248 400364 193254
rect 400312 193190 400364 193196
rect 400588 193248 400640 193254
rect 400588 193190 400640 193196
rect 400600 186266 400628 193190
rect 400508 186238 400628 186266
rect 400508 176746 400536 186238
rect 400416 176718 400536 176746
rect 400416 176662 400444 176718
rect 400404 176656 400456 176662
rect 400404 176598 400456 176604
rect 400588 176656 400640 176662
rect 400588 176598 400640 176604
rect 400600 173890 400628 176598
rect 400416 173862 400628 173890
rect 400416 164286 400444 173862
rect 400312 164280 400364 164286
rect 400312 164222 400364 164228
rect 400404 164280 400456 164286
rect 400404 164222 400456 164228
rect 400324 154737 400352 164222
rect 400310 154728 400366 154737
rect 400310 154663 400366 154672
rect 400494 154592 400550 154601
rect 400494 154527 400550 154536
rect 400508 153202 400536 154527
rect 400496 153196 400548 153202
rect 400496 153138 400548 153144
rect 400496 147620 400548 147626
rect 400496 147562 400548 147568
rect 400508 143546 400536 147562
rect 400404 143540 400456 143546
rect 400404 143482 400456 143488
rect 400496 143540 400548 143546
rect 400496 143482 400548 143488
rect 400416 128382 400444 143482
rect 400404 128376 400456 128382
rect 400404 128318 400456 128324
rect 400496 128308 400548 128314
rect 400496 128250 400548 128256
rect 400508 124166 400536 128250
rect 400496 124160 400548 124166
rect 400496 124102 400548 124108
rect 400312 114572 400364 114578
rect 400312 114514 400364 114520
rect 400324 106321 400352 114514
rect 400310 106312 400366 106321
rect 400310 106247 400366 106256
rect 400494 106312 400550 106321
rect 400494 106247 400550 106256
rect 400508 101402 400536 106247
rect 400324 101374 400536 101402
rect 400324 96665 400352 101374
rect 400310 96656 400366 96665
rect 400310 96591 400366 96600
rect 400586 96656 400642 96665
rect 400586 96591 400642 96600
rect 400600 89706 400628 96591
rect 400416 89678 400628 89706
rect 400416 86970 400444 89678
rect 400404 86964 400456 86970
rect 400404 86906 400456 86912
rect 400312 77308 400364 77314
rect 400312 77250 400364 77256
rect 400324 70394 400352 77250
rect 400324 70366 400536 70394
rect 400508 51202 400536 70366
rect 400496 51196 400548 51202
rect 400496 51138 400548 51144
rect 400404 48408 400456 48414
rect 400404 48350 400456 48356
rect 400416 48278 400444 48350
rect 400404 48272 400456 48278
rect 400404 48214 400456 48220
rect 400772 48272 400824 48278
rect 400772 48214 400824 48220
rect 400784 38706 400812 48214
rect 400692 38678 400812 38706
rect 400692 31822 400720 38678
rect 400680 31816 400732 31822
rect 400680 31758 400732 31764
rect 400680 29096 400732 29102
rect 400600 29044 400680 29050
rect 400600 29038 400732 29044
rect 400600 29022 400720 29038
rect 400600 27606 400628 29022
rect 400588 27600 400640 27606
rect 400588 27542 400640 27548
rect 400588 18012 400640 18018
rect 400588 17954 400640 17960
rect 400600 17882 400628 17954
rect 400588 17876 400640 17882
rect 400588 17818 400640 17824
rect 400404 8356 400456 8362
rect 400404 8298 400456 8304
rect 399024 4344 399076 4350
rect 399024 4286 399076 4292
rect 400416 4282 400444 8298
rect 400404 4276 400456 4282
rect 400404 4218 400456 4224
rect 400220 4140 400272 4146
rect 400220 4082 400272 4088
rect 399024 3800 399076 3806
rect 399024 3742 399076 3748
rect 399036 480 399064 3742
rect 400232 480 400260 4082
rect 400876 3942 400904 335430
rect 401704 8974 401732 340054
rect 402624 338026 402652 340068
rect 403084 340054 403282 340082
rect 402612 338020 402664 338026
rect 402612 337962 402664 337968
rect 401692 8968 401744 8974
rect 401692 8910 401744 8916
rect 401324 5500 401376 5506
rect 401324 5442 401376 5448
rect 400864 3936 400916 3942
rect 400864 3878 400916 3884
rect 401336 480 401364 5442
rect 403084 4214 403112 340054
rect 403912 337346 403940 340068
rect 403900 337340 403952 337346
rect 403900 337282 403952 337288
rect 404464 336870 404492 340068
rect 404556 340054 405122 340082
rect 405766 340054 405872 340082
rect 404452 336864 404504 336870
rect 404452 336806 404504 336812
rect 404556 4758 404584 340054
rect 405004 338088 405056 338094
rect 405004 338030 405056 338036
rect 404544 4752 404596 4758
rect 404544 4694 404596 4700
rect 404912 4752 404964 4758
rect 404912 4694 404964 4700
rect 403072 4208 403124 4214
rect 403072 4150 403124 4156
rect 403532 4072 403584 4078
rect 403584 4020 403664 4026
rect 403532 4014 403664 4020
rect 403544 3998 403664 4014
rect 402520 3460 402572 3466
rect 402520 3402 402572 3408
rect 402532 480 402560 3402
rect 403636 3126 403664 3998
rect 403716 3868 403768 3874
rect 403716 3810 403768 3816
rect 403624 3120 403676 3126
rect 403624 3062 403676 3068
rect 403728 480 403756 3810
rect 404924 480 404952 4694
rect 405016 4214 405044 338030
rect 405648 40384 405700 40390
rect 405646 40352 405648 40361
rect 405700 40352 405702 40361
rect 405646 40287 405702 40296
rect 405844 7614 405872 340054
rect 406304 337822 406332 340068
rect 406672 340054 406962 340082
rect 406292 337816 406344 337822
rect 406292 337758 406344 337764
rect 406672 335646 406700 340054
rect 407500 337278 407528 340068
rect 407764 337952 407816 337958
rect 407764 337894 407816 337900
rect 407488 337272 407540 337278
rect 407488 337214 407540 337220
rect 405924 335640 405976 335646
rect 405924 335582 405976 335588
rect 406660 335640 406712 335646
rect 406660 335582 406712 335588
rect 405832 7608 405884 7614
rect 405832 7550 405884 7556
rect 405936 4690 405964 335582
rect 407776 4876 407804 337894
rect 408144 336802 408172 340068
rect 408512 340054 408802 340082
rect 408132 336796 408184 336802
rect 408132 336738 408184 336744
rect 408408 16856 408460 16862
rect 408406 16824 408408 16833
rect 408460 16824 408462 16833
rect 408406 16759 408462 16768
rect 408512 4894 408540 340054
rect 408880 331242 408908 340190
rect 409788 337816 409840 337822
rect 409788 337758 409840 337764
rect 409144 337340 409196 337346
rect 409144 337282 409196 337288
rect 408696 331214 408908 331242
rect 408696 321638 408724 331214
rect 408684 321632 408736 321638
rect 408684 321574 408736 321580
rect 408776 321496 408828 321502
rect 408776 321438 408828 321444
rect 408788 312066 408816 321438
rect 408788 312038 408908 312066
rect 408880 307850 408908 312038
rect 408788 307822 408908 307850
rect 408788 302258 408816 307822
rect 408776 302252 408828 302258
rect 408776 302194 408828 302200
rect 408776 298172 408828 298178
rect 408776 298114 408828 298120
rect 408788 293078 408816 298114
rect 408776 293072 408828 293078
rect 408776 293014 408828 293020
rect 408776 282804 408828 282810
rect 408776 282746 408828 282752
rect 408788 278730 408816 282746
rect 408776 278724 408828 278730
rect 408776 278666 408828 278672
rect 408776 263492 408828 263498
rect 408776 263434 408828 263440
rect 408788 259457 408816 263434
rect 408774 259448 408830 259457
rect 408774 259383 408830 259392
rect 408958 259448 409014 259457
rect 408958 259383 409014 259392
rect 408972 244186 409000 259383
rect 408776 244180 408828 244186
rect 408776 244122 408828 244128
rect 408960 244180 409012 244186
rect 408960 244122 409012 244128
rect 408788 234734 408816 244122
rect 408776 234728 408828 234734
rect 408776 234670 408828 234676
rect 408684 234592 408736 234598
rect 408684 234534 408736 234540
rect 408696 231810 408724 234534
rect 408684 231804 408736 231810
rect 408684 231746 408736 231752
rect 408776 222216 408828 222222
rect 408776 222158 408828 222164
rect 408788 215422 408816 222158
rect 408776 215416 408828 215422
rect 408776 215358 408828 215364
rect 408684 215280 408736 215286
rect 408684 215222 408736 215228
rect 408696 212498 408724 215222
rect 408684 212492 408736 212498
rect 408684 212434 408736 212440
rect 408776 202904 408828 202910
rect 408776 202846 408828 202852
rect 408788 196110 408816 202846
rect 408776 196104 408828 196110
rect 408776 196046 408828 196052
rect 408684 195968 408736 195974
rect 408684 195910 408736 195916
rect 408696 193225 408724 195910
rect 408682 193216 408738 193225
rect 408682 193151 408738 193160
rect 408958 193216 409014 193225
rect 408958 193151 409014 193160
rect 408972 183598 409000 193151
rect 408776 183592 408828 183598
rect 408776 183534 408828 183540
rect 408960 183592 409012 183598
rect 408960 183534 409012 183540
rect 408788 176798 408816 183534
rect 408776 176792 408828 176798
rect 408776 176734 408828 176740
rect 408776 176588 408828 176594
rect 408776 176530 408828 176536
rect 408788 166954 408816 176530
rect 408604 166926 408816 166954
rect 408604 157418 408632 166926
rect 408592 157412 408644 157418
rect 408592 157354 408644 157360
rect 408684 157276 408736 157282
rect 408684 157218 408736 157224
rect 408696 154562 408724 157218
rect 408684 154556 408736 154562
rect 408684 154498 408736 154504
rect 408684 147620 408736 147626
rect 408684 147562 408736 147568
rect 408696 144922 408724 147562
rect 408696 144894 408816 144922
rect 408788 138106 408816 144894
rect 408776 138100 408828 138106
rect 408776 138042 408828 138048
rect 408684 137964 408736 137970
rect 408684 137906 408736 137912
rect 408696 135250 408724 137906
rect 408684 135244 408736 135250
rect 408684 135186 408736 135192
rect 408684 128308 408736 128314
rect 408684 128250 408736 128256
rect 408696 125610 408724 128250
rect 408696 125582 408816 125610
rect 408788 118794 408816 125582
rect 408776 118788 408828 118794
rect 408776 118730 408828 118736
rect 408684 118652 408736 118658
rect 408684 118594 408736 118600
rect 408696 109070 408724 118594
rect 408684 109064 408736 109070
rect 408684 109006 408736 109012
rect 408776 108996 408828 109002
rect 408776 108938 408828 108944
rect 408788 104854 408816 108938
rect 408776 104848 408828 104854
rect 408776 104790 408828 104796
rect 408684 95260 408736 95266
rect 408684 95202 408736 95208
rect 408696 89758 408724 95202
rect 408684 89752 408736 89758
rect 408684 89694 408736 89700
rect 408776 89616 408828 89622
rect 408776 89558 408828 89564
rect 408788 82142 408816 89558
rect 408776 82136 408828 82142
rect 408776 82078 408828 82084
rect 408776 77308 408828 77314
rect 408776 77250 408828 77256
rect 408788 70446 408816 77250
rect 408776 70440 408828 70446
rect 408776 70382 408828 70388
rect 408776 67652 408828 67658
rect 408776 67594 408828 67600
rect 408788 62830 408816 67594
rect 408776 62824 408828 62830
rect 408776 62766 408828 62772
rect 408776 57996 408828 58002
rect 408776 57938 408828 57944
rect 408788 51202 408816 57938
rect 408776 51196 408828 51202
rect 408776 51138 408828 51144
rect 408684 48408 408736 48414
rect 408736 48356 408816 48362
rect 408684 48350 408816 48356
rect 408696 48334 408816 48350
rect 408788 46918 408816 48334
rect 408776 46912 408828 46918
rect 408776 46854 408828 46860
rect 408868 38548 408920 38554
rect 408868 38490 408920 38496
rect 408880 31634 408908 38490
rect 408788 31606 408908 31634
rect 408788 22166 408816 31606
rect 408776 22160 408828 22166
rect 408776 22102 408828 22108
rect 408684 22092 408736 22098
rect 408684 22034 408736 22040
rect 408696 12458 408724 22034
rect 408696 12430 408816 12458
rect 408788 6866 408816 12430
rect 408776 6860 408828 6866
rect 408776 6802 408828 6808
rect 407408 4848 407804 4876
rect 408500 4888 408552 4894
rect 405924 4684 405976 4690
rect 405924 4626 405976 4632
rect 405004 4208 405056 4214
rect 405004 4150 405056 4156
rect 407408 3448 407436 4848
rect 408500 4830 408552 4836
rect 408684 4276 408736 4282
rect 408684 4218 408736 4224
rect 408592 4208 408644 4214
rect 408512 4156 408592 4162
rect 408512 4150 408644 4156
rect 408408 4140 408460 4146
rect 408408 4082 408460 4088
rect 408512 4134 408632 4150
rect 408420 3913 408448 4082
rect 408406 3904 408462 3913
rect 408406 3839 408462 3848
rect 408512 3670 408540 4134
rect 408696 4010 408724 4218
rect 409156 4078 409184 337282
rect 409144 4072 409196 4078
rect 409144 4014 409196 4020
rect 408684 4004 408736 4010
rect 408684 3946 408736 3952
rect 408592 3936 408644 3942
rect 408590 3904 408592 3913
rect 408644 3904 408646 3913
rect 408590 3839 408646 3848
rect 408316 3664 408368 3670
rect 408314 3632 408316 3641
rect 408500 3664 408552 3670
rect 408368 3632 408370 3641
rect 408592 3664 408644 3670
rect 408500 3606 408552 3612
rect 408590 3632 408592 3641
rect 408644 3632 408646 3641
rect 408314 3567 408370 3576
rect 408590 3567 408646 3576
rect 409800 3466 409828 337758
rect 409984 337754 410012 340068
rect 410076 340054 410642 340082
rect 409972 337748 410024 337754
rect 409972 337690 410024 337696
rect 410076 4826 410104 340054
rect 411180 337210 411208 340068
rect 411824 338094 411852 340068
rect 411916 340054 412482 340082
rect 411812 338088 411864 338094
rect 411812 338030 411864 338036
rect 411168 337204 411220 337210
rect 411168 337146 411220 337152
rect 410524 337000 410576 337006
rect 410524 336942 410576 336948
rect 410064 4820 410116 4826
rect 410064 4762 410116 4768
rect 410536 4146 410564 336942
rect 410616 336796 410668 336802
rect 410616 336738 410668 336744
rect 410524 4140 410576 4146
rect 410524 4082 410576 4088
rect 407132 3420 407436 3448
rect 408500 3460 408552 3466
rect 407132 3330 407160 3420
rect 408500 3402 408552 3408
rect 409788 3460 409840 3466
rect 409788 3402 409840 3408
rect 407120 3324 407172 3330
rect 407120 3266 407172 3272
rect 407304 3324 407356 3330
rect 407304 3266 407356 3272
rect 406108 2984 406160 2990
rect 406108 2926 406160 2932
rect 406120 480 406148 2926
rect 407316 480 407344 3266
rect 408512 480 408540 3402
rect 410628 3369 410656 336738
rect 411916 335594 411944 340054
rect 412088 338088 412140 338094
rect 412088 338030 412140 338036
rect 411364 335566 411944 335594
rect 410706 17096 410762 17105
rect 410706 17031 410762 17040
rect 410720 16862 410748 17031
rect 410708 16856 410760 16862
rect 410708 16798 410760 16804
rect 411364 6050 411392 335566
rect 412100 331242 412128 338030
rect 412548 337748 412600 337754
rect 412548 337690 412600 337696
rect 411916 331214 412128 331242
rect 411352 6044 411404 6050
rect 411352 5986 411404 5992
rect 411916 4146 411944 331214
rect 412560 4146 412588 337690
rect 413020 336802 413048 340068
rect 413468 337476 413520 337482
rect 413468 337418 413520 337424
rect 413376 337272 413428 337278
rect 413376 337214 413428 337220
rect 413284 336864 413336 336870
rect 413284 336806 413336 336812
rect 413008 336796 413060 336802
rect 413008 336738 413060 336744
rect 411904 4140 411956 4146
rect 411904 4082 411956 4088
rect 412088 4140 412140 4146
rect 412088 4082 412140 4088
rect 412548 4140 412600 4146
rect 412548 4082 412600 4088
rect 410892 4072 410944 4078
rect 410892 4014 410944 4020
rect 410614 3360 410670 3369
rect 409696 3324 409748 3330
rect 410614 3295 410670 3304
rect 409696 3266 409748 3272
rect 409144 2984 409196 2990
rect 409420 2984 409472 2990
rect 409196 2932 409420 2938
rect 409144 2926 409472 2932
rect 409156 2910 409460 2926
rect 409708 480 409736 3266
rect 410904 480 410932 4014
rect 412100 480 412128 4082
rect 413296 4078 413324 336806
rect 413284 4072 413336 4078
rect 413284 4014 413336 4020
rect 412640 3460 412692 3466
rect 412640 3402 412692 3408
rect 412652 3058 412680 3402
rect 413388 3262 413416 337214
rect 413480 3466 413508 337418
rect 413664 337142 413692 340068
rect 414124 340054 414322 340082
rect 413652 337136 413704 337142
rect 413652 337078 413704 337084
rect 414124 4962 414152 340054
rect 414664 337136 414716 337142
rect 414664 337078 414716 337084
rect 414112 4956 414164 4962
rect 414112 4898 414164 4904
rect 414480 4140 414532 4146
rect 414480 4082 414532 4088
rect 413468 3460 413520 3466
rect 413468 3402 413520 3408
rect 413376 3256 413428 3262
rect 413376 3198 413428 3204
rect 412640 3052 412692 3058
rect 412640 2994 412692 3000
rect 413284 604 413336 610
rect 413284 546 413336 552
rect 413296 480 413324 546
rect 414492 480 414520 4082
rect 414676 3126 414704 337078
rect 414860 337074 414888 340068
rect 415504 337958 415532 340068
rect 415596 340054 416162 340082
rect 416424 340054 416714 340082
rect 415492 337952 415544 337958
rect 415492 337894 415544 337900
rect 414848 337068 414900 337074
rect 414848 337010 414900 337016
rect 415306 134328 415362 134337
rect 415306 134263 415362 134272
rect 415320 134201 415348 134263
rect 415306 134192 415362 134201
rect 415306 134127 415362 134136
rect 415596 5914 415624 340054
rect 416044 337952 416096 337958
rect 416044 337894 416096 337900
rect 415584 5908 415636 5914
rect 415584 5850 415636 5856
rect 416056 4146 416084 337894
rect 416424 337006 416452 340054
rect 416688 338020 416740 338026
rect 416688 337962 416740 337968
rect 416412 337000 416464 337006
rect 416412 336942 416464 336948
rect 416136 336796 416188 336802
rect 416136 336738 416188 336744
rect 416044 4140 416096 4146
rect 416044 4082 416096 4088
rect 414664 3120 414716 3126
rect 414664 3062 414716 3068
rect 415676 3120 415728 3126
rect 415676 3062 415728 3068
rect 415688 480 415716 3062
rect 416148 2938 416176 336738
rect 416700 3126 416728 337962
rect 417344 337210 417372 340068
rect 417436 340054 418002 340082
rect 417332 337204 417384 337210
rect 417332 337146 417384 337152
rect 417436 335594 417464 340054
rect 418540 337686 418568 340068
rect 419184 338094 419212 340068
rect 419644 340054 419842 340082
rect 419172 338088 419224 338094
rect 419172 338030 419224 338036
rect 418528 337680 418580 337686
rect 418528 337622 418580 337628
rect 417608 337204 417660 337210
rect 417608 337146 417660 337152
rect 416792 335566 417464 335594
rect 416792 331226 416820 335566
rect 417620 334234 417648 337146
rect 417436 334206 417648 334234
rect 416780 331220 416832 331226
rect 416780 331162 416832 331168
rect 416964 331220 417016 331226
rect 416964 331162 417016 331168
rect 416976 328438 417004 331162
rect 416964 328432 417016 328438
rect 416964 328374 417016 328380
rect 416872 318844 416924 318850
rect 416872 318786 416924 318792
rect 416884 311930 416912 318786
rect 416792 311902 416912 311930
rect 416792 311846 416820 311902
rect 416780 311840 416832 311846
rect 416780 311782 416832 311788
rect 416964 311840 417016 311846
rect 416964 311782 417016 311788
rect 416976 309126 417004 311782
rect 416964 309120 417016 309126
rect 416964 309062 417016 309068
rect 416872 299532 416924 299538
rect 416872 299474 416924 299480
rect 416884 294658 416912 299474
rect 416884 294630 417004 294658
rect 416976 282826 417004 294630
rect 416884 282798 417004 282826
rect 416884 280158 416912 282798
rect 416872 280152 416924 280158
rect 416872 280094 416924 280100
rect 416964 270564 417016 270570
rect 416964 270506 417016 270512
rect 416976 263514 417004 270506
rect 416884 263486 417004 263514
rect 416884 260846 416912 263486
rect 416872 260840 416924 260846
rect 416872 260782 416924 260788
rect 416964 251252 417016 251258
rect 416964 251194 417016 251200
rect 416976 244202 417004 251194
rect 416884 244174 417004 244202
rect 416884 241505 416912 244174
rect 416870 241496 416926 241505
rect 416870 241431 416926 241440
rect 417146 241496 417202 241505
rect 417146 241431 417202 241440
rect 417160 231878 417188 241431
rect 416964 231872 417016 231878
rect 416964 231814 417016 231820
rect 417148 231872 417200 231878
rect 417148 231814 417200 231820
rect 416976 224890 417004 231814
rect 416884 224862 417004 224890
rect 416884 222193 416912 224862
rect 416870 222184 416926 222193
rect 416870 222119 416926 222128
rect 417146 222184 417202 222193
rect 417146 222119 417202 222128
rect 417160 212566 417188 222119
rect 416964 212560 417016 212566
rect 416964 212502 417016 212508
rect 417148 212560 417200 212566
rect 417148 212502 417200 212508
rect 416976 205578 417004 212502
rect 416884 205550 417004 205578
rect 416884 202881 416912 205550
rect 416870 202872 416926 202881
rect 416870 202807 416926 202816
rect 417146 202872 417202 202881
rect 417146 202807 417202 202816
rect 417160 193254 417188 202807
rect 416964 193248 417016 193254
rect 416964 193190 417016 193196
rect 417148 193248 417200 193254
rect 417148 193190 417200 193196
rect 416976 186266 417004 193190
rect 416884 186238 417004 186266
rect 416884 183569 416912 186238
rect 416870 183560 416926 183569
rect 416870 183495 416926 183504
rect 417146 183560 417202 183569
rect 417146 183495 417202 183504
rect 417160 173942 417188 183495
rect 416964 173936 417016 173942
rect 416964 173878 417016 173884
rect 417148 173936 417200 173942
rect 417148 173878 417200 173884
rect 416976 166954 417004 173878
rect 416884 166926 417004 166954
rect 416884 164218 416912 166926
rect 416872 164212 416924 164218
rect 416872 164154 416924 164160
rect 417148 164212 417200 164218
rect 417148 164154 417200 164160
rect 417160 154601 417188 164154
rect 416962 154592 417018 154601
rect 416962 154527 417018 154536
rect 417146 154592 417202 154601
rect 417146 154527 417202 154536
rect 416976 147642 417004 154527
rect 416884 147614 417004 147642
rect 416884 138038 416912 147614
rect 416872 138032 416924 138038
rect 416872 137974 416924 137980
rect 416780 137964 416832 137970
rect 416780 137906 416832 137912
rect 416792 135289 416820 137906
rect 416778 135280 416834 135289
rect 416778 135215 416834 135224
rect 416962 135280 417018 135289
rect 416962 135215 417018 135224
rect 416976 128330 417004 135215
rect 416884 128302 417004 128330
rect 416884 118726 416912 128302
rect 416872 118720 416924 118726
rect 416872 118662 416924 118668
rect 416780 118652 416832 118658
rect 416780 118594 416832 118600
rect 416792 115977 416820 118594
rect 416778 115968 416834 115977
rect 416778 115903 416834 115912
rect 416962 115968 417018 115977
rect 416962 115903 417018 115912
rect 416976 109018 417004 115903
rect 416884 108990 417004 109018
rect 416884 99414 416912 108990
rect 416872 99408 416924 99414
rect 416872 99350 416924 99356
rect 416780 99340 416832 99346
rect 416780 99282 416832 99288
rect 416792 96665 416820 99282
rect 416778 96656 416834 96665
rect 416778 96591 416834 96600
rect 416962 96656 417018 96665
rect 416962 96591 417018 96600
rect 416976 89706 417004 96591
rect 416884 89678 417004 89706
rect 416884 82090 416912 89678
rect 416792 82062 416912 82090
rect 416792 77382 416820 82062
rect 416780 77376 416832 77382
rect 416780 77318 416832 77324
rect 416964 77376 417016 77382
rect 416964 77318 417016 77324
rect 416976 77246 417004 77318
rect 416964 77240 417016 77246
rect 416964 77182 417016 77188
rect 416872 67652 416924 67658
rect 416872 67594 416924 67600
rect 416884 60738 416912 67594
rect 416792 60722 416912 60738
rect 416780 60716 416912 60722
rect 416832 60710 416912 60716
rect 416964 60716 417016 60722
rect 416780 60658 416832 60664
rect 416964 60658 417016 60664
rect 416976 57934 417004 60658
rect 416964 57928 417016 57934
rect 416964 57870 417016 57876
rect 416872 48408 416924 48414
rect 416872 48350 416924 48356
rect 416884 48278 416912 48350
rect 416872 48272 416924 48278
rect 416872 48214 416924 48220
rect 417056 48272 417108 48278
rect 417056 48214 417108 48220
rect 417068 38706 417096 48214
rect 416976 38678 417096 38706
rect 416976 38622 417004 38678
rect 416964 38616 417016 38622
rect 416964 38558 417016 38564
rect 416872 29028 416924 29034
rect 416872 28970 416924 28976
rect 416884 22114 416912 28970
rect 416792 22098 416912 22114
rect 416780 22092 416912 22098
rect 416832 22086 416912 22092
rect 416964 22092 417016 22098
rect 416780 22034 416832 22040
rect 416964 22034 417016 22040
rect 416976 19310 417004 22034
rect 416964 19304 417016 19310
rect 416964 19246 417016 19252
rect 416964 12300 417016 12306
rect 416964 12242 417016 12248
rect 416976 5030 417004 12242
rect 416964 5024 417016 5030
rect 416964 4966 417016 4972
rect 417436 3398 417464 334206
rect 418066 169960 418122 169969
rect 418066 169895 418122 169904
rect 418080 169561 418108 169895
rect 418066 169552 418122 169561
rect 418066 169487 418122 169496
rect 418066 40352 418122 40361
rect 418066 40287 418122 40296
rect 418080 40202 418108 40287
rect 418158 40216 418214 40225
rect 418080 40174 418158 40202
rect 418158 40151 418214 40160
rect 418066 17096 418122 17105
rect 418066 17031 418122 17040
rect 418080 16946 418108 17031
rect 418250 16960 418306 16969
rect 418080 16918 418250 16946
rect 418250 16895 418306 16904
rect 419644 5846 419672 340054
rect 420380 337482 420408 340068
rect 420828 337680 420880 337686
rect 420828 337622 420880 337628
rect 420368 337476 420420 337482
rect 420368 337418 420420 337424
rect 420276 337068 420328 337074
rect 420276 337010 420328 337016
rect 420184 337000 420236 337006
rect 420184 336942 420236 336948
rect 419632 5840 419684 5846
rect 419632 5782 419684 5788
rect 420196 4146 420224 336942
rect 419172 4140 419224 4146
rect 419172 4082 419224 4088
rect 420184 4140 420236 4146
rect 420184 4082 420236 4088
rect 417424 3392 417476 3398
rect 417424 3334 417476 3340
rect 417976 3392 418028 3398
rect 417976 3334 418028 3340
rect 416872 3256 416924 3262
rect 416872 3198 416924 3204
rect 416688 3120 416740 3126
rect 416688 3062 416740 3068
rect 416056 2922 416176 2938
rect 416044 2916 416176 2922
rect 416096 2910 416176 2916
rect 416044 2858 416096 2864
rect 416884 480 416912 3198
rect 417988 480 418016 3334
rect 419184 480 419212 4082
rect 420288 4010 420316 337010
rect 420840 4146 420868 337622
rect 421024 337414 421052 340068
rect 421116 340054 421682 340082
rect 421944 340054 422234 340082
rect 421012 337408 421064 337414
rect 421012 337350 421064 337356
rect 421116 6186 421144 340054
rect 421944 336938 421972 340054
rect 422208 337272 422260 337278
rect 422208 337214 422260 337220
rect 421932 336932 421984 336938
rect 421932 336874 421984 336880
rect 422114 27568 422170 27577
rect 422114 27503 422170 27512
rect 422128 19242 422156 27503
rect 422116 19236 422168 19242
rect 422116 19178 422168 19184
rect 421104 6180 421156 6186
rect 421104 6122 421156 6128
rect 420368 4140 420420 4146
rect 420368 4082 420420 4088
rect 420828 4140 420880 4146
rect 420828 4082 420880 4088
rect 420276 4004 420328 4010
rect 420276 3946 420328 3952
rect 420380 480 420408 4082
rect 422220 2922 422248 337214
rect 422864 337142 422892 340068
rect 423232 340054 423522 340082
rect 422852 337136 422904 337142
rect 422852 337078 422904 337084
rect 423232 335646 423260 340054
rect 424060 337210 424088 340068
rect 424048 337204 424100 337210
rect 424048 337146 424100 337152
rect 423588 337136 423640 337142
rect 423588 337078 423640 337084
rect 422300 335640 422352 335646
rect 422300 335582 422352 335588
rect 423220 335640 423272 335646
rect 423220 335582 423272 335588
rect 422312 331226 422340 335582
rect 422300 331220 422352 331226
rect 422300 331162 422352 331168
rect 422484 331220 422536 331226
rect 422484 331162 422536 331168
rect 422496 328438 422524 331162
rect 422484 328432 422536 328438
rect 422484 328374 422536 328380
rect 422392 318844 422444 318850
rect 422392 318786 422444 318792
rect 422404 311930 422432 318786
rect 422312 311902 422432 311930
rect 422312 311846 422340 311902
rect 422300 311840 422352 311846
rect 422300 311782 422352 311788
rect 422484 311840 422536 311846
rect 422484 311782 422536 311788
rect 422496 309126 422524 311782
rect 422484 309120 422536 309126
rect 422484 309062 422536 309068
rect 422484 299940 422536 299946
rect 422484 299882 422536 299888
rect 422496 282946 422524 299882
rect 422300 282940 422352 282946
rect 422300 282882 422352 282888
rect 422484 282940 422536 282946
rect 422484 282882 422536 282888
rect 422312 282826 422340 282882
rect 422312 282798 422432 282826
rect 422404 273306 422432 282798
rect 422404 273278 422524 273306
rect 422496 263634 422524 273278
rect 422300 263628 422352 263634
rect 422300 263570 422352 263576
rect 422484 263628 422536 263634
rect 422484 263570 422536 263576
rect 422312 263514 422340 263570
rect 422312 263486 422432 263514
rect 422404 253994 422432 263486
rect 422404 253966 422524 253994
rect 422496 244322 422524 253966
rect 422300 244316 422352 244322
rect 422300 244258 422352 244264
rect 422484 244316 422536 244322
rect 422484 244258 422536 244264
rect 422312 244202 422340 244258
rect 422312 244174 422432 244202
rect 422404 234682 422432 244174
rect 422404 234654 422524 234682
rect 422496 225010 422524 234654
rect 422300 225004 422352 225010
rect 422300 224946 422352 224952
rect 422484 225004 422536 225010
rect 422484 224946 422536 224952
rect 422312 224890 422340 224946
rect 422312 224862 422432 224890
rect 422404 215370 422432 224862
rect 422404 215342 422524 215370
rect 422496 205698 422524 215342
rect 422300 205692 422352 205698
rect 422300 205634 422352 205640
rect 422484 205692 422536 205698
rect 422484 205634 422536 205640
rect 422312 205578 422340 205634
rect 422312 205550 422432 205578
rect 422404 196058 422432 205550
rect 422404 196030 422524 196058
rect 422496 186386 422524 196030
rect 422300 186380 422352 186386
rect 422300 186322 422352 186328
rect 422484 186380 422536 186386
rect 422484 186322 422536 186328
rect 422312 186266 422340 186322
rect 422312 186238 422432 186266
rect 422404 183569 422432 186238
rect 422390 183560 422446 183569
rect 422390 183495 422446 183504
rect 422666 183560 422722 183569
rect 422666 183495 422722 183504
rect 422680 173942 422708 183495
rect 422484 173936 422536 173942
rect 422484 173878 422536 173884
rect 422668 173936 422720 173942
rect 422668 173878 422720 173884
rect 422496 167074 422524 173878
rect 422300 167068 422352 167074
rect 422300 167010 422352 167016
rect 422484 167068 422536 167074
rect 422484 167010 422536 167016
rect 422312 166954 422340 167010
rect 422312 166926 422432 166954
rect 422404 164218 422432 166926
rect 422392 164212 422444 164218
rect 422392 164154 422444 164160
rect 422392 157344 422444 157350
rect 422392 157286 422444 157292
rect 422404 154578 422432 157286
rect 422404 154550 422524 154578
rect 422496 147694 422524 154550
rect 422300 147688 422352 147694
rect 422484 147688 422536 147694
rect 422352 147636 422432 147642
rect 422300 147630 422432 147636
rect 422484 147630 422536 147636
rect 422312 147614 422432 147630
rect 422404 144906 422432 147614
rect 422392 144900 422444 144906
rect 422392 144842 422444 144848
rect 422392 137964 422444 137970
rect 422392 137906 422444 137912
rect 422404 135266 422432 137906
rect 422404 135238 422524 135266
rect 422496 128382 422524 135238
rect 422300 128376 422352 128382
rect 422484 128376 422536 128382
rect 422352 128324 422432 128330
rect 422300 128318 422432 128324
rect 422484 128318 422536 128324
rect 422312 128302 422432 128318
rect 422404 125594 422432 128302
rect 422392 125588 422444 125594
rect 422392 125530 422444 125536
rect 422392 118652 422444 118658
rect 422392 118594 422444 118600
rect 422404 115954 422432 118594
rect 422404 115926 422524 115954
rect 422496 109070 422524 115926
rect 422300 109064 422352 109070
rect 422484 109064 422536 109070
rect 422352 109012 422432 109018
rect 422300 109006 422432 109012
rect 422484 109006 422536 109012
rect 422312 108990 422432 109006
rect 422404 106282 422432 108990
rect 422392 106276 422444 106282
rect 422392 106218 422444 106224
rect 422392 99340 422444 99346
rect 422392 99282 422444 99288
rect 422404 96642 422432 99282
rect 422404 96614 422524 96642
rect 422496 89758 422524 96614
rect 422300 89752 422352 89758
rect 422484 89752 422536 89758
rect 422352 89700 422432 89706
rect 422300 89694 422432 89700
rect 422484 89694 422536 89700
rect 422312 89678 422432 89694
rect 422404 86970 422432 89678
rect 422392 86964 422444 86970
rect 422392 86906 422444 86912
rect 422484 77308 422536 77314
rect 422484 77250 422536 77256
rect 422496 70258 422524 77250
rect 422404 70230 422524 70258
rect 422404 60738 422432 70230
rect 422404 60710 422524 60738
rect 422496 48346 422524 60710
rect 422392 48340 422444 48346
rect 422392 48282 422444 48288
rect 422484 48340 422536 48346
rect 422484 48282 422536 48288
rect 422404 41426 422432 48282
rect 422404 41398 422524 41426
rect 422496 38622 422524 41398
rect 422484 38616 422536 38622
rect 422484 38558 422536 38564
rect 422392 27668 422444 27674
rect 422392 27610 422444 27616
rect 422298 27568 422354 27577
rect 422404 27554 422432 27610
rect 422354 27526 422432 27554
rect 422298 27503 422354 27512
rect 422484 19236 422536 19242
rect 422484 19178 422536 19184
rect 422496 9722 422524 19178
rect 422300 9716 422352 9722
rect 422300 9658 422352 9664
rect 422484 9716 422536 9722
rect 422484 9658 422536 9664
rect 422312 5098 422340 9658
rect 422300 5092 422352 5098
rect 422300 5034 422352 5040
rect 423600 4146 423628 337078
rect 424416 337000 424468 337006
rect 424416 336942 424468 336948
rect 424324 336796 424376 336802
rect 424324 336738 424376 336744
rect 422760 4140 422812 4146
rect 422760 4082 422812 4088
rect 423588 4140 423640 4146
rect 423588 4082 423640 4088
rect 423956 4140 424008 4146
rect 423956 4082 424008 4088
rect 421564 2916 421616 2922
rect 421564 2858 421616 2864
rect 422208 2916 422260 2922
rect 422208 2858 422260 2864
rect 421576 480 421604 2858
rect 422772 480 422800 4082
rect 423968 480 423996 4082
rect 424336 3126 424364 336738
rect 424428 4010 424456 336942
rect 424704 336870 424732 340068
rect 425164 340054 425270 340082
rect 424968 337272 425020 337278
rect 424968 337214 425020 337220
rect 424692 336864 424744 336870
rect 424692 336806 424744 336812
rect 424980 4146 425008 337214
rect 425060 169856 425112 169862
rect 425058 169824 425060 169833
rect 425112 169824 425114 169833
rect 425058 169759 425114 169768
rect 425164 6254 425192 340054
rect 425900 336802 425928 340068
rect 426558 340054 426664 340082
rect 425888 336796 425940 336802
rect 425888 336738 425940 336744
rect 425152 6248 425204 6254
rect 425152 6190 425204 6196
rect 424968 4140 425020 4146
rect 424968 4082 425020 4088
rect 424416 4004 424468 4010
rect 424416 3946 424468 3952
rect 425152 3936 425204 3942
rect 425152 3878 425204 3884
rect 424324 3120 424376 3126
rect 424324 3062 424376 3068
rect 425164 480 425192 3878
rect 426348 3528 426400 3534
rect 426348 3470 426400 3476
rect 426360 480 426388 3470
rect 426636 2990 426664 340054
rect 426728 340054 427110 340082
rect 427464 340054 427754 340082
rect 426728 5166 426756 340054
rect 427464 338094 427492 340054
rect 427452 338088 427504 338094
rect 427452 338030 427504 338036
rect 428384 337346 428412 340068
rect 428476 340054 428950 340082
rect 428372 337340 428424 337346
rect 428372 337282 428424 337288
rect 427084 336932 427136 336938
rect 427084 336874 427136 336880
rect 426716 5160 426768 5166
rect 426716 5102 426768 5108
rect 427096 3058 427124 336874
rect 428476 331378 428504 340054
rect 429108 337544 429160 337550
rect 429108 337486 429160 337492
rect 428556 337340 428608 337346
rect 428556 337282 428608 337288
rect 428384 331350 428504 331378
rect 428384 328681 428412 331350
rect 428568 331242 428596 337282
rect 428476 331214 428596 331242
rect 428370 328672 428426 328681
rect 428370 328607 428426 328616
rect 428002 328536 428058 328545
rect 428002 328471 428058 328480
rect 428016 328438 428044 328471
rect 428004 328432 428056 328438
rect 428004 328374 428056 328380
rect 427912 318844 427964 318850
rect 427912 318786 427964 318792
rect 427924 311930 427952 318786
rect 427832 311902 427952 311930
rect 427832 311846 427860 311902
rect 427820 311840 427872 311846
rect 427820 311782 427872 311788
rect 428004 311840 428056 311846
rect 428004 311782 428056 311788
rect 428016 309126 428044 311782
rect 428004 309120 428056 309126
rect 428004 309062 428056 309068
rect 428004 299532 428056 299538
rect 428004 299474 428056 299480
rect 428016 282946 428044 299474
rect 427820 282940 427872 282946
rect 427820 282882 427872 282888
rect 428004 282940 428056 282946
rect 428004 282882 428056 282888
rect 427832 282826 427860 282882
rect 427832 282798 427952 282826
rect 427924 273306 427952 282798
rect 427924 273278 428044 273306
rect 428016 263634 428044 273278
rect 427820 263628 427872 263634
rect 427820 263570 427872 263576
rect 428004 263628 428056 263634
rect 428004 263570 428056 263576
rect 427832 263514 427860 263570
rect 427832 263486 427952 263514
rect 427924 253994 427952 263486
rect 427924 253966 428044 253994
rect 428016 244322 428044 253966
rect 427820 244316 427872 244322
rect 427820 244258 427872 244264
rect 428004 244316 428056 244322
rect 428004 244258 428056 244264
rect 427832 244202 427860 244258
rect 427832 244174 427952 244202
rect 427924 234682 427952 244174
rect 427924 234654 428044 234682
rect 428016 225010 428044 234654
rect 427820 225004 427872 225010
rect 427820 224946 427872 224952
rect 428004 225004 428056 225010
rect 428004 224946 428056 224952
rect 427832 224890 427860 224946
rect 427832 224862 427952 224890
rect 427924 215370 427952 224862
rect 427924 215342 428044 215370
rect 428016 205698 428044 215342
rect 427820 205692 427872 205698
rect 427820 205634 427872 205640
rect 428004 205692 428056 205698
rect 428004 205634 428056 205640
rect 427832 205578 427860 205634
rect 427832 205550 427952 205578
rect 427924 196058 427952 205550
rect 427924 196030 428044 196058
rect 428016 183546 428044 196030
rect 427924 183518 428044 183546
rect 427924 176730 427952 183518
rect 427912 176724 427964 176730
rect 427912 176666 427964 176672
rect 427912 173936 427964 173942
rect 427912 173878 427964 173884
rect 427924 167090 427952 173878
rect 427832 167062 427952 167090
rect 427832 166954 427860 167062
rect 427832 166926 427952 166954
rect 427924 164218 427952 166926
rect 427912 164212 427964 164218
rect 427912 164154 427964 164160
rect 427912 157344 427964 157350
rect 427912 157286 427964 157292
rect 427924 154578 427952 157286
rect 427924 154550 428044 154578
rect 428016 147694 428044 154550
rect 427820 147688 427872 147694
rect 428004 147688 428056 147694
rect 427872 147636 428004 147642
rect 427820 147630 428056 147636
rect 427832 147614 428044 147630
rect 428016 138106 428044 147614
rect 428004 138100 428056 138106
rect 428004 138042 428056 138048
rect 427912 135312 427964 135318
rect 427912 135254 427964 135260
rect 427542 134192 427598 134201
rect 427726 134192 427782 134201
rect 427598 134150 427726 134178
rect 427542 134127 427598 134136
rect 427726 134127 427782 134136
rect 427924 128466 427952 135254
rect 427832 128438 427952 128466
rect 427832 128330 427860 128438
rect 427832 128302 427952 128330
rect 427924 125594 427952 128302
rect 427912 125588 427964 125594
rect 427912 125530 427964 125536
rect 427912 118652 427964 118658
rect 427912 118594 427964 118600
rect 427924 115954 427952 118594
rect 427924 115926 428044 115954
rect 428016 109070 428044 115926
rect 427820 109064 427872 109070
rect 428004 109064 428056 109070
rect 427872 109012 427952 109018
rect 427820 109006 427952 109012
rect 428004 109006 428056 109012
rect 427832 108990 427952 109006
rect 427924 106282 427952 108990
rect 427912 106276 427964 106282
rect 427912 106218 427964 106224
rect 427912 99340 427964 99346
rect 427912 99282 427964 99288
rect 427924 96642 427952 99282
rect 427924 96614 428044 96642
rect 428016 89758 428044 96614
rect 427820 89752 427872 89758
rect 428004 89752 428056 89758
rect 427872 89700 427952 89706
rect 427820 89694 427952 89700
rect 428004 89694 428056 89700
rect 427832 89678 427952 89694
rect 427924 86970 427952 89678
rect 427912 86964 427964 86970
rect 427912 86906 427964 86912
rect 428004 77308 428056 77314
rect 428004 77250 428056 77256
rect 428016 70258 428044 77250
rect 427924 70230 428044 70258
rect 427924 60738 427952 70230
rect 427924 60710 428044 60738
rect 428016 51082 428044 60710
rect 427832 51054 428044 51082
rect 427832 50946 427860 51054
rect 427832 50918 427952 50946
rect 427924 31822 427952 50918
rect 427912 31816 427964 31822
rect 427912 31758 427964 31764
rect 427820 31748 427872 31754
rect 427820 31690 427872 31696
rect 427832 26330 427860 31690
rect 427832 26302 427952 26330
rect 427924 24857 427952 26302
rect 427910 24848 427966 24857
rect 427910 24783 427966 24792
rect 428094 24848 428150 24857
rect 428094 24783 428150 24792
rect 428108 12374 428136 24783
rect 427912 12368 427964 12374
rect 427912 12310 427964 12316
rect 428096 12368 428148 12374
rect 428096 12310 428148 12316
rect 427924 5234 427952 12310
rect 427912 5228 427964 5234
rect 427912 5170 427964 5176
rect 427544 4004 427596 4010
rect 427544 3946 427596 3952
rect 427084 3052 427136 3058
rect 427084 2994 427136 3000
rect 426624 2984 426676 2990
rect 426624 2926 426676 2932
rect 427556 480 427584 3946
rect 428476 3534 428504 331214
rect 428464 3528 428516 3534
rect 428464 3470 428516 3476
rect 429120 626 429148 337486
rect 429580 337414 429608 340068
rect 429764 340054 430238 340082
rect 430684 340054 430790 340082
rect 431144 340054 431434 340082
rect 429568 337408 429620 337414
rect 429568 337350 429620 337356
rect 429764 331242 429792 340054
rect 430488 337408 430540 337414
rect 430488 337350 430540 337356
rect 429304 331214 429792 331242
rect 429304 4146 429332 331214
rect 430500 4146 430528 337350
rect 430580 335640 430632 335646
rect 430580 335582 430632 335588
rect 429292 4140 429344 4146
rect 429292 4082 429344 4088
rect 429936 4140 429988 4146
rect 429936 4082 429988 4088
rect 430488 4140 430540 4146
rect 430488 4082 430540 4088
rect 428752 598 429148 626
rect 428752 480 428780 598
rect 429948 480 429976 4082
rect 430592 3194 430620 335582
rect 430684 5302 430712 340054
rect 431144 335646 431172 340054
rect 432064 337618 432092 340068
rect 432156 340054 432630 340082
rect 432052 337612 432104 337618
rect 432052 337554 432104 337560
rect 431868 337068 431920 337074
rect 431868 337010 431920 337016
rect 431224 336864 431276 336870
rect 431224 336806 431276 336812
rect 431132 335640 431184 335646
rect 431132 335582 431184 335588
rect 430672 5296 430724 5302
rect 430672 5238 430724 5244
rect 431132 4140 431184 4146
rect 431132 4082 431184 4088
rect 430580 3188 430632 3194
rect 430580 3130 430632 3136
rect 431144 480 431172 4082
rect 431236 3330 431264 336806
rect 431880 4146 431908 337010
rect 432156 5370 432184 340054
rect 433260 337210 433288 340068
rect 433352 340054 433918 340082
rect 434180 340054 434470 340082
rect 434824 340054 435114 340082
rect 433248 337204 433300 337210
rect 433248 337146 433300 337152
rect 432604 336796 432656 336802
rect 432604 336738 432656 336744
rect 432144 5364 432196 5370
rect 432144 5306 432196 5312
rect 431868 4140 431920 4146
rect 431868 4082 431920 4088
rect 432616 3670 432644 336738
rect 433248 164212 433300 164218
rect 433248 164154 433300 164160
rect 433260 154601 433288 164154
rect 433246 154592 433302 154601
rect 433246 154527 433302 154536
rect 432604 3664 432656 3670
rect 432604 3606 432656 3612
rect 433352 3602 433380 340054
rect 434180 333334 434208 340054
rect 434628 337612 434680 337618
rect 434628 337554 434680 337560
rect 433708 333328 433760 333334
rect 433708 333270 433760 333276
rect 434168 333328 434220 333334
rect 434168 333270 434220 333276
rect 433720 328438 433748 333270
rect 433708 328432 433760 328438
rect 433708 328374 433760 328380
rect 433800 318844 433852 318850
rect 433800 318786 433852 318792
rect 433812 311914 433840 318786
rect 433432 311908 433484 311914
rect 433432 311850 433484 311856
rect 433800 311908 433852 311914
rect 433800 311850 433852 311856
rect 433444 309126 433472 311850
rect 433432 309120 433484 309126
rect 433432 309062 433484 309068
rect 433708 299532 433760 299538
rect 433708 299474 433760 299480
rect 433720 285002 433748 299474
rect 433628 284974 433748 285002
rect 433628 280158 433656 284974
rect 433616 280152 433668 280158
rect 433616 280094 433668 280100
rect 433708 270564 433760 270570
rect 433708 270506 433760 270512
rect 433720 263514 433748 270506
rect 433628 263486 433748 263514
rect 433628 260846 433656 263486
rect 433616 260840 433668 260846
rect 433616 260782 433668 260788
rect 433708 251252 433760 251258
rect 433708 251194 433760 251200
rect 433720 244202 433748 251194
rect 433628 244174 433748 244202
rect 433628 241505 433656 244174
rect 433430 241496 433486 241505
rect 433430 241431 433486 241440
rect 433614 241496 433670 241505
rect 433614 241431 433670 241440
rect 433444 231878 433472 241431
rect 433432 231872 433484 231878
rect 433432 231814 433484 231820
rect 433708 231872 433760 231878
rect 433708 231814 433760 231820
rect 433720 224890 433748 231814
rect 433628 224862 433748 224890
rect 433628 222193 433656 224862
rect 433430 222184 433486 222193
rect 433430 222119 433486 222128
rect 433614 222184 433670 222193
rect 433614 222119 433670 222128
rect 433444 212566 433472 222119
rect 433432 212560 433484 212566
rect 433432 212502 433484 212508
rect 433708 212560 433760 212566
rect 433708 212502 433760 212508
rect 433720 205578 433748 212502
rect 433628 205550 433748 205578
rect 433628 202881 433656 205550
rect 433430 202872 433486 202881
rect 433430 202807 433486 202816
rect 433614 202872 433670 202881
rect 433614 202807 433670 202816
rect 433444 193254 433472 202807
rect 433432 193248 433484 193254
rect 433432 193190 433484 193196
rect 433708 193248 433760 193254
rect 433708 193190 433760 193196
rect 433720 186266 433748 193190
rect 433628 186238 433748 186266
rect 433628 176662 433656 186238
rect 433616 176656 433668 176662
rect 433616 176598 433668 176604
rect 433616 173936 433668 173942
rect 433616 173878 433668 173884
rect 433628 166954 433656 173878
rect 434534 170096 434590 170105
rect 434534 170031 434590 170040
rect 434548 169862 434576 170031
rect 434536 169856 434588 169862
rect 434536 169798 434588 169804
rect 433444 166926 433656 166954
rect 433444 164218 433472 166926
rect 433432 164212 433484 164218
rect 433432 164154 433484 164160
rect 433706 154592 433762 154601
rect 433706 154527 433762 154536
rect 433720 147642 433748 154527
rect 433628 147614 433748 147642
rect 433628 144906 433656 147614
rect 433616 144900 433668 144906
rect 433616 144842 433668 144848
rect 433800 144900 433852 144906
rect 433800 144842 433852 144848
rect 433812 135289 433840 144842
rect 433614 135280 433670 135289
rect 433614 135215 433670 135224
rect 433798 135280 433854 135289
rect 433798 135215 433854 135224
rect 433628 125594 433656 135215
rect 433616 125588 433668 125594
rect 433616 125530 433668 125536
rect 433616 118652 433668 118658
rect 433616 118594 433668 118600
rect 433628 115954 433656 118594
rect 433628 115926 433748 115954
rect 433720 109018 433748 115926
rect 433628 108990 433748 109018
rect 433628 101402 433656 108990
rect 433444 101374 433656 101402
rect 433444 96665 433472 101374
rect 433430 96656 433486 96665
rect 433430 96591 433486 96600
rect 433706 96656 433762 96665
rect 433706 96591 433762 96600
rect 433720 89706 433748 96591
rect 433536 89678 433748 89706
rect 433536 86970 433564 89678
rect 433524 86964 433576 86970
rect 433524 86906 433576 86912
rect 433432 77308 433484 77314
rect 433432 77250 433484 77256
rect 433444 67658 433472 77250
rect 433432 67652 433484 67658
rect 433432 67594 433484 67600
rect 433524 67652 433576 67658
rect 433524 67594 433576 67600
rect 433536 60722 433564 67594
rect 433524 60716 433576 60722
rect 433524 60658 433576 60664
rect 433708 60716 433760 60722
rect 433708 60658 433760 60664
rect 433720 57934 433748 60658
rect 433708 57928 433760 57934
rect 433708 57870 433760 57876
rect 433616 48340 433668 48346
rect 433616 48282 433668 48288
rect 433628 41342 433656 48282
rect 433616 41336 433668 41342
rect 433616 41278 433668 41284
rect 433524 37392 433576 37398
rect 433576 37340 433656 37346
rect 433524 37334 433656 37340
rect 433536 37318 433656 37334
rect 433628 37262 433656 37318
rect 433616 37256 433668 37262
rect 433616 37198 433668 37204
rect 433708 27668 433760 27674
rect 433708 27610 433760 27616
rect 433720 22794 433748 27610
rect 433628 22766 433748 22794
rect 433628 5438 433656 22766
rect 433616 5432 433668 5438
rect 433616 5374 433668 5380
rect 434640 4146 434668 337554
rect 433524 4140 433576 4146
rect 433524 4082 433576 4088
rect 434628 4140 434680 4146
rect 434628 4082 434680 4088
rect 433340 3596 433392 3602
rect 433340 3538 433392 3544
rect 432328 3528 432380 3534
rect 432328 3470 432380 3476
rect 431224 3324 431276 3330
rect 431224 3266 431276 3272
rect 432340 480 432368 3470
rect 433536 480 433564 4082
rect 434824 3806 434852 340054
rect 435364 336864 435416 336870
rect 435364 336806 435416 336812
rect 434812 3800 434864 3806
rect 434812 3742 434864 3748
rect 434536 3732 434588 3738
rect 434536 3674 434588 3680
rect 434548 1850 434576 3674
rect 435376 3398 435404 336806
rect 435744 336802 435772 340068
rect 436204 340054 436310 340082
rect 436008 337068 436060 337074
rect 436008 337010 436060 337016
rect 435732 336796 435784 336802
rect 435732 336738 435784 336744
rect 435364 3392 435416 3398
rect 435364 3334 435416 3340
rect 434548 1822 434668 1850
rect 434640 480 434668 1822
rect 436020 610 436048 337010
rect 436204 5506 436232 340054
rect 436940 336802 436968 340068
rect 437598 340054 437704 340082
rect 436928 336796 436980 336802
rect 436928 336738 436980 336744
rect 436192 5500 436244 5506
rect 436192 5442 436244 5448
rect 437020 4140 437072 4146
rect 437020 4082 437072 4088
rect 435824 604 435876 610
rect 435824 546 435876 552
rect 436008 604 436060 610
rect 436008 546 436060 552
rect 435836 480 435864 546
rect 437032 480 437060 4082
rect 437676 3874 437704 340054
rect 437768 340054 438150 340082
rect 437768 4758 437796 340054
rect 438780 337006 438808 340068
rect 438964 340054 439438 340082
rect 438768 337000 438820 337006
rect 438768 336942 438820 336948
rect 438124 336796 438176 336802
rect 438124 336738 438176 336744
rect 437756 4752 437808 4758
rect 437756 4694 437808 4700
rect 437664 3868 437716 3874
rect 437664 3810 437716 3816
rect 438136 3262 438164 336738
rect 438964 4078 438992 340054
rect 439976 337822 440004 340068
rect 439964 337816 440016 337822
rect 439964 337758 440016 337764
rect 440620 336938 440648 340068
rect 441264 337890 441292 340068
rect 441252 337884 441304 337890
rect 441252 337826 441304 337832
rect 441816 337754 441844 340068
rect 441804 337748 441856 337754
rect 441804 337690 441856 337696
rect 442356 337748 442408 337754
rect 442356 337690 442408 337696
rect 442264 337340 442316 337346
rect 442264 337282 442316 337288
rect 440608 336932 440660 336938
rect 440608 336874 440660 336880
rect 438952 4072 439004 4078
rect 438952 4014 439004 4020
rect 440608 4072 440660 4078
rect 440608 4014 440660 4020
rect 438216 3800 438268 3806
rect 438216 3742 438268 3748
rect 438124 3256 438176 3262
rect 438124 3198 438176 3204
rect 438228 480 438256 3742
rect 439412 3596 439464 3602
rect 439412 3538 439464 3544
rect 439424 480 439452 3538
rect 440620 480 440648 4014
rect 442276 3942 442304 337282
rect 442368 4146 442396 337690
rect 442460 336870 442488 340068
rect 443012 337958 443040 340068
rect 443656 338026 443684 340068
rect 443644 338020 443696 338026
rect 443644 337962 443696 337968
rect 443000 337952 443052 337958
rect 443000 337894 443052 337900
rect 442448 336864 442500 336870
rect 442448 336806 442500 336812
rect 444300 336802 444328 340068
rect 444576 340054 444866 340082
rect 444288 336796 444340 336802
rect 444288 336738 444340 336744
rect 442356 4140 442408 4146
rect 442356 4082 442408 4088
rect 442264 3936 442316 3942
rect 442264 3878 442316 3884
rect 443000 3664 443052 3670
rect 443000 3606 443052 3612
rect 441804 3324 441856 3330
rect 441804 3266 441856 3272
rect 441816 480 441844 3266
rect 443012 480 443040 3606
rect 444196 3460 444248 3466
rect 444196 3402 444248 3408
rect 444208 480 444236 3402
rect 444576 3398 444604 340054
rect 445496 338094 445524 340068
rect 445484 338088 445536 338094
rect 445484 338030 445536 338036
rect 445024 337816 445076 337822
rect 445024 337758 445076 337764
rect 445036 4078 445064 337758
rect 446140 337686 446168 340068
rect 446128 337680 446180 337686
rect 446128 337622 446180 337628
rect 446692 337550 446720 340068
rect 446680 337544 446732 337550
rect 446680 337486 446732 337492
rect 446404 337476 446456 337482
rect 446404 337418 446456 337424
rect 445024 4072 445076 4078
rect 445024 4014 445076 4020
rect 446416 3466 446444 337418
rect 447336 337414 447364 340068
rect 447324 337408 447376 337414
rect 447324 337350 447376 337356
rect 447980 337278 448008 340068
rect 448428 337408 448480 337414
rect 448428 337350 448480 337356
rect 447968 337272 448020 337278
rect 447968 337214 448020 337220
rect 446496 336796 446548 336802
rect 446496 336738 446548 336744
rect 447784 336796 447836 336802
rect 447784 336738 447836 336744
rect 446508 3738 446536 336738
rect 447796 3806 447824 336738
rect 447784 3800 447836 3806
rect 447784 3742 447836 3748
rect 446496 3732 446548 3738
rect 446496 3674 446548 3680
rect 448440 3602 448468 337350
rect 448532 4010 448560 340068
rect 449176 337210 449204 340068
rect 449256 337680 449308 337686
rect 449256 337622 449308 337628
rect 449164 337204 449216 337210
rect 449164 337146 449216 337152
rect 449268 334506 449296 337622
rect 449820 337346 449848 340068
rect 450372 338026 450400 340068
rect 450360 338020 450412 338026
rect 450360 337962 450412 337968
rect 451016 337890 451044 340068
rect 451004 337884 451056 337890
rect 451004 337826 451056 337832
rect 451188 337544 451240 337550
rect 451188 337486 451240 337492
rect 449808 337340 449860 337346
rect 449808 337282 449860 337288
rect 449176 334478 449296 334506
rect 448520 4004 448572 4010
rect 448520 3946 448572 3952
rect 448980 3868 449032 3874
rect 448980 3810 449032 3816
rect 447784 3596 447836 3602
rect 447784 3538 447836 3544
rect 448428 3596 448480 3602
rect 448428 3538 448480 3544
rect 446404 3460 446456 3466
rect 446404 3402 446456 3408
rect 446588 3460 446640 3466
rect 446588 3402 446640 3408
rect 444564 3392 444616 3398
rect 444564 3334 444616 3340
rect 445392 3052 445444 3058
rect 445392 2994 445444 3000
rect 445404 480 445432 2994
rect 446600 480 446628 3402
rect 447796 480 447824 3538
rect 448992 480 449020 3810
rect 449176 3330 449204 334478
rect 451200 3738 451228 337486
rect 451660 337142 451688 340068
rect 451752 338094 451780 340190
rect 451740 338088 451792 338094
rect 451740 338030 451792 338036
rect 451924 338020 451976 338026
rect 451924 337962 451976 337968
rect 451648 337136 451700 337142
rect 451648 337078 451700 337084
rect 451556 330540 451608 330546
rect 451556 330482 451608 330488
rect 451568 325689 451596 330482
rect 451554 325680 451610 325689
rect 451554 325615 451610 325624
rect 451738 325680 451794 325689
rect 451738 325615 451794 325624
rect 451752 316130 451780 325615
rect 451556 316124 451608 316130
rect 451556 316066 451608 316072
rect 451740 316124 451792 316130
rect 451740 316066 451792 316072
rect 451568 315994 451596 316066
rect 451556 315988 451608 315994
rect 451556 315930 451608 315936
rect 451556 302116 451608 302122
rect 451556 302058 451608 302064
rect 451568 292670 451596 302058
rect 451556 292664 451608 292670
rect 451556 292606 451608 292612
rect 451464 292528 451516 292534
rect 451464 292470 451516 292476
rect 451476 288425 451504 292470
rect 451278 288416 451334 288425
rect 451278 288351 451334 288360
rect 451462 288416 451518 288425
rect 451462 288351 451518 288360
rect 451292 278798 451320 288351
rect 451280 278792 451332 278798
rect 451280 278734 451332 278740
rect 451556 278792 451608 278798
rect 451556 278734 451608 278740
rect 451568 273766 451596 278734
rect 451556 273760 451608 273766
rect 451556 273702 451608 273708
rect 451556 263492 451608 263498
rect 451556 263434 451608 263440
rect 451568 259418 451596 263434
rect 451556 259412 451608 259418
rect 451556 259354 451608 259360
rect 451556 244180 451608 244186
rect 451556 244122 451608 244128
rect 451568 234734 451596 244122
rect 451556 234728 451608 234734
rect 451556 234670 451608 234676
rect 451464 234592 451516 234598
rect 451464 234534 451516 234540
rect 451476 231849 451504 234534
rect 451278 231840 451334 231849
rect 451278 231775 451334 231784
rect 451462 231840 451518 231849
rect 451462 231775 451518 231784
rect 451292 222222 451320 231775
rect 451280 222216 451332 222222
rect 451280 222158 451332 222164
rect 451556 222216 451608 222222
rect 451556 222158 451608 222164
rect 451568 215422 451596 222158
rect 451556 215416 451608 215422
rect 451556 215358 451608 215364
rect 451464 215280 451516 215286
rect 451464 215222 451516 215228
rect 451476 212537 451504 215222
rect 451278 212528 451334 212537
rect 451278 212463 451334 212472
rect 451462 212528 451518 212537
rect 451462 212463 451518 212472
rect 451292 202910 451320 212463
rect 451280 202904 451332 202910
rect 451280 202846 451332 202852
rect 451556 202904 451608 202910
rect 451556 202846 451608 202852
rect 451568 196110 451596 202846
rect 451556 196104 451608 196110
rect 451556 196046 451608 196052
rect 451464 195968 451516 195974
rect 451464 195910 451516 195916
rect 451476 186318 451504 195910
rect 451464 186312 451516 186318
rect 451464 186254 451516 186260
rect 451648 186312 451700 186318
rect 451648 186254 451700 186260
rect 451660 183530 451688 186254
rect 451648 183524 451700 183530
rect 451648 183466 451700 183472
rect 451740 173936 451792 173942
rect 451740 173878 451792 173884
rect 451752 166954 451780 173878
rect 451660 166926 451780 166954
rect 451660 157350 451688 166926
rect 451648 157344 451700 157350
rect 451648 157286 451700 157292
rect 451648 157208 451700 157214
rect 451648 157150 451700 157156
rect 451660 154562 451688 157150
rect 451648 154556 451700 154562
rect 451648 154498 451700 154504
rect 451648 147620 451700 147626
rect 451648 147562 451700 147568
rect 451660 144922 451688 147562
rect 451660 144894 451780 144922
rect 451752 135318 451780 144894
rect 451648 135312 451700 135318
rect 451568 135260 451648 135266
rect 451568 135254 451700 135260
rect 451740 135312 451792 135318
rect 451740 135254 451792 135260
rect 451568 135238 451688 135254
rect 451568 128466 451596 135238
rect 451568 128438 451688 128466
rect 451660 128194 451688 128438
rect 451476 128166 451688 128194
rect 451476 124166 451504 128166
rect 451464 124160 451516 124166
rect 451464 124102 451516 124108
rect 451556 114572 451608 114578
rect 451556 114514 451608 114520
rect 451568 104854 451596 114514
rect 451556 104848 451608 104854
rect 451556 104790 451608 104796
rect 451556 95260 451608 95266
rect 451556 95202 451608 95208
rect 451568 85542 451596 95202
rect 451556 85536 451608 85542
rect 451556 85478 451608 85484
rect 451464 67652 451516 67658
rect 451464 67594 451516 67600
rect 451476 66230 451504 67594
rect 451464 66224 451516 66230
rect 451464 66166 451516 66172
rect 451648 60716 451700 60722
rect 451648 60658 451700 60664
rect 451660 56574 451688 60658
rect 451648 56568 451700 56574
rect 451648 56510 451700 56516
rect 451832 46980 451884 46986
rect 451832 46922 451884 46928
rect 451844 46866 451872 46922
rect 451660 46838 451872 46866
rect 451660 31754 451688 46838
rect 451648 31748 451700 31754
rect 451648 31690 451700 31696
rect 451832 31748 451884 31754
rect 451832 31690 451884 31696
rect 451844 28966 451872 31690
rect 451832 28960 451884 28966
rect 451832 28902 451884 28908
rect 451740 19372 451792 19378
rect 451740 19314 451792 19320
rect 451752 12458 451780 19314
rect 451568 12430 451780 12458
rect 451280 4140 451332 4146
rect 451280 4082 451332 4088
rect 450176 3732 450228 3738
rect 450176 3674 450228 3680
rect 451188 3732 451240 3738
rect 451188 3674 451240 3680
rect 449164 3324 449216 3330
rect 449164 3266 449216 3272
rect 450188 480 450216 3674
rect 451292 480 451320 4082
rect 451568 3534 451596 12430
rect 451556 3528 451608 3534
rect 451556 3470 451608 3476
rect 451936 3058 451964 337962
rect 452856 337618 452884 340068
rect 453304 337884 453356 337890
rect 453304 337826 453356 337832
rect 452844 337612 452896 337618
rect 452844 337554 452896 337560
rect 453316 4146 453344 337826
rect 453396 337204 453448 337210
rect 453396 337146 453448 337152
rect 453304 4140 453356 4146
rect 453304 4082 453356 4088
rect 453408 3874 453436 337146
rect 453500 336938 453528 340068
rect 453948 337612 454000 337618
rect 453948 337554 454000 337560
rect 453488 336932 453540 336938
rect 453488 336874 453540 336880
rect 453396 3868 453448 3874
rect 453396 3810 453448 3816
rect 452476 3460 452528 3466
rect 452476 3402 452528 3408
rect 451924 3052 451976 3058
rect 451924 2994 451976 3000
rect 452488 480 452516 3402
rect 453960 610 453988 337554
rect 454052 337074 454080 340068
rect 454696 337754 454724 340068
rect 454684 337748 454736 337754
rect 454684 337690 454736 337696
rect 454040 337068 454092 337074
rect 454040 337010 454092 337016
rect 455340 336802 455368 340068
rect 455616 340054 455906 340082
rect 455328 336796 455380 336802
rect 455328 336738 455380 336744
rect 454868 4140 454920 4146
rect 454868 4082 454920 4088
rect 453672 604 453724 610
rect 453672 546 453724 552
rect 453948 604 454000 610
rect 453948 546 454000 552
rect 453684 480 453712 546
rect 454880 480 454908 4082
rect 455616 3806 455644 340054
rect 456536 337822 456564 340068
rect 456524 337816 456576 337822
rect 456524 337758 456576 337764
rect 456064 337748 456116 337754
rect 456064 337690 456116 337696
rect 456076 4146 456104 337690
rect 457180 337686 457208 340068
rect 457168 337680 457220 337686
rect 457168 337622 457220 337628
rect 457272 331242 457300 340190
rect 458376 337482 458404 340068
rect 459020 338026 459048 340068
rect 459586 340054 459784 340082
rect 459008 338020 459060 338026
rect 459008 337962 459060 337968
rect 458364 337476 458416 337482
rect 458364 337418 458416 337424
rect 457444 336796 457496 336802
rect 457444 336738 457496 336744
rect 456904 331214 457300 331242
rect 456798 40352 456854 40361
rect 456798 40287 456854 40296
rect 456706 40216 456762 40225
rect 456812 40202 456840 40287
rect 456762 40174 456840 40202
rect 456706 40151 456762 40160
rect 456798 16960 456854 16969
rect 456798 16895 456854 16904
rect 456706 16824 456762 16833
rect 456812 16810 456840 16895
rect 456762 16782 456840 16810
rect 456706 16759 456762 16768
rect 456064 4140 456116 4146
rect 456064 4082 456116 4088
rect 455604 3800 455656 3806
rect 455604 3742 455656 3748
rect 456904 3670 456932 331214
rect 457260 3732 457312 3738
rect 457260 3674 457312 3680
rect 456892 3664 456944 3670
rect 456892 3606 456944 3612
rect 456064 2780 456116 2786
rect 456064 2722 456116 2728
rect 456076 480 456104 2722
rect 457272 480 457300 3674
rect 457456 3466 457484 336738
rect 458822 134056 458878 134065
rect 458822 133991 458878 134000
rect 458836 133793 458864 133991
rect 458822 133784 458878 133793
rect 458822 133719 458878 133728
rect 458456 4004 458508 4010
rect 458456 3946 458508 3952
rect 457444 3460 457496 3466
rect 457444 3402 457496 3408
rect 458468 480 458496 3946
rect 459756 3534 459784 340054
rect 460216 337414 460244 340068
rect 460204 337408 460256 337414
rect 460204 337350 460256 337356
rect 460768 337210 460796 340068
rect 461412 337550 461440 340068
rect 462056 337890 462084 340068
rect 462044 337884 462096 337890
rect 462044 337826 462096 337832
rect 461400 337544 461452 337550
rect 461400 337486 461452 337492
rect 460848 337408 460900 337414
rect 460848 337350 460900 337356
rect 460756 337204 460808 337210
rect 460756 337146 460808 337152
rect 460204 336932 460256 336938
rect 460204 336874 460256 336880
rect 459744 3528 459796 3534
rect 459744 3470 459796 3476
rect 459652 3392 459704 3398
rect 459652 3334 459704 3340
rect 459664 480 459692 3334
rect 460216 2854 460244 336874
rect 460204 2848 460256 2854
rect 460204 2790 460256 2796
rect 460860 480 460888 337350
rect 462608 336802 462636 340068
rect 463252 337618 463280 340068
rect 463608 337884 463660 337890
rect 463608 337826 463660 337832
rect 463240 337612 463292 337618
rect 463240 337554 463292 337560
rect 462596 336796 462648 336802
rect 462596 336738 462648 336744
rect 462044 3460 462096 3466
rect 462044 3402 462096 3408
rect 462056 480 462084 3402
rect 463620 2854 463648 337826
rect 463896 337754 463924 340068
rect 463884 337748 463936 337754
rect 463884 337690 463936 337696
rect 464448 336938 464476 340068
rect 465106 340054 465396 340082
rect 464988 337816 465040 337822
rect 464988 337758 465040 337764
rect 464436 336932 464488 336938
rect 464436 336874 464488 336880
rect 464344 336864 464396 336870
rect 464344 336806 464396 336812
rect 464356 3398 464384 336806
rect 464436 336796 464488 336802
rect 464436 336738 464488 336744
rect 464448 4010 464476 336738
rect 464436 4004 464488 4010
rect 464436 3946 464488 3952
rect 464344 3392 464396 3398
rect 464344 3334 464396 3340
rect 465000 3330 465028 337758
rect 465368 3738 465396 340054
rect 465736 336802 465764 340068
rect 466288 336870 466316 340068
rect 466368 337680 466420 337686
rect 466368 337622 466420 337628
rect 466276 336864 466328 336870
rect 466276 336806 466328 336812
rect 465724 336796 465776 336802
rect 465724 336738 465776 336744
rect 465356 3732 465408 3738
rect 465356 3674 465408 3680
rect 464436 3324 464488 3330
rect 464436 3266 464488 3272
rect 464988 3324 465040 3330
rect 464988 3266 465040 3272
rect 463240 2848 463292 2854
rect 463240 2790 463292 2796
rect 463608 2848 463660 2854
rect 463608 2790 463660 2796
rect 463252 480 463280 2790
rect 464448 480 464476 3266
rect 466380 2922 466408 337622
rect 466932 337414 466960 340068
rect 467116 340054 467590 340082
rect 466920 337408 466972 337414
rect 466920 337350 466972 337356
rect 467116 333334 467144 340054
rect 468128 337890 468156 340068
rect 468116 337884 468168 337890
rect 468116 337826 468168 337832
rect 468772 337822 468800 340068
rect 468760 337816 468812 337822
rect 468760 337758 468812 337764
rect 469416 337686 469444 340068
rect 469404 337680 469456 337686
rect 469404 337622 469456 337628
rect 469968 336870 469996 340068
rect 470626 340054 470824 340082
rect 467748 336864 467800 336870
rect 467748 336806 467800 336812
rect 469956 336864 470008 336870
rect 469956 336806 470008 336812
rect 466552 333328 466604 333334
rect 466552 333270 466604 333276
rect 467104 333328 467156 333334
rect 467104 333270 467156 333276
rect 466564 321638 466592 333270
rect 466552 321632 466604 321638
rect 466552 321574 466604 321580
rect 466552 318844 466604 318850
rect 466552 318786 466604 318792
rect 466564 311930 466592 318786
rect 466472 311902 466592 311930
rect 466472 311846 466500 311902
rect 466460 311840 466512 311846
rect 466460 311782 466512 311788
rect 466644 311840 466696 311846
rect 466644 311782 466696 311788
rect 466656 309126 466684 311782
rect 466644 309120 466696 309126
rect 466644 309062 466696 309068
rect 466552 299532 466604 299538
rect 466552 299474 466604 299480
rect 466564 292618 466592 299474
rect 466472 292590 466592 292618
rect 466472 292534 466500 292590
rect 466460 292528 466512 292534
rect 466460 292470 466512 292476
rect 466644 292528 466696 292534
rect 466644 292470 466696 292476
rect 466656 280242 466684 292470
rect 466564 280214 466684 280242
rect 466564 280158 466592 280214
rect 466552 280152 466604 280158
rect 466552 280094 466604 280100
rect 466644 270564 466696 270570
rect 466644 270506 466696 270512
rect 466656 263514 466684 270506
rect 466564 263486 466684 263514
rect 466564 260846 466592 263486
rect 466552 260840 466604 260846
rect 466552 260782 466604 260788
rect 466644 251252 466696 251258
rect 466644 251194 466696 251200
rect 466656 244202 466684 251194
rect 466564 244174 466684 244202
rect 466564 241466 466592 244174
rect 466552 241460 466604 241466
rect 466552 241402 466604 241408
rect 466644 241460 466696 241466
rect 466644 241402 466696 241408
rect 466656 224890 466684 241402
rect 466564 224862 466684 224890
rect 466564 222154 466592 224862
rect 466552 222148 466604 222154
rect 466552 222090 466604 222096
rect 466644 222148 466696 222154
rect 466644 222090 466696 222096
rect 466656 205578 466684 222090
rect 466564 205550 466684 205578
rect 466564 202842 466592 205550
rect 466552 202836 466604 202842
rect 466552 202778 466604 202784
rect 466644 202836 466696 202842
rect 466644 202778 466696 202784
rect 466656 186266 466684 202778
rect 466564 186238 466684 186266
rect 466564 183530 466592 186238
rect 466552 183524 466604 183530
rect 466552 183466 466604 183472
rect 466644 183524 466696 183530
rect 466644 183466 466696 183472
rect 466656 166954 466684 183466
rect 466564 166926 466684 166954
rect 466564 157298 466592 166926
rect 466564 157270 466684 157298
rect 466656 154630 466684 157270
rect 466552 154624 466604 154630
rect 466552 154566 466604 154572
rect 466644 154624 466696 154630
rect 466644 154566 466696 154572
rect 466564 154494 466592 154566
rect 466552 154488 466604 154494
rect 466552 154430 466604 154436
rect 466552 147620 466604 147626
rect 466552 147562 466604 147568
rect 466564 144922 466592 147562
rect 466564 144894 466684 144922
rect 466656 138038 466684 144894
rect 466460 138032 466512 138038
rect 466460 137974 466512 137980
rect 466644 138032 466696 138038
rect 466644 137974 466696 137980
rect 466472 128382 466500 137974
rect 466460 128376 466512 128382
rect 466460 128318 466512 128324
rect 466552 128308 466604 128314
rect 466552 128250 466604 128256
rect 466564 125610 466592 128250
rect 466564 125594 466684 125610
rect 466564 125588 466696 125594
rect 466564 125582 466644 125588
rect 466644 125530 466696 125536
rect 466736 125588 466788 125594
rect 466736 125530 466788 125536
rect 466748 124166 466776 125530
rect 466736 124160 466788 124166
rect 466736 124102 466788 124108
rect 466644 114572 466696 114578
rect 466644 114514 466696 114520
rect 466656 109070 466684 114514
rect 466644 109064 466696 109070
rect 466644 109006 466696 109012
rect 466552 108996 466604 109002
rect 466552 108938 466604 108944
rect 466564 99414 466592 108938
rect 466552 99408 466604 99414
rect 466552 99350 466604 99356
rect 466460 99340 466512 99346
rect 466460 99282 466512 99288
rect 466472 96665 466500 99282
rect 466458 96656 466514 96665
rect 466458 96591 466514 96600
rect 466642 96656 466698 96665
rect 466642 96591 466698 96600
rect 466656 89706 466684 96591
rect 466564 89678 466684 89706
rect 466564 85542 466592 89678
rect 466552 85536 466604 85542
rect 466552 85478 466604 85484
rect 466644 75948 466696 75954
rect 466644 75890 466696 75896
rect 466656 67674 466684 75890
rect 466472 67646 466684 67674
rect 466472 66230 466500 67646
rect 466460 66224 466512 66230
rect 466460 66166 466512 66172
rect 466828 56636 466880 56642
rect 466828 56578 466880 56584
rect 466840 48346 466868 56578
rect 466644 48340 466696 48346
rect 466644 48282 466696 48288
rect 466828 48340 466880 48346
rect 466828 48282 466880 48288
rect 466656 29034 466684 48282
rect 466552 29028 466604 29034
rect 466552 28970 466604 28976
rect 466644 29028 466696 29034
rect 466644 28970 466696 28976
rect 466564 22114 466592 28970
rect 466564 22086 466684 22114
rect 466656 12458 466684 22086
rect 466472 12430 466684 12458
rect 466472 3466 466500 12430
rect 467760 3738 467788 336806
rect 469864 336796 469916 336802
rect 469864 336738 469916 336744
rect 469876 4146 469904 336738
rect 470692 335640 470744 335646
rect 470692 335582 470744 335588
rect 469128 4140 469180 4146
rect 469128 4082 469180 4088
rect 469864 4140 469916 4146
rect 469864 4082 469916 4088
rect 466828 3732 466880 3738
rect 466828 3674 466880 3680
rect 467748 3732 467800 3738
rect 467748 3674 467800 3680
rect 466460 3460 466512 3466
rect 466460 3402 466512 3408
rect 465632 2916 465684 2922
rect 465632 2858 465684 2864
rect 466368 2916 466420 2922
rect 466368 2858 466420 2864
rect 465644 480 465672 2858
rect 466840 480 466868 3674
rect 467932 3596 467984 3602
rect 467932 3538 467984 3544
rect 467944 480 467972 3538
rect 469140 480 469168 4082
rect 470704 3126 470732 335582
rect 470796 3602 470824 340054
rect 471256 336802 471284 340068
rect 471440 340054 471822 340082
rect 471992 340054 472466 340082
rect 472544 340054 473110 340082
rect 473372 340054 473662 340082
rect 474306 340054 474688 340082
rect 471244 336796 471296 336802
rect 471244 336738 471296 336744
rect 471440 335646 471468 340054
rect 471992 336818 472020 340054
rect 471900 336790 472020 336818
rect 471428 335640 471480 335646
rect 471428 335582 471480 335588
rect 470784 3596 470836 3602
rect 470784 3538 470836 3544
rect 470324 3120 470376 3126
rect 470324 3062 470376 3068
rect 470692 3120 470744 3126
rect 470692 3062 470744 3068
rect 470336 480 470364 3062
rect 471900 2854 471928 336790
rect 472544 333282 472572 340054
rect 472176 333254 472572 333282
rect 472176 328438 472204 333254
rect 472164 328432 472216 328438
rect 472164 328374 472216 328380
rect 472072 318844 472124 318850
rect 472072 318786 472124 318792
rect 472084 311930 472112 318786
rect 471992 311902 472112 311930
rect 471992 311846 472020 311902
rect 471980 311840 472032 311846
rect 471980 311782 472032 311788
rect 472164 311840 472216 311846
rect 472164 311782 472216 311788
rect 472176 309126 472204 311782
rect 472164 309120 472216 309126
rect 472164 309062 472216 309068
rect 472072 299532 472124 299538
rect 472072 299474 472124 299480
rect 472084 292618 472112 299474
rect 471992 292590 472112 292618
rect 471992 292534 472020 292590
rect 471980 292528 472032 292534
rect 471980 292470 472032 292476
rect 472164 292528 472216 292534
rect 472164 292470 472216 292476
rect 472176 280242 472204 292470
rect 472084 280214 472204 280242
rect 472084 280158 472112 280214
rect 472072 280152 472124 280158
rect 472072 280094 472124 280100
rect 472164 270564 472216 270570
rect 472164 270506 472216 270512
rect 472176 263514 472204 270506
rect 472084 263486 472204 263514
rect 472084 260846 472112 263486
rect 472072 260840 472124 260846
rect 472072 260782 472124 260788
rect 472164 251252 472216 251258
rect 472164 251194 472216 251200
rect 472176 244202 472204 251194
rect 472084 244174 472204 244202
rect 472084 241505 472112 244174
rect 472070 241496 472126 241505
rect 472070 241431 472126 241440
rect 472346 241496 472402 241505
rect 472346 241431 472402 241440
rect 472360 231878 472388 241431
rect 472164 231872 472216 231878
rect 472164 231814 472216 231820
rect 472348 231872 472400 231878
rect 472348 231814 472400 231820
rect 472176 224890 472204 231814
rect 472084 224862 472204 224890
rect 472084 222193 472112 224862
rect 472070 222184 472126 222193
rect 472070 222119 472126 222128
rect 472346 222184 472402 222193
rect 472346 222119 472402 222128
rect 472360 212566 472388 222119
rect 472164 212560 472216 212566
rect 472164 212502 472216 212508
rect 472348 212560 472400 212566
rect 472348 212502 472400 212508
rect 472176 205578 472204 212502
rect 472084 205550 472204 205578
rect 472084 202881 472112 205550
rect 472070 202872 472126 202881
rect 472070 202807 472126 202816
rect 472346 202872 472402 202881
rect 472346 202807 472402 202816
rect 472360 193254 472388 202807
rect 472164 193248 472216 193254
rect 472164 193190 472216 193196
rect 472348 193248 472400 193254
rect 472348 193190 472400 193196
rect 472176 186266 472204 193190
rect 472084 186238 472204 186266
rect 472084 183569 472112 186238
rect 472070 183560 472126 183569
rect 472070 183495 472126 183504
rect 472346 183560 472402 183569
rect 472346 183495 472402 183504
rect 472360 173942 472388 183495
rect 472164 173936 472216 173942
rect 472164 173878 472216 173884
rect 472348 173936 472400 173942
rect 472348 173878 472400 173884
rect 472176 166954 472204 173878
rect 472084 166926 472204 166954
rect 472084 164218 472112 166926
rect 472072 164212 472124 164218
rect 472072 164154 472124 164160
rect 472348 164212 472400 164218
rect 472348 164154 472400 164160
rect 472360 154601 472388 164154
rect 472162 154592 472218 154601
rect 472162 154527 472218 154536
rect 472346 154592 472402 154601
rect 472346 154527 472402 154536
rect 472176 147642 472204 154527
rect 472084 147614 472204 147642
rect 472084 143546 472112 147614
rect 472072 143540 472124 143546
rect 472072 143482 472124 143488
rect 472072 128308 472124 128314
rect 472072 128250 472124 128256
rect 472084 118726 472112 128250
rect 472072 118720 472124 118726
rect 472072 118662 472124 118668
rect 471980 118652 472032 118658
rect 471980 118594 472032 118600
rect 471992 115977 472020 118594
rect 471978 115968 472034 115977
rect 471978 115903 472034 115912
rect 472162 115968 472218 115977
rect 472162 115903 472218 115912
rect 472176 109018 472204 115903
rect 472084 108990 472204 109018
rect 472084 99414 472112 108990
rect 472072 99408 472124 99414
rect 472072 99350 472124 99356
rect 471980 99340 472032 99346
rect 471980 99282 472032 99288
rect 471992 96665 472020 99282
rect 471978 96656 472034 96665
rect 471978 96591 472034 96600
rect 472162 96656 472218 96665
rect 472162 96591 472218 96600
rect 472176 89706 472204 96591
rect 472084 89678 472204 89706
rect 472084 80782 472112 89678
rect 472072 80776 472124 80782
rect 472072 80718 472124 80724
rect 472072 67652 472124 67658
rect 472072 67594 472124 67600
rect 472084 60738 472112 67594
rect 471992 60722 472112 60738
rect 471980 60716 472112 60722
rect 472032 60710 472112 60716
rect 472164 60716 472216 60722
rect 471980 60658 472032 60664
rect 472164 60658 472216 60664
rect 472176 57934 472204 60658
rect 472164 57928 472216 57934
rect 472164 57870 472216 57876
rect 472072 48340 472124 48346
rect 472072 48282 472124 48288
rect 472084 41426 472112 48282
rect 471992 41410 472112 41426
rect 471980 41404 472112 41410
rect 472032 41398 472112 41404
rect 472164 41404 472216 41410
rect 471980 41346 472032 41352
rect 472164 41346 472216 41352
rect 472176 38622 472204 41346
rect 472164 38616 472216 38622
rect 472164 38558 472216 38564
rect 472072 29028 472124 29034
rect 472072 28970 472124 28976
rect 472084 24154 472112 28970
rect 472084 24126 472204 24154
rect 472176 4146 472204 24126
rect 473372 4146 473400 340054
rect 474660 4146 474688 340054
rect 474936 336802 474964 340068
rect 475488 337686 475516 340068
rect 475476 337680 475528 337686
rect 475476 337622 475528 337628
rect 476132 336938 476160 340068
rect 476790 340054 477264 340082
rect 477236 337736 477264 340054
rect 477328 338026 477356 340068
rect 477316 338020 477368 338026
rect 477316 337962 477368 337968
rect 477972 337754 478000 340068
rect 477960 337748 478012 337754
rect 477236 337708 477448 337736
rect 476120 336932 476172 336938
rect 476120 336874 476172 336880
rect 474924 336796 474976 336802
rect 474924 336738 474976 336744
rect 476028 336796 476080 336802
rect 476028 336738 476080 336744
rect 475934 169960 475990 169969
rect 475934 169895 475936 169904
rect 475988 169895 475990 169904
rect 475936 169866 475988 169872
rect 475936 40248 475988 40254
rect 475934 40216 475936 40225
rect 475988 40216 475990 40225
rect 475934 40151 475990 40160
rect 475936 16856 475988 16862
rect 475934 16824 475936 16833
rect 475988 16824 475990 16833
rect 475934 16759 475990 16768
rect 472164 4140 472216 4146
rect 472164 4082 472216 4088
rect 472716 4140 472768 4146
rect 472716 4082 472768 4088
rect 473360 4140 473412 4146
rect 473360 4082 473412 4088
rect 473912 4140 473964 4146
rect 473912 4082 473964 4088
rect 474648 4140 474700 4146
rect 474648 4082 474700 4088
rect 475108 4140 475160 4146
rect 475108 4082 475160 4088
rect 471520 2848 471572 2854
rect 471520 2790 471572 2796
rect 471888 2848 471940 2854
rect 471888 2790 471940 2796
rect 471532 480 471560 2790
rect 472728 480 472756 4082
rect 473924 480 473952 4082
rect 475120 480 475148 4082
rect 476040 3482 476068 336738
rect 476040 3454 476344 3482
rect 476316 480 476344 3454
rect 477420 3058 477448 337708
rect 477960 337690 478012 337696
rect 477592 337680 477644 337686
rect 477592 337622 477644 337628
rect 477500 16856 477552 16862
rect 477498 16824 477500 16833
rect 477552 16824 477554 16833
rect 477498 16759 477554 16768
rect 477604 3482 477632 337622
rect 478524 337618 478552 340068
rect 479168 337754 479196 340068
rect 478788 337748 478840 337754
rect 478788 337690 478840 337696
rect 479156 337748 479208 337754
rect 479156 337690 479208 337696
rect 478512 337612 478564 337618
rect 478512 337554 478564 337560
rect 477776 336932 477828 336938
rect 477776 336874 477828 336880
rect 477512 3454 477632 3482
rect 477408 3052 477460 3058
rect 477408 2994 477460 3000
rect 477512 480 477540 3454
rect 477788 610 477816 336874
rect 478142 169960 478198 169969
rect 478142 169895 478144 169904
rect 478196 169895 478198 169904
rect 478144 169866 478196 169872
rect 478236 40248 478288 40254
rect 478234 40216 478236 40225
rect 478288 40216 478290 40225
rect 478234 40151 478290 40160
rect 478800 3670 478828 337690
rect 479812 337550 479840 340068
rect 480260 338020 480312 338026
rect 480260 337962 480312 337968
rect 480272 337634 480300 337962
rect 480364 337754 480392 340068
rect 480352 337748 480404 337754
rect 480352 337690 480404 337696
rect 480272 337606 480392 337634
rect 479800 337544 479852 337550
rect 479800 337486 479852 337492
rect 478788 3664 478840 3670
rect 478788 3606 478840 3612
rect 479892 3052 479944 3058
rect 479892 2994 479944 3000
rect 477776 604 477828 610
rect 477776 546 477828 552
rect 478696 604 478748 610
rect 478696 546 478748 552
rect 478708 480 478736 546
rect 479904 480 479932 2994
rect 480364 610 480392 337606
rect 481008 337482 481036 340068
rect 481548 337748 481600 337754
rect 481548 337690 481600 337696
rect 480996 337476 481048 337482
rect 480996 337418 481048 337424
rect 481560 3330 481588 337690
rect 481652 337550 481680 340068
rect 482218 340054 482784 340082
rect 482756 337668 482784 340054
rect 482848 337822 482876 340068
rect 482836 337816 482888 337822
rect 482836 337758 482888 337764
rect 483492 337686 483520 340068
rect 484058 340054 484348 340082
rect 483480 337680 483532 337686
rect 482756 337640 482968 337668
rect 481640 337544 481692 337550
rect 481640 337486 481692 337492
rect 482836 337544 482888 337550
rect 482836 337486 482888 337492
rect 482284 3664 482336 3670
rect 482284 3606 482336 3612
rect 481548 3324 481600 3330
rect 481548 3266 481600 3272
rect 480352 604 480404 610
rect 480352 546 480404 552
rect 481088 604 481140 610
rect 481088 546 481140 552
rect 481100 480 481128 546
rect 482296 480 482324 3606
rect 482848 3398 482876 337486
rect 482940 3874 482968 337640
rect 483480 337622 483532 337628
rect 484216 337680 484268 337686
rect 484216 337622 484268 337628
rect 483204 337612 483256 337618
rect 483204 337554 483256 337560
rect 482928 3868 482980 3874
rect 482928 3810 482980 3816
rect 482836 3392 482888 3398
rect 482836 3334 482888 3340
rect 483216 626 483244 337554
rect 484228 3670 484256 337622
rect 484216 3664 484268 3670
rect 484216 3606 484268 3612
rect 484320 3602 484348 340054
rect 484584 337612 484636 337618
rect 484584 337554 484636 337560
rect 484308 3596 484360 3602
rect 484308 3538 484360 3544
rect 483216 598 483520 626
rect 483492 480 483520 598
rect 484596 480 484624 337554
rect 484688 337414 484716 340068
rect 485332 337482 485360 340068
rect 485884 337686 485912 340068
rect 486542 340054 487108 340082
rect 485872 337680 485924 337686
rect 485872 337622 485924 337628
rect 485044 337476 485096 337482
rect 485044 337418 485096 337424
rect 485320 337476 485372 337482
rect 485320 337418 485372 337424
rect 484676 337408 484728 337414
rect 484676 337350 484728 337356
rect 485056 3262 485084 337418
rect 485688 337408 485740 337414
rect 485688 337350 485740 337356
rect 485700 3738 485728 337350
rect 485964 337340 486016 337346
rect 485964 337282 486016 337288
rect 485688 3732 485740 3738
rect 485688 3674 485740 3680
rect 485044 3256 485096 3262
rect 485044 3198 485096 3204
rect 485976 626 486004 337282
rect 487080 3534 487108 340054
rect 487172 337890 487200 340068
rect 487160 337884 487212 337890
rect 487160 337826 487212 337832
rect 487724 337074 487752 340068
rect 487712 337068 487764 337074
rect 487712 337010 487764 337016
rect 487068 3528 487120 3534
rect 487068 3470 487120 3476
rect 488368 3330 488396 340068
rect 489012 337754 489040 340068
rect 489578 340054 489868 340082
rect 489000 337748 489052 337754
rect 489000 337690 489052 337696
rect 489184 337680 489236 337686
rect 489184 337622 489236 337628
rect 488448 337068 488500 337074
rect 488448 337010 488500 337016
rect 488460 3466 488488 337010
rect 489196 3806 489224 337622
rect 489184 3800 489236 3806
rect 489184 3742 489236 3748
rect 488448 3460 488500 3466
rect 488448 3402 488500 3408
rect 489368 3392 489420 3398
rect 489368 3334 489420 3340
rect 486976 3324 487028 3330
rect 486976 3266 487028 3272
rect 488356 3324 488408 3330
rect 488356 3266 488408 3272
rect 485792 598 486004 626
rect 485792 480 485820 598
rect 486988 480 487016 3266
rect 488172 3256 488224 3262
rect 488172 3198 488224 3204
rect 488184 480 488212 3198
rect 489380 480 489408 3334
rect 489840 3262 489868 340054
rect 490208 337958 490236 340068
rect 490852 338094 490880 340068
rect 490840 338088 490892 338094
rect 490840 338030 490892 338036
rect 490196 337952 490248 337958
rect 490196 337894 490248 337900
rect 491404 337686 491432 340068
rect 492062 340054 492536 340082
rect 491392 337680 491444 337686
rect 491392 337622 491444 337628
rect 491484 337408 491536 337414
rect 491484 337350 491536 337356
rect 490564 3868 490616 3874
rect 490564 3810 490616 3816
rect 489828 3256 489880 3262
rect 489828 3198 489880 3204
rect 490576 480 490604 3810
rect 491496 626 491524 337350
rect 492508 4078 492536 340054
rect 492588 337680 492640 337686
rect 492588 337622 492640 337628
rect 492496 4072 492548 4078
rect 492496 4014 492548 4020
rect 492600 3398 492628 337622
rect 492692 337618 492720 340068
rect 493244 337686 493272 340068
rect 493232 337680 493284 337686
rect 493232 337622 493284 337628
rect 492680 337612 492732 337618
rect 492680 337554 492732 337560
rect 493324 337476 493376 337482
rect 493324 337418 493376 337424
rect 492956 3664 493008 3670
rect 492956 3606 493008 3612
rect 492588 3392 492640 3398
rect 492588 3334 492640 3340
rect 491496 598 491708 626
rect 491680 592 491708 598
rect 491680 564 491800 592
rect 491772 480 491800 564
rect 492968 480 492996 3606
rect 493336 3194 493364 337418
rect 493888 4010 493916 340068
rect 493968 337680 494020 337686
rect 493968 337622 494020 337628
rect 493980 4146 494008 337622
rect 494532 337550 494560 340068
rect 494520 337544 494572 337550
rect 494520 337486 494572 337492
rect 495084 337074 495112 340068
rect 495728 337618 495756 340068
rect 495716 337612 495768 337618
rect 495716 337554 495768 337560
rect 496280 337482 496308 340068
rect 496924 337686 496952 340068
rect 497568 337822 497596 340068
rect 497556 337816 497608 337822
rect 497556 337758 497608 337764
rect 496912 337680 496964 337686
rect 496912 337622 496964 337628
rect 496728 337612 496780 337618
rect 496728 337554 496780 337560
rect 496268 337476 496320 337482
rect 496268 337418 496320 337424
rect 495072 337068 495124 337074
rect 495072 337010 495124 337016
rect 496084 337068 496136 337074
rect 496084 337010 496136 337016
rect 493968 4140 494020 4146
rect 493968 4082 494020 4088
rect 493876 4004 493928 4010
rect 493876 3946 493928 3952
rect 496096 3942 496124 337010
rect 496084 3936 496136 3942
rect 496084 3878 496136 3884
rect 496740 3874 496768 337554
rect 498120 337414 498148 340068
rect 498764 338026 498792 340068
rect 498752 338020 498804 338026
rect 498752 337962 498804 337968
rect 498844 337680 498896 337686
rect 498844 337622 498896 337628
rect 498108 337408 498160 337414
rect 498108 337350 498160 337356
rect 496728 3868 496780 3874
rect 496728 3810 496780 3816
rect 498856 3806 498884 337622
rect 497740 3800 497792 3806
rect 497740 3742 497792 3748
rect 498844 3800 498896 3806
rect 498844 3742 498896 3748
rect 495348 3732 495400 3738
rect 495348 3674 495400 3680
rect 494152 3596 494204 3602
rect 494152 3538 494204 3544
rect 493324 3188 493376 3194
rect 493324 3130 493376 3136
rect 494164 480 494192 3538
rect 495360 480 495388 3674
rect 496544 3188 496596 3194
rect 496544 3130 496596 3136
rect 496556 480 496584 3130
rect 497752 480 497780 3742
rect 499408 3602 499436 340068
rect 499488 338020 499540 338026
rect 499488 337962 499540 337968
rect 499500 3738 499528 337962
rect 499764 337884 499816 337890
rect 499764 337826 499816 337832
rect 499488 3732 499540 3738
rect 499488 3674 499540 3680
rect 499396 3596 499448 3602
rect 499396 3538 499448 3544
rect 498936 3528 498988 3534
rect 498936 3470 498988 3476
rect 498948 480 498976 3470
rect 499776 610 499804 337826
rect 499960 337754 499988 340068
rect 500618 340054 500908 340082
rect 499948 337748 500000 337754
rect 499948 337690 500000 337696
rect 500776 337748 500828 337754
rect 500776 337690 500828 337696
rect 500788 3670 500816 337690
rect 500776 3664 500828 3670
rect 500776 3606 500828 3612
rect 500880 3534 500908 340054
rect 501248 337890 501276 340068
rect 501814 340054 502288 340082
rect 501604 337952 501656 337958
rect 501604 337894 501656 337900
rect 501236 337884 501288 337890
rect 501236 337826 501288 337832
rect 500868 3528 500920 3534
rect 500868 3470 500920 3476
rect 501236 3460 501288 3466
rect 501236 3402 501288 3408
rect 499764 604 499816 610
rect 499764 546 499816 552
rect 500132 604 500184 610
rect 500132 546 500184 552
rect 500144 480 500172 546
rect 501248 480 501276 3402
rect 501616 3126 501644 337894
rect 502260 3466 502288 340054
rect 502444 337686 502472 340068
rect 503102 340054 503576 340082
rect 503444 337952 503496 337958
rect 503444 337894 503496 337900
rect 502616 337748 502668 337754
rect 502616 337690 502668 337696
rect 502432 337680 502484 337686
rect 502432 337622 502484 337628
rect 502248 3460 502300 3466
rect 502248 3402 502300 3408
rect 502432 3324 502484 3330
rect 502432 3266 502484 3272
rect 501604 3120 501656 3126
rect 501604 3062 501656 3068
rect 502444 480 502472 3266
rect 502628 3210 502656 337690
rect 503456 337006 503484 337894
rect 503548 337770 503576 340054
rect 503640 337958 503668 340068
rect 503628 337952 503680 337958
rect 503628 337894 503680 337900
rect 503548 337742 503668 337770
rect 504284 337754 504312 340068
rect 503536 337680 503588 337686
rect 503536 337622 503588 337628
rect 503444 337000 503496 337006
rect 503444 336942 503496 336948
rect 503548 4962 503576 337622
rect 503536 4956 503588 4962
rect 503536 4898 503588 4904
rect 503640 3584 503668 337742
rect 504272 337748 504324 337754
rect 504272 337690 504324 337696
rect 504928 336938 504956 340068
rect 505480 337754 505508 340068
rect 506138 340054 506336 340082
rect 505008 337748 505060 337754
rect 505008 337690 505060 337696
rect 505468 337748 505520 337754
rect 505468 337690 505520 337696
rect 504916 336932 504968 336938
rect 504916 336874 504968 336880
rect 503640 3556 503760 3584
rect 502628 3182 503668 3210
rect 503640 480 503668 3182
rect 503732 2854 503760 3556
rect 504824 3256 504876 3262
rect 504824 3198 504876 3204
rect 503720 2848 503772 2854
rect 503720 2790 503772 2796
rect 504836 480 504864 3198
rect 505020 2922 505048 337690
rect 506308 4826 506336 340054
rect 506768 337754 506796 340068
rect 506388 337748 506440 337754
rect 506388 337690 506440 337696
rect 506756 337748 506808 337754
rect 506756 337690 506808 337696
rect 506296 4820 506348 4826
rect 506296 4762 506348 4768
rect 506020 3120 506072 3126
rect 506020 3062 506072 3068
rect 505008 2916 505060 2922
rect 505008 2858 505060 2864
rect 506032 480 506060 3062
rect 506400 2990 506428 337690
rect 506664 337340 506716 337346
rect 506664 337282 506716 337288
rect 506388 2984 506440 2990
rect 506388 2926 506440 2932
rect 506676 610 506704 337282
rect 507320 337142 507348 340068
rect 507964 337754 507992 340068
rect 507768 337748 507820 337754
rect 507768 337690 507820 337696
rect 507952 337748 508004 337754
rect 507952 337690 508004 337696
rect 507308 337136 507360 337142
rect 507308 337078 507360 337084
rect 507780 3058 507808 337690
rect 508608 337278 508636 340068
rect 509160 338094 509188 340068
rect 509148 338088 509200 338094
rect 509148 338030 509200 338036
rect 509148 337748 509200 337754
rect 509148 337690 509200 337696
rect 508596 337272 508648 337278
rect 508596 337214 508648 337220
rect 509160 4894 509188 337690
rect 509804 337074 509832 340068
rect 510462 340054 510568 340082
rect 509884 337816 509936 337822
rect 509884 337758 509936 337764
rect 509792 337068 509844 337074
rect 509792 337010 509844 337016
rect 509148 4888 509200 4894
rect 509148 4830 509200 4836
rect 509608 4072 509660 4078
rect 509608 4014 509660 4020
rect 508412 3392 508464 3398
rect 508412 3334 508464 3340
rect 507768 3052 507820 3058
rect 507768 2994 507820 3000
rect 506664 604 506716 610
rect 506664 546 506716 552
rect 507216 604 507268 610
rect 507216 546 507268 552
rect 507228 480 507256 546
rect 508424 480 508452 3334
rect 509620 480 509648 4014
rect 509896 3942 509924 337758
rect 509884 3936 509936 3942
rect 509884 3878 509936 3884
rect 510540 3194 510568 340054
rect 511000 337754 511028 340068
rect 511658 340054 511856 340082
rect 510988 337748 511040 337754
rect 510988 337690 511040 337696
rect 510804 337612 510856 337618
rect 510804 337554 510856 337560
rect 510528 3188 510580 3194
rect 510528 3130 510580 3136
rect 510816 480 510844 337554
rect 511828 3262 511856 340054
rect 512288 337958 512316 340068
rect 512840 338026 512868 340068
rect 513498 340054 513880 340082
rect 512828 338020 512880 338026
rect 512828 337962 512880 337968
rect 512276 337952 512328 337958
rect 512276 337894 512328 337900
rect 511908 337748 511960 337754
rect 511908 337690 511960 337696
rect 511816 3256 511868 3262
rect 511816 3198 511868 3204
rect 511920 3126 511948 337690
rect 513852 337550 513880 340054
rect 514588 337736 514616 340190
rect 514680 337890 514708 340068
rect 514668 337884 514720 337890
rect 514668 337826 514720 337832
rect 514588 337708 514708 337736
rect 513564 337544 513616 337550
rect 513564 337486 513616 337492
rect 513840 337544 513892 337550
rect 513840 337486 513892 337492
rect 512000 4140 512052 4146
rect 512000 4082 512052 4088
rect 511908 3120 511960 3126
rect 511908 3062 511960 3068
rect 512012 480 512040 4082
rect 513196 4004 513248 4010
rect 513196 3946 513248 3952
rect 513208 480 513236 3946
rect 513576 610 513604 337486
rect 514576 134088 514628 134094
rect 514574 134056 514576 134065
rect 514628 134056 514630 134065
rect 514574 133991 514630 134000
rect 514576 40248 514628 40254
rect 514574 40216 514576 40225
rect 514628 40216 514630 40225
rect 514574 40151 514630 40160
rect 514574 16824 514630 16833
rect 514574 16759 514630 16768
rect 514588 16425 514616 16759
rect 514574 16416 514630 16425
rect 514574 16351 514630 16360
rect 514680 3330 514708 337708
rect 515324 337210 515352 340068
rect 515876 337822 515904 340068
rect 515864 337816 515916 337822
rect 515864 337758 515916 337764
rect 516520 337754 516548 340068
rect 516508 337748 516560 337754
rect 516508 337690 516560 337696
rect 516784 337680 516836 337686
rect 516784 337622 516836 337628
rect 515312 337204 515364 337210
rect 515312 337146 515364 337152
rect 514852 134088 514904 134094
rect 514850 134056 514852 134065
rect 514904 134056 514906 134065
rect 514850 133991 514906 134000
rect 514852 40248 514904 40254
rect 514850 40216 514852 40225
rect 514904 40216 514906 40225
rect 514850 40151 514906 40160
rect 516796 3874 516824 337622
rect 517164 337346 517192 340068
rect 517428 337748 517480 337754
rect 517428 337690 517480 337696
rect 517152 337340 517204 337346
rect 517152 337282 517204 337288
rect 515588 3868 515640 3874
rect 515588 3810 515640 3816
rect 516784 3868 516836 3874
rect 516784 3810 516836 3816
rect 514668 3324 514720 3330
rect 514668 3266 514720 3272
rect 513564 604 513616 610
rect 513564 546 513616 552
rect 514392 604 514444 610
rect 514392 546 514444 552
rect 514404 480 514432 546
rect 515600 480 515628 3810
rect 517440 3398 517468 337690
rect 517716 337618 517744 340068
rect 518360 337686 518388 340068
rect 518348 337680 518400 337686
rect 518348 337622 518400 337628
rect 519004 337618 519032 340068
rect 517704 337612 517756 337618
rect 517704 337554 517756 337560
rect 518808 337612 518860 337618
rect 518808 337554 518860 337560
rect 518992 337612 519044 337618
rect 518992 337554 519044 337560
rect 517612 337476 517664 337482
rect 517612 337418 517664 337424
rect 516784 3392 516836 3398
rect 516784 3334 516836 3340
rect 517428 3392 517480 3398
rect 517428 3334 517480 3340
rect 516796 480 516824 3334
rect 517624 626 517652 337418
rect 518820 4146 518848 337554
rect 519556 337482 519584 340068
rect 520096 337612 520148 337618
rect 520096 337554 520148 337560
rect 519544 337476 519596 337482
rect 519544 337418 519596 337424
rect 518808 4140 518860 4146
rect 518808 4082 518860 4088
rect 520108 4078 520136 337554
rect 520096 4072 520148 4078
rect 520096 4014 520148 4020
rect 520200 4010 520228 340068
rect 520844 337890 520872 340068
rect 521410 340054 521608 340082
rect 520832 337884 520884 337890
rect 520832 337826 520884 337832
rect 520372 337408 520424 337414
rect 520372 337350 520424 337356
rect 520188 4004 520240 4010
rect 520188 3946 520240 3952
rect 520280 3936 520332 3942
rect 520280 3878 520332 3884
rect 519084 3800 519136 3806
rect 519084 3742 519136 3748
rect 517624 598 517928 626
rect 517900 480 517928 598
rect 519096 480 519124 3742
rect 520292 480 520320 3878
rect 520384 610 520412 337350
rect 521580 3942 521608 340054
rect 522040 337618 522068 340068
rect 522698 340054 522988 340082
rect 522028 337612 522080 337618
rect 522028 337554 522080 337560
rect 521658 170368 521714 170377
rect 521658 170303 521714 170312
rect 521672 169833 521700 170303
rect 521658 169824 521714 169833
rect 521658 169759 521714 169768
rect 521658 22264 521714 22273
rect 521658 22199 521714 22208
rect 521672 22001 521700 22199
rect 521658 21992 521714 22001
rect 521658 21927 521714 21936
rect 521660 16720 521712 16726
rect 521658 16688 521660 16697
rect 521712 16688 521714 16697
rect 521658 16623 521714 16632
rect 521568 3936 521620 3942
rect 521568 3878 521620 3884
rect 522960 3806 522988 340054
rect 523236 337414 523264 340068
rect 523894 340054 524368 340082
rect 523224 337408 523276 337414
rect 523224 337350 523276 337356
rect 522948 3800 523000 3806
rect 522948 3742 523000 3748
rect 524340 3738 524368 340054
rect 524524 336802 524552 340068
rect 525090 340054 525564 340082
rect 524512 336796 524564 336802
rect 524512 336738 524564 336744
rect 524510 16960 524566 16969
rect 524510 16895 524566 16904
rect 524524 16726 524552 16895
rect 524512 16720 524564 16726
rect 524512 16662 524564 16668
rect 525064 3868 525116 3874
rect 525064 3810 525116 3816
rect 522672 3732 522724 3738
rect 522672 3674 522724 3680
rect 524328 3732 524380 3738
rect 524328 3674 524380 3680
rect 520372 604 520424 610
rect 520372 546 520424 552
rect 521476 604 521528 610
rect 521476 546 521528 552
rect 521488 480 521516 546
rect 522684 480 522712 3674
rect 523868 3596 523920 3602
rect 523868 3538 523920 3544
rect 523880 480 523908 3538
rect 525076 480 525104 3810
rect 525536 3670 525564 340054
rect 525616 336796 525668 336802
rect 525616 336738 525668 336744
rect 525628 3874 525656 336738
rect 525616 3868 525668 3874
rect 525616 3810 525668 3816
rect 525524 3664 525576 3670
rect 525524 3606 525576 3612
rect 525720 3369 525748 340068
rect 526378 340054 526852 340082
rect 526824 337210 526852 340054
rect 526916 337414 526944 340068
rect 526904 337408 526956 337414
rect 526904 337350 526956 337356
rect 526812 337204 526864 337210
rect 526812 337146 526864 337152
rect 527560 336802 527588 340068
rect 528204 337385 528232 340068
rect 528190 337376 528246 337385
rect 528190 337311 528246 337320
rect 528756 337210 528784 340068
rect 528744 337204 528796 337210
rect 528744 337146 528796 337152
rect 529400 336802 529428 340068
rect 527548 336796 527600 336802
rect 527548 336738 527600 336744
rect 528468 336796 528520 336802
rect 528468 336738 528520 336744
rect 529388 336796 529440 336802
rect 529388 336738 529440 336744
rect 527454 336560 527510 336569
rect 527454 336495 527510 336504
rect 527468 319025 527496 336495
rect 527454 319016 527510 319025
rect 527454 318951 527510 318960
rect 527638 309088 527694 309097
rect 527638 309023 527694 309032
rect 527652 302161 527680 309023
rect 527638 302152 527694 302161
rect 527638 302087 527694 302096
rect 527638 289776 527694 289785
rect 527638 289711 527694 289720
rect 527652 280401 527680 289711
rect 527638 280392 527694 280401
rect 527638 280327 527694 280336
rect 527454 270464 527510 270473
rect 527454 270399 527510 270408
rect 527468 261089 527496 270399
rect 527454 261080 527510 261089
rect 527454 261015 527510 261024
rect 527454 251152 527510 251161
rect 527454 251087 527510 251096
rect 527468 241777 527496 251087
rect 527454 241768 527510 241777
rect 527454 241703 527510 241712
rect 527638 231840 527694 231849
rect 527638 231775 527694 231784
rect 527652 222329 527680 231775
rect 527638 222320 527694 222329
rect 527638 222255 527694 222264
rect 527454 212528 527510 212537
rect 527454 212463 527510 212472
rect 527468 203153 527496 212463
rect 527454 203144 527510 203153
rect 527454 203079 527510 203088
rect 527454 193216 527510 193225
rect 527454 193151 527510 193160
rect 527468 183841 527496 193151
rect 527454 183832 527510 183841
rect 527454 183767 527510 183776
rect 527270 173904 527326 173913
rect 527270 173839 527326 173848
rect 527284 164257 527312 173839
rect 527270 164248 527326 164257
rect 527270 164183 527326 164192
rect 527270 154320 527326 154329
rect 527270 154255 527326 154264
rect 527284 144945 527312 154255
rect 527270 144936 527326 144945
rect 527270 144871 527326 144880
rect 527822 135144 527878 135153
rect 527822 135079 527878 135088
rect 527836 125633 527864 135079
rect 527822 125624 527878 125633
rect 527822 125559 527878 125568
rect 527454 96520 527510 96529
rect 527454 96455 527510 96464
rect 527468 87009 527496 96455
rect 527454 87000 527510 87009
rect 527454 86935 527510 86944
rect 527270 57760 527326 57769
rect 527270 57695 527326 57704
rect 527284 48385 527312 57695
rect 527270 48376 527326 48385
rect 527270 48311 527326 48320
rect 527454 38584 527510 38593
rect 527454 38519 527510 38528
rect 527468 29209 527496 38519
rect 527454 29200 527510 29209
rect 527454 29135 527510 29144
rect 527456 3596 527508 3602
rect 527456 3538 527508 3544
rect 526260 3528 526312 3534
rect 526260 3470 526312 3476
rect 525706 3360 525762 3369
rect 525706 3295 525762 3304
rect 526272 480 526300 3470
rect 527468 480 527496 3538
rect 528480 3534 528508 336738
rect 529492 64870 529520 640902
rect 529584 111790 529612 641038
rect 529662 638344 529718 638353
rect 529662 638279 529718 638288
rect 529676 158710 529704 638279
rect 529768 487150 529796 641378
rect 529860 534070 529888 641514
rect 530228 627910 530256 641582
rect 530306 638616 530362 638625
rect 530306 638551 530362 638560
rect 530216 627904 530268 627910
rect 530216 627846 530268 627852
rect 530320 604450 530348 638551
rect 530308 604444 530360 604450
rect 530308 604386 530360 604392
rect 530412 557530 530440 642738
rect 532148 642728 532200 642734
rect 532148 642670 532200 642676
rect 532056 642660 532108 642666
rect 532056 642602 532108 642608
rect 531044 642592 531096 642598
rect 531044 642534 531096 642540
rect 530676 642524 530728 642530
rect 530676 642466 530728 642472
rect 530492 641504 530544 641510
rect 530492 641446 530544 641452
rect 530400 557524 530452 557530
rect 530400 557466 530452 557472
rect 529848 534064 529900 534070
rect 529848 534006 529900 534012
rect 530504 510610 530532 641446
rect 530584 641164 530636 641170
rect 530584 641106 530636 641112
rect 530492 510604 530544 510610
rect 530492 510546 530544 510552
rect 529756 487144 529808 487150
rect 529756 487086 529808 487092
rect 529756 337204 529808 337210
rect 529756 337146 529808 337152
rect 529664 158704 529716 158710
rect 529664 158646 529716 158652
rect 529572 111784 529624 111790
rect 529572 111726 529624 111732
rect 529480 64864 529532 64870
rect 529480 64806 529532 64812
rect 529664 4956 529716 4962
rect 529664 4898 529716 4904
rect 528468 3528 528520 3534
rect 528468 3470 528520 3476
rect 528652 3460 528704 3466
rect 528652 3402 528704 3408
rect 528664 480 528692 3402
rect 529676 3346 529704 4898
rect 529768 3466 529796 337146
rect 529848 336796 529900 336802
rect 529848 336738 529900 336744
rect 529860 3602 529888 336738
rect 530596 205630 530624 641106
rect 530688 252550 530716 642466
rect 530952 641300 531004 641306
rect 530952 641242 531004 641248
rect 530768 641232 530820 641238
rect 530768 641174 530820 641180
rect 530780 264926 530808 641174
rect 530860 639872 530912 639878
rect 530860 639814 530912 639820
rect 530872 322930 530900 639814
rect 530964 346390 530992 641242
rect 531056 393310 531084 642534
rect 531964 641368 532016 641374
rect 531964 641310 532016 641316
rect 531136 640144 531188 640150
rect 531136 640086 531188 640092
rect 531148 416770 531176 640086
rect 531226 638480 531282 638489
rect 531226 638415 531282 638424
rect 531240 440230 531268 638415
rect 531228 440224 531280 440230
rect 531228 440166 531280 440172
rect 531136 416764 531188 416770
rect 531136 416706 531188 416712
rect 531976 405686 532004 641310
rect 532068 463690 532096 642602
rect 532160 499526 532188 642670
rect 532252 546446 532280 642806
rect 532344 593366 532372 642874
rect 532332 593360 532384 593366
rect 532332 593302 532384 593308
rect 532240 546440 532292 546446
rect 532240 546382 532292 546388
rect 532148 499520 532200 499526
rect 532148 499462 532200 499468
rect 532056 463684 532108 463690
rect 532056 463626 532108 463632
rect 531964 405680 532016 405686
rect 531964 405622 532016 405628
rect 531044 393304 531096 393310
rect 531044 393246 531096 393252
rect 530952 346384 531004 346390
rect 530952 346326 531004 346332
rect 542360 338088 542412 338094
rect 542360 338030 542412 338036
rect 540244 337272 540296 337278
rect 540244 337214 540296 337220
rect 538220 337136 538272 337142
rect 538220 337078 538272 337084
rect 534080 336932 534132 336938
rect 534080 336874 534132 336880
rect 531320 336796 531372 336802
rect 531320 336738 531372 336744
rect 530860 322924 530912 322930
rect 530860 322866 530912 322872
rect 530768 264920 530820 264926
rect 530768 264862 530820 264868
rect 530676 252544 530728 252550
rect 530676 252486 530728 252492
rect 530584 205624 530636 205630
rect 530584 205566 530636 205572
rect 529848 3596 529900 3602
rect 529848 3538 529900 3544
rect 529756 3460 529808 3466
rect 529756 3402 529808 3408
rect 531332 3346 531360 336738
rect 534092 3346 534120 336874
rect 536932 4820 536984 4826
rect 536932 4762 536984 4768
rect 529676 3318 529888 3346
rect 531332 3318 532280 3346
rect 534092 3318 534580 3346
rect 529860 480 529888 3318
rect 531044 2848 531096 2854
rect 531044 2790 531096 2796
rect 531056 480 531084 2790
rect 532252 480 532280 3318
rect 533436 2916 533488 2922
rect 533436 2858 533488 2864
rect 533448 480 533476 2858
rect 534552 480 534580 3318
rect 535736 2984 535788 2990
rect 535736 2926 535788 2932
rect 535748 480 535776 2926
rect 536944 480 536972 4762
rect 538232 3346 538260 337078
rect 538232 3318 539364 3346
rect 538128 3052 538180 3058
rect 538128 2994 538180 3000
rect 538140 480 538168 2994
rect 539336 480 539364 3318
rect 540256 3262 540284 337214
rect 540336 337068 540388 337074
rect 540336 337010 540388 337016
rect 540244 3256 540296 3262
rect 540244 3198 540296 3204
rect 540348 3194 540376 337010
rect 540886 170232 540942 170241
rect 540886 170167 540942 170176
rect 540900 169969 540928 170167
rect 540886 169960 540942 169969
rect 540886 169895 540942 169904
rect 540980 133952 541032 133958
rect 540978 133920 540980 133929
rect 541032 133920 541034 133929
rect 540978 133855 541034 133864
rect 540980 40112 541032 40118
rect 540978 40080 540980 40089
rect 541032 40080 541034 40089
rect 540978 40015 541034 40024
rect 540886 17232 540942 17241
rect 540886 17167 540942 17176
rect 540900 16833 540928 17167
rect 540886 16824 540942 16833
rect 540886 16759 540942 16768
rect 540520 4888 540572 4894
rect 540520 4830 540572 4836
rect 540336 3188 540388 3194
rect 540336 3130 540388 3136
rect 540532 480 540560 4830
rect 542372 3346 542400 338030
rect 547144 338020 547196 338026
rect 547144 337962 547196 337968
rect 545764 337000 545816 337006
rect 545764 336942 545816 336948
rect 543004 336864 543056 336870
rect 543004 336806 543056 336812
rect 542372 3318 542952 3346
rect 541716 3256 541768 3262
rect 541716 3198 541768 3204
rect 541728 480 541756 3198
rect 542924 480 542952 3318
rect 543016 2854 543044 336806
rect 544108 3188 544160 3194
rect 544108 3130 544160 3136
rect 543004 2848 543056 2854
rect 543004 2790 543056 2796
rect 544120 480 544148 3130
rect 545776 3126 545804 336942
rect 545854 134056 545910 134065
rect 545854 133991 545910 134000
rect 545868 133958 545896 133991
rect 545856 133952 545908 133958
rect 545856 133894 545908 133900
rect 545854 40216 545910 40225
rect 545854 40151 545910 40160
rect 545868 40118 545896 40151
rect 545856 40112 545908 40118
rect 545856 40054 545908 40060
rect 547156 3262 547184 337962
rect 547236 337952 547288 337958
rect 547236 337894 547288 337900
rect 547144 3256 547196 3262
rect 547144 3198 547196 3204
rect 545304 3120 545356 3126
rect 545304 3062 545356 3068
rect 545764 3120 545816 3126
rect 545764 3062 545816 3068
rect 545316 480 545344 3062
rect 547248 3058 547276 337894
rect 556804 337884 556856 337890
rect 556804 337826 556856 337832
rect 553400 337816 553452 337822
rect 553400 337758 553452 337764
rect 549904 337340 549956 337346
rect 549904 337282 549956 337288
rect 549916 3058 549944 337282
rect 553412 3346 553440 337758
rect 554872 337748 554924 337754
rect 554872 337690 554924 337696
rect 554502 134192 554558 134201
rect 554502 134127 554558 134136
rect 554516 133793 554544 134127
rect 554502 133784 554558 133793
rect 554502 133719 554558 133728
rect 554502 40352 554558 40361
rect 554502 40287 554558 40296
rect 554516 39953 554544 40287
rect 554502 39944 554558 39953
rect 554502 39879 554558 39888
rect 554884 3346 554912 337690
rect 552388 3324 552440 3330
rect 553412 3318 553624 3346
rect 554884 3318 556016 3346
rect 556816 3330 556844 337826
rect 560300 337680 560352 337686
rect 560300 337622 560352 337628
rect 558184 337204 558236 337210
rect 558184 337146 558236 337152
rect 558196 3398 558224 337146
rect 560206 170504 560262 170513
rect 560206 170439 560262 170448
rect 560220 170105 560248 170439
rect 560206 170096 560262 170105
rect 560206 170031 560262 170040
rect 560206 17368 560262 17377
rect 560206 17303 560262 17312
rect 560220 16969 560248 17303
rect 560206 16960 560262 16969
rect 560206 16895 560262 16904
rect 559564 4140 559616 4146
rect 559564 4082 559616 4088
rect 557172 3392 557224 3398
rect 557172 3334 557224 3340
rect 558184 3392 558236 3398
rect 558184 3334 558236 3340
rect 552388 3266 552440 3272
rect 550088 3256 550140 3262
rect 550088 3198 550140 3204
rect 546500 3052 546552 3058
rect 546500 2994 546552 3000
rect 547236 3052 547288 3058
rect 547236 2994 547288 3000
rect 548892 3052 548944 3058
rect 548892 2994 548944 3000
rect 549904 3052 549956 3058
rect 549904 2994 549956 3000
rect 546512 480 546540 2994
rect 547696 2984 547748 2990
rect 547696 2926 547748 2932
rect 547708 480 547736 2926
rect 548904 480 548932 2994
rect 550100 480 550128 3198
rect 551192 2984 551244 2990
rect 551192 2926 551244 2932
rect 551204 480 551232 2926
rect 552400 480 552428 3266
rect 553596 480 553624 3318
rect 554780 3120 554832 3126
rect 554780 3062 554832 3068
rect 554792 480 554820 3062
rect 555988 480 556016 3318
rect 556804 3324 556856 3330
rect 556804 3266 556856 3272
rect 557184 480 557212 3334
rect 558368 3256 558420 3262
rect 558368 3198 558420 3204
rect 558380 480 558408 3198
rect 559576 480 559604 4082
rect 560312 3482 560340 337622
rect 563152 337612 563204 337618
rect 563152 337554 563204 337560
rect 561956 4072 562008 4078
rect 561956 4014 562008 4020
rect 560312 3454 560800 3482
rect 560772 480 560800 3454
rect 561968 480 561996 4014
rect 563164 480 563192 337554
rect 567200 337544 567252 337550
rect 567200 337486 567252 337492
rect 565082 337376 565138 337385
rect 565082 337311 565138 337320
rect 565096 4010 565124 337311
rect 564348 4004 564400 4010
rect 564348 3946 564400 3952
rect 565084 4004 565136 4010
rect 565084 3946 565136 3952
rect 564360 480 564388 3946
rect 566740 3936 566792 3942
rect 566740 3878 566792 3884
rect 565544 3324 565596 3330
rect 565544 3266 565596 3272
rect 565556 480 565584 3266
rect 566752 480 566780 3878
rect 567212 3482 567240 337486
rect 569224 337476 569276 337482
rect 569224 337418 569276 337424
rect 569040 3800 569092 3806
rect 569040 3742 569092 3748
rect 567212 3454 567884 3482
rect 567856 480 567884 3454
rect 569052 480 569080 3742
rect 569236 3398 569264 337418
rect 571984 337408 572036 337414
rect 571984 337350 572036 337356
rect 571432 3732 571484 3738
rect 571432 3674 571484 3680
rect 569224 3392 569276 3398
rect 569224 3334 569276 3340
rect 570236 3392 570288 3398
rect 570236 3334 570288 3340
rect 570248 480 570276 3334
rect 571444 480 571472 3674
rect 571996 3058 572024 337350
rect 577516 218006 577544 670686
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 580908 642456 580960 642462
rect 580908 642398 580960 642404
rect 580632 642388 580684 642394
rect 580632 642330 580684 642336
rect 579802 642288 579858 642297
rect 579802 642223 579858 642232
rect 579618 639840 579674 639849
rect 579618 639775 579674 639784
rect 579632 639169 579660 639775
rect 579816 639198 579844 642223
rect 580356 641708 580408 641714
rect 580356 641650 580408 641656
rect 580080 641028 580132 641034
rect 580080 640970 580132 640976
rect 579896 640892 579948 640898
rect 579896 640834 579948 640840
rect 579804 639192 579856 639198
rect 579618 639160 579674 639169
rect 579804 639134 579856 639140
rect 579618 639095 579674 639104
rect 579804 627904 579856 627910
rect 579804 627846 579856 627852
rect 579816 627745 579844 627846
rect 579802 627736 579858 627745
rect 579802 627671 579858 627680
rect 579804 604444 579856 604450
rect 579804 604386 579856 604392
rect 579816 604217 579844 604386
rect 579802 604208 579858 604217
rect 579802 604143 579858 604152
rect 579804 593360 579856 593366
rect 579804 593302 579856 593308
rect 579816 592521 579844 593302
rect 579802 592512 579858 592521
rect 579802 592447 579858 592456
rect 579804 557524 579856 557530
rect 579804 557466 579856 557472
rect 579816 557297 579844 557466
rect 579802 557288 579858 557297
rect 579802 557223 579858 557232
rect 579804 546440 579856 546446
rect 579804 546382 579856 546388
rect 579816 545601 579844 546382
rect 579802 545592 579858 545601
rect 579802 545527 579858 545536
rect 579804 534064 579856 534070
rect 579804 534006 579856 534012
rect 579816 533905 579844 534006
rect 579802 533896 579858 533905
rect 579802 533831 579858 533840
rect 579804 510604 579856 510610
rect 579804 510546 579856 510552
rect 579816 510377 579844 510546
rect 579802 510368 579858 510377
rect 579802 510303 579858 510312
rect 579804 499520 579856 499526
rect 579804 499462 579856 499468
rect 579816 498681 579844 499462
rect 579802 498672 579858 498681
rect 579802 498607 579858 498616
rect 579804 487144 579856 487150
rect 579804 487086 579856 487092
rect 579816 486849 579844 487086
rect 579802 486840 579858 486849
rect 579802 486775 579858 486784
rect 579804 463684 579856 463690
rect 579804 463626 579856 463632
rect 579816 463457 579844 463626
rect 579802 463448 579858 463457
rect 579802 463383 579858 463392
rect 579908 451761 579936 640834
rect 579988 640212 580040 640218
rect 579988 640154 580040 640160
rect 579894 451752 579950 451761
rect 579894 451687 579950 451696
rect 579896 440224 579948 440230
rect 579896 440166 579948 440172
rect 579908 439929 579936 440166
rect 579894 439920 579950 439929
rect 579894 439855 579950 439864
rect 579896 416764 579948 416770
rect 579896 416706 579948 416712
rect 579908 416537 579936 416706
rect 579894 416528 579950 416537
rect 579894 416463 579950 416472
rect 579896 405680 579948 405686
rect 579896 405622 579948 405628
rect 579908 404841 579936 405622
rect 579894 404832 579950 404841
rect 579894 404767 579950 404776
rect 579896 393304 579948 393310
rect 579896 393246 579948 393252
rect 579908 393009 579936 393246
rect 579894 393000 579950 393009
rect 579894 392935 579950 392944
rect 580000 369617 580028 640154
rect 579986 369608 580042 369617
rect 579986 369543 580042 369552
rect 580092 357921 580120 640970
rect 580172 640076 580224 640082
rect 580172 640018 580224 640024
rect 580184 639441 580212 640018
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580368 639282 580396 641650
rect 580540 639940 580592 639946
rect 580540 639882 580592 639888
rect 580184 639254 580396 639282
rect 580446 639296 580502 639305
rect 580078 357912 580134 357921
rect 580078 357847 580134 357856
rect 579804 346384 579856 346390
rect 579804 346326 579856 346332
rect 579816 346089 579844 346326
rect 579802 346080 579858 346089
rect 579802 346015 579858 346024
rect 580080 322924 580132 322930
rect 580080 322866 580132 322872
rect 580092 322697 580120 322866
rect 580078 322688 580134 322697
rect 580078 322623 580134 322632
rect 580184 310865 580212 639254
rect 580446 639231 580502 639240
rect 580356 639192 580408 639198
rect 580262 639160 580318 639169
rect 580356 639134 580408 639140
rect 580262 639095 580318 639104
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 579620 252544 579672 252550
rect 579620 252486 579672 252492
rect 579632 252249 579660 252486
rect 579618 252240 579674 252249
rect 579618 252175 579674 252184
rect 577504 218000 577556 218006
rect 577504 217942 577556 217948
rect 579620 218000 579672 218006
rect 579620 217942 579672 217948
rect 579632 217025 579660 217942
rect 579618 217016 579674 217025
rect 579618 216951 579674 216960
rect 580172 205624 580224 205630
rect 580172 205566 580224 205572
rect 580184 205329 580212 205566
rect 580170 205320 580226 205329
rect 580170 205255 580226 205264
rect 572626 169960 572682 169969
rect 572626 169895 572682 169904
rect 572640 169810 572668 169895
rect 572718 169824 572774 169833
rect 572640 169782 572718 169810
rect 572718 169759 572774 169768
rect 579712 158704 579764 158710
rect 579712 158646 579764 158652
rect 579724 158409 579752 158646
rect 579710 158400 579766 158409
rect 579710 158335 579766 158344
rect 572626 134056 572682 134065
rect 572626 133991 572682 134000
rect 572640 133906 572668 133991
rect 572718 133920 572774 133929
rect 572640 133878 572718 133906
rect 572718 133855 572774 133864
rect 580172 111784 580224 111790
rect 580172 111726 580224 111732
rect 580184 111489 580212 111726
rect 580170 111480 580226 111489
rect 580170 111415 580226 111424
rect 580172 64864 580224 64870
rect 580172 64806 580224 64812
rect 580184 64569 580212 64806
rect 580170 64560 580226 64569
rect 580170 64495 580226 64504
rect 572626 40216 572682 40225
rect 572626 40151 572682 40160
rect 572640 40066 572668 40151
rect 572718 40080 572774 40089
rect 572640 40038 572718 40066
rect 572718 40015 572774 40024
rect 580276 29345 580304 639095
rect 580368 87961 580396 639134
rect 580354 87952 580410 87961
rect 580354 87887 580410 87896
rect 580460 76265 580488 639231
rect 580552 123185 580580 639882
rect 580644 181937 580672 642330
rect 580724 640280 580776 640286
rect 580724 640222 580776 640228
rect 580736 228857 580764 640222
rect 580816 639804 580868 639810
rect 580816 639746 580868 639752
rect 580828 275777 580856 639746
rect 580920 299169 580948 642398
rect 580906 299160 580962 299169
rect 580906 299095 580962 299104
rect 580814 275768 580870 275777
rect 580814 275703 580870 275712
rect 580722 228848 580778 228857
rect 580722 228783 580778 228792
rect 580630 181928 580686 181937
rect 580630 181863 580686 181872
rect 580538 123176 580594 123185
rect 580538 123111 580594 123120
rect 580446 76256 580502 76265
rect 580446 76191 580502 76200
rect 580262 29336 580318 29345
rect 580262 29271 580318 29280
rect 572626 16824 572682 16833
rect 572626 16759 572682 16768
rect 572640 16674 572668 16759
rect 572718 16688 572774 16697
rect 572640 16646 572718 16674
rect 572718 16623 572774 16632
rect 579804 4004 579856 4010
rect 579804 3946 579856 3952
rect 572628 3868 572680 3874
rect 572628 3810 572680 3816
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572640 480 572668 3810
rect 573824 3664 573876 3670
rect 573824 3606 573876 3612
rect 573836 480 573864 3606
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 575018 3360 575074 3369
rect 575018 3295 575074 3304
rect 575032 480 575060 3295
rect 576216 3256 576268 3262
rect 576216 3198 576268 3204
rect 576228 480 576256 3198
rect 577412 3052 577464 3058
rect 577412 2994 577464 3000
rect 577424 480 577452 2994
rect 578620 480 578648 3470
rect 579816 480 579844 3946
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3514 643048 3570 643104
rect 3238 624860 3240 624880
rect 3240 624860 3292 624880
rect 3292 624860 3294 624880
rect 3238 624824 3294 624860
rect 2778 610408 2834 610464
rect 3238 596028 3240 596048
rect 3240 596028 3292 596048
rect 3292 596028 3294 596048
rect 3238 595992 3294 596028
rect 3238 567296 3294 567352
rect 2778 553052 2780 553072
rect 2780 553052 2832 553072
rect 2832 553052 2834 553072
rect 2778 553016 2834 553052
rect 3238 538600 3294 538656
rect 3238 509904 3294 509960
rect 2778 495488 2834 495544
rect 3238 481108 3240 481128
rect 3240 481108 3292 481128
rect 3292 481108 3294 481128
rect 3238 481072 3294 481108
rect 3146 452412 3148 452432
rect 3148 452412 3200 452432
rect 3200 452412 3202 452432
rect 3146 452376 3202 452412
rect 3146 437960 3202 438016
rect 3422 639512 3478 639568
rect 3330 423680 3386 423736
rect 3146 394984 3202 395040
rect 2778 380604 2780 380624
rect 2780 380604 2832 380624
rect 2832 380604 2834 380624
rect 2778 380568 2834 380604
rect 3330 366152 3386 366208
rect 3238 337456 3294 337512
rect 2778 323040 2834 323096
rect 3330 294380 3332 294400
rect 3332 294380 3384 294400
rect 3384 294380 3386 294400
rect 3330 294344 3386 294380
rect 3146 280100 3148 280120
rect 3148 280100 3200 280120
rect 3200 280100 3202 280120
rect 3146 280064 3202 280100
rect 3330 265648 3386 265704
rect 3146 252456 3202 252512
rect 3146 251232 3202 251288
rect 2778 236952 2834 237008
rect 3146 193840 3202 193896
rect 2778 179460 2780 179480
rect 2780 179460 2832 179480
rect 2832 179460 2834 179480
rect 2778 179424 2834 179460
rect 2778 78920 2834 78976
rect 259918 642912 259974 642968
rect 258722 642776 258778 642832
rect 4894 641960 4950 642016
rect 3698 641824 3754 641880
rect 3606 638968 3662 639024
rect 3606 107616 3662 107672
rect 3882 639648 3938 639704
rect 3790 638152 3846 638208
rect 4158 639784 4214 639840
rect 4066 222536 4122 222592
rect 3974 150728 4030 150784
rect 3882 136312 3938 136368
rect 3790 122032 3846 122088
rect 3698 93200 3754 93256
rect 3514 64504 3570 64560
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 4066 7112 4122 7168
rect 72422 642096 72478 642152
rect 5538 639532 5594 639568
rect 5538 639512 5540 639532
rect 5540 639512 5592 639532
rect 5592 639512 5594 639532
rect 6182 639104 6238 639160
rect 41602 641552 41658 641608
rect 53102 641552 53158 641608
rect 60922 641552 60978 641608
rect 68466 641552 68522 641608
rect 41602 640872 41658 640928
rect 53102 640872 53158 640928
rect 60922 640872 60978 640928
rect 68466 640872 68522 640928
rect 23386 639512 23442 639568
rect 50802 639376 50858 639432
rect 51078 639376 51134 639432
rect 60646 639376 60702 639432
rect 70122 639376 70178 639432
rect 70398 639376 70454 639432
rect 66166 639260 66222 639296
rect 66166 639240 66168 639260
rect 66168 639240 66220 639260
rect 66220 639240 66222 639260
rect 10322 337320 10378 337376
rect 6458 3304 6514 3360
rect 48134 6160 48190 6216
rect 60646 10240 60702 10296
rect 79966 639376 80022 639432
rect 80150 639376 80206 639432
rect 91742 641552 91798 641608
rect 99562 641552 99618 641608
rect 118882 641552 118938 641608
rect 130382 641552 130438 641608
rect 146114 641552 146170 641608
rect 157522 641552 157578 641608
rect 176842 641552 176898 641608
rect 188342 641552 188398 641608
rect 193954 641552 194010 641608
rect 207662 641552 207718 641608
rect 91742 640872 91798 640928
rect 99562 640872 99618 640928
rect 118882 640872 118938 640928
rect 130382 640872 130438 640928
rect 146114 640872 146170 640928
rect 157522 640872 157578 640928
rect 176842 640872 176898 640928
rect 188342 640872 188398 640928
rect 193954 640872 194010 640928
rect 207662 640872 207718 640928
rect 109682 639784 109738 639840
rect 119342 639784 119398 639840
rect 162858 639784 162914 639840
rect 177302 639784 177358 639840
rect 89442 639376 89498 639432
rect 89718 639376 89774 639432
rect 147770 639512 147826 639568
rect 156326 639532 156382 639568
rect 156326 639512 156328 639532
rect 156328 639512 156380 639532
rect 156380 639512 156382 639532
rect 119342 639376 119398 639432
rect 147586 639376 147642 639432
rect 186318 639512 186374 639568
rect 177302 639376 177358 639432
rect 186042 639376 186098 639432
rect 220818 639512 220874 639568
rect 201498 639376 201554 639432
rect 109682 639240 109738 639296
rect 211066 639240 211122 639296
rect 136086 8880 136142 8936
rect 134890 7520 134946 7576
rect 219346 4800 219402 4856
rect 231398 639920 231454 639976
rect 241518 642232 241574 642288
rect 243542 641552 243598 641608
rect 243542 640872 243598 640928
rect 244186 640056 244242 640112
rect 275282 641552 275338 641608
rect 275282 640872 275338 640928
rect 233974 639784 234030 639840
rect 235262 639784 235318 639840
rect 249522 639784 249578 639840
rect 254950 639784 255006 639840
rect 302054 640056 302110 640112
rect 325698 642912 325754 642968
rect 328182 639920 328238 639976
rect 290002 639784 290058 639840
rect 340786 639784 340842 639840
rect 340970 639784 341026 639840
rect 414018 700304 414074 700360
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 520462 643048 520518 643104
rect 429014 642096 429070 642152
rect 340786 639648 340842 639704
rect 340970 639648 341026 639704
rect 463422 640056 463478 640112
rect 463238 639920 463294 639976
rect 471058 639920 471114 639976
rect 504638 642776 504694 642832
rect 483662 642640 483718 642696
rect 491482 642504 491538 642560
rect 499394 642368 499450 642424
rect 494150 641960 494206 642016
rect 507306 642096 507362 642152
rect 509974 641824 510030 641880
rect 515862 641688 515918 641744
rect 515862 640192 515918 640248
rect 525706 641688 525762 641744
rect 462962 639648 463018 639704
rect 463238 639648 463294 639704
rect 463422 639648 463478 639704
rect 470138 639648 470194 639704
rect 471058 639648 471114 639704
rect 485134 639648 485190 639704
rect 496634 639648 496690 639704
rect 512274 639648 512330 639704
rect 528098 639648 528154 639704
rect 232410 337320 232466 337376
rect 230662 231784 230718 231840
rect 230846 231784 230902 231840
rect 231766 220768 231822 220824
rect 231950 220768 232006 220824
rect 230662 212472 230718 212528
rect 230846 212472 230902 212528
rect 230662 193160 230718 193216
rect 230846 193160 230902 193216
rect 230662 154536 230718 154592
rect 230846 154556 230902 154592
rect 230846 154536 230848 154556
rect 230848 154536 230900 154556
rect 230900 154536 230902 154556
rect 230754 144880 230810 144936
rect 231030 144880 231086 144936
rect 231950 143540 232006 143576
rect 231950 143520 231952 143540
rect 231952 143520 232004 143540
rect 232004 143520 232006 143540
rect 232226 143520 232282 143576
rect 230754 125568 230810 125624
rect 231030 125568 231086 125624
rect 230754 106256 230810 106312
rect 231030 106256 231086 106312
rect 231950 86944 232006 87000
rect 232226 86944 232282 87000
rect 231950 3304 232006 3360
rect 236458 288360 236514 288416
rect 236642 288360 236698 288416
rect 236274 230424 236330 230480
rect 236458 230424 236514 230480
rect 236274 211112 236330 211168
rect 236550 211112 236606 211168
rect 236274 106256 236330 106312
rect 236458 106256 236514 106312
rect 236366 96600 236422 96656
rect 236550 96600 236606 96656
rect 236366 87080 236422 87136
rect 236274 86944 236330 87000
rect 238758 170332 238814 170368
rect 238758 170312 238760 170332
rect 238760 170312 238812 170332
rect 238812 170312 238814 170332
rect 240138 164212 240194 164248
rect 240138 164192 240140 164212
rect 240140 164192 240192 164212
rect 240192 164192 240194 164212
rect 240322 164212 240378 164248
rect 240322 164192 240324 164212
rect 240324 164192 240376 164212
rect 240376 164192 240378 164212
rect 240138 143656 240194 143712
rect 240138 143520 240194 143576
rect 242806 270544 242862 270600
rect 242806 251232 242862 251288
rect 241794 183504 241850 183560
rect 241978 183504 242034 183560
rect 241794 115912 241850 115968
rect 241978 115912 242034 115968
rect 241794 96600 241850 96656
rect 241978 96600 242034 96656
rect 243542 327256 243598 327312
rect 243082 327120 243138 327176
rect 243174 270408 243230 270464
rect 242990 251096 243046 251152
rect 242990 241476 242992 241496
rect 242992 241476 243044 241496
rect 243044 241476 243046 241496
rect 242990 241440 243046 241476
rect 243174 241476 243176 241496
rect 243176 241476 243228 241496
rect 243228 241476 243230 241496
rect 243174 241440 243230 241476
rect 244462 182144 244518 182200
rect 244646 182144 244702 182200
rect 243174 171128 243230 171184
rect 243358 171128 243414 171184
rect 243266 77424 243322 77480
rect 243082 75928 243138 75984
rect 244186 16768 244242 16824
rect 244370 16768 244426 16824
rect 248326 170040 248382 170096
rect 249246 307672 249302 307728
rect 249246 298288 249302 298344
rect 249246 279792 249302 279848
rect 249246 270544 249302 270600
rect 249246 270408 249302 270464
rect 249246 260888 249302 260944
rect 249246 251096 249302 251152
rect 249246 241712 249302 241768
rect 249430 222128 249486 222184
rect 249430 214512 249486 214568
rect 249522 199824 249578 199880
rect 249522 185544 249578 185600
rect 249614 179288 249670 179344
rect 249614 169904 249670 169960
rect 252466 212472 252522 212528
rect 252558 154536 252614 154592
rect 252558 135224 252614 135280
rect 252742 231784 252798 231840
rect 252926 231784 252982 231840
rect 252742 212508 252744 212528
rect 252744 212508 252796 212528
rect 252796 212508 252798 212528
rect 252742 212472 252798 212508
rect 252742 154536 252798 154592
rect 252742 135224 252798 135280
rect 252742 115912 252798 115968
rect 252926 115912 252982 115968
rect 255594 315968 255650 316024
rect 255778 315968 255834 316024
rect 254306 296656 254362 296712
rect 254490 296656 254546 296712
rect 254030 259392 254086 259448
rect 254214 259392 254270 259448
rect 254030 241476 254032 241496
rect 254032 241476 254084 241496
rect 254084 241476 254086 241496
rect 254030 241440 254086 241476
rect 254214 241476 254216 241496
rect 254216 241476 254268 241496
rect 254268 241476 254270 241496
rect 254214 241440 254270 241476
rect 254122 193196 254124 193216
rect 254124 193196 254176 193216
rect 254176 193196 254178 193216
rect 254122 193160 254178 193196
rect 254306 193196 254308 193216
rect 254308 193196 254360 193216
rect 254360 193196 254362 193216
rect 254306 193160 254362 193196
rect 254306 154536 254362 154592
rect 254306 154400 254362 154456
rect 254122 135224 254178 135280
rect 254306 135224 254362 135280
rect 254122 115932 254178 115968
rect 254122 115912 254124 115932
rect 254124 115912 254176 115932
rect 254176 115912 254178 115932
rect 254306 115912 254362 115968
rect 253938 6160 253994 6216
rect 259366 277344 259422 277400
rect 259366 170312 259422 170368
rect 259366 169904 259422 169960
rect 261022 318960 261078 319016
rect 261022 318824 261078 318880
rect 261022 307672 261078 307728
rect 261206 307672 261262 307728
rect 259734 277344 259790 277400
rect 259550 259392 259606 259448
rect 259734 259392 259790 259448
rect 259550 241476 259552 241496
rect 259552 241476 259604 241496
rect 259604 241476 259606 241496
rect 259550 241440 259606 241476
rect 259734 241476 259736 241496
rect 259736 241476 259788 241496
rect 259788 241476 259790 241496
rect 259734 241440 259790 241476
rect 259642 182280 259698 182336
rect 259734 182164 259790 182200
rect 259734 182144 259736 182164
rect 259736 182144 259788 182164
rect 259788 182144 259790 182164
rect 259642 172488 259698 172544
rect 259918 172488 259974 172544
rect 259642 135244 259698 135280
rect 259642 135224 259644 135244
rect 259644 135224 259696 135244
rect 259696 135224 259698 135244
rect 259826 135244 259882 135280
rect 259826 135224 259828 135244
rect 259828 135224 259880 135244
rect 259880 135224 259882 135244
rect 259642 115932 259698 115968
rect 259642 115912 259644 115932
rect 259644 115912 259696 115932
rect 259696 115912 259698 115932
rect 259826 115932 259882 115968
rect 259826 115912 259828 115932
rect 259828 115912 259880 115932
rect 259880 115912 259882 115932
rect 259642 96600 259698 96656
rect 259826 96600 259882 96656
rect 259826 10240 259882 10296
rect 265162 269048 265218 269104
rect 265438 269048 265494 269104
rect 265162 230424 265218 230480
rect 265346 230424 265402 230480
rect 266358 202816 266414 202872
rect 266542 202816 266598 202872
rect 267002 183504 267058 183560
rect 267186 183504 267242 183560
rect 265162 164328 265218 164384
rect 265254 164192 265310 164248
rect 267738 169924 267794 169960
rect 267738 169904 267740 169924
rect 267740 169904 267792 169924
rect 267792 169904 267794 169924
rect 265254 143520 265310 143576
rect 265438 143384 265494 143440
rect 265162 115932 265218 115968
rect 265162 115912 265164 115932
rect 265164 115912 265216 115932
rect 265216 115912 265218 115932
rect 265346 115912 265402 115968
rect 266726 115912 266782 115968
rect 267094 115912 267150 115968
rect 267278 115912 267334 115968
rect 266542 115776 266598 115832
rect 269026 17176 269082 17232
rect 269026 16768 269082 16824
rect 270406 182144 270462 182200
rect 270774 260752 270830 260808
rect 270590 260616 270646 260672
rect 270590 203088 270646 203144
rect 270774 202952 270830 203008
rect 271970 183504 272026 183560
rect 272246 183368 272302 183424
rect 270590 182164 270646 182200
rect 270590 182144 270592 182164
rect 270592 182144 270644 182164
rect 270644 182144 270646 182164
rect 270682 172488 270738 172544
rect 270866 172488 270922 172544
rect 272062 164212 272118 164248
rect 272062 164192 272064 164212
rect 272064 164192 272116 164212
rect 272116 164192 272118 164212
rect 272246 164212 272302 164248
rect 272246 164192 272248 164212
rect 272248 164192 272300 164212
rect 272300 164192 272302 164212
rect 270866 154672 270922 154728
rect 270682 154556 270738 154592
rect 270682 154536 270684 154556
rect 270684 154536 270736 154556
rect 270736 154536 270738 154556
rect 272062 154556 272118 154592
rect 272062 154536 272064 154556
rect 272064 154536 272116 154556
rect 272116 154536 272118 154556
rect 272246 154536 272302 154592
rect 271786 144880 271842 144936
rect 271970 144900 272026 144936
rect 271970 144880 271972 144900
rect 271972 144880 272024 144900
rect 272024 144880 272026 144900
rect 270682 135244 270738 135280
rect 270682 135224 270684 135244
rect 270684 135224 270736 135244
rect 270736 135224 270738 135244
rect 270866 135224 270922 135280
rect 273074 40296 273130 40352
rect 273258 40296 273314 40352
rect 277674 335280 277730 335336
rect 277950 335280 278006 335336
rect 277674 325624 277730 325680
rect 277858 325624 277914 325680
rect 278686 169768 278742 169824
rect 277398 154536 277454 154592
rect 277674 154536 277730 154592
rect 278778 16924 278834 16960
rect 278778 16904 278780 16924
rect 278780 16904 278832 16924
rect 278832 16904 278834 16924
rect 277490 8472 277546 8528
rect 277582 8336 277638 8392
rect 281630 289720 281686 289776
rect 281906 289720 281962 289776
rect 281722 280064 281778 280120
rect 281814 279928 281870 279984
rect 281814 260752 281870 260808
rect 281998 260752 282054 260808
rect 282918 241440 282974 241496
rect 283102 241440 283158 241496
rect 281722 211132 281778 211168
rect 281722 211112 281724 211132
rect 281724 211112 281776 211132
rect 281776 211112 281778 211132
rect 281906 211112 281962 211168
rect 282918 183504 282974 183560
rect 283102 183504 283158 183560
rect 283470 169904 283526 169960
rect 283470 169496 283526 169552
rect 281630 143520 281686 143576
rect 281814 143520 281870 143576
rect 281814 67632 281870 67688
rect 281998 67632 282054 67688
rect 284298 134036 284300 134056
rect 284300 134036 284352 134056
rect 284352 134036 284354 134056
rect 284298 134000 284354 134036
rect 287242 231784 287298 231840
rect 287426 231784 287482 231840
rect 287242 193160 287298 193216
rect 287426 193160 287482 193216
rect 287242 154536 287298 154592
rect 287426 154536 287482 154592
rect 289634 169940 289636 169960
rect 289636 169940 289688 169960
rect 289688 169940 289690 169960
rect 289634 169904 289690 169940
rect 289818 40160 289874 40216
rect 289818 40024 289874 40080
rect 288346 16632 288402 16688
rect 292486 55256 292542 55312
rect 292946 170040 293002 170096
rect 293774 134272 293830 134328
rect 292762 55256 292818 55312
rect 294050 335280 294106 335336
rect 294326 335280 294382 335336
rect 294142 201592 294198 201648
rect 294142 201456 294198 201512
rect 295246 134272 295302 134328
rect 295246 133864 295302 133920
rect 295430 190440 295486 190496
rect 295614 190440 295670 190496
rect 295706 131280 295762 131336
rect 295522 131144 295578 131200
rect 298282 278704 298338 278760
rect 298558 278704 298614 278760
rect 298190 170040 298246 170096
rect 298190 169904 298246 169960
rect 299294 16632 299350 16688
rect 299294 16496 299350 16552
rect 298282 7520 298338 7576
rect 299570 8880 299626 8936
rect 302146 40044 302202 40080
rect 302146 40024 302148 40044
rect 302148 40024 302200 40044
rect 302200 40024 302202 40044
rect 305182 241440 305238 241496
rect 305366 241440 305422 241496
rect 305182 222128 305238 222184
rect 305366 222128 305422 222184
rect 305182 202816 305238 202872
rect 305366 202816 305422 202872
rect 305182 183504 305238 183560
rect 305366 183504 305422 183560
rect 307298 40160 307354 40216
rect 308034 183504 308090 183560
rect 308310 183504 308366 183560
rect 308034 154536 308090 154592
rect 308310 154536 308366 154592
rect 308126 135224 308182 135280
rect 308310 135224 308366 135280
rect 308034 115912 308090 115968
rect 308310 115912 308366 115968
rect 308034 96600 308090 96656
rect 308218 96600 308274 96656
rect 309046 16768 309102 16824
rect 309046 16360 309102 16416
rect 309414 299376 309470 299432
rect 309598 299376 309654 299432
rect 309414 280064 309470 280120
rect 309598 280064 309654 280120
rect 309322 251096 309378 251152
rect 309506 251096 309562 251152
rect 309230 183776 309286 183832
rect 309414 183640 309470 183696
rect 310426 28872 310482 28928
rect 310702 241440 310758 241496
rect 310886 241440 310942 241496
rect 310702 222128 310758 222184
rect 310886 222128 310942 222184
rect 310702 202816 310758 202872
rect 310886 202816 310942 202872
rect 310702 154536 310758 154592
rect 310886 154536 310942 154592
rect 310702 135224 310758 135280
rect 310886 135224 310942 135280
rect 310702 48456 310758 48512
rect 310610 48320 310666 48376
rect 310610 28872 310666 28928
rect 314566 134408 314622 134464
rect 314566 134136 314622 134192
rect 317510 170040 317566 170096
rect 317510 169768 317566 169824
rect 324226 318688 324282 318744
rect 324226 182144 324282 182200
rect 324226 171128 324282 171184
rect 324226 122712 324282 122768
rect 323582 16904 323638 16960
rect 323490 16768 323546 16824
rect 324410 318688 324466 318744
rect 324502 289720 324558 289776
rect 324686 289720 324742 289776
rect 324502 182144 324558 182200
rect 324410 171128 324466 171184
rect 325606 133884 325662 133920
rect 325606 133864 325608 133884
rect 325608 133864 325660 133884
rect 325660 133864 325662 133884
rect 324410 122712 324466 122768
rect 324502 95240 324558 95296
rect 324686 95240 324742 95296
rect 326066 169804 326068 169824
rect 326068 169804 326120 169824
rect 326120 169804 326122 169824
rect 326066 169768 326122 169804
rect 327446 328616 327502 328672
rect 327170 328480 327226 328536
rect 327170 124208 327226 124264
rect 327170 123936 327226 123992
rect 331126 270544 331182 270600
rect 331126 251232 331182 251288
rect 331126 251096 331182 251152
rect 331126 209752 331182 209808
rect 331310 270408 331366 270464
rect 331494 209752 331550 209808
rect 330206 135224 330262 135280
rect 329930 135088 329986 135144
rect 329930 45600 329986 45656
rect 330114 45464 330170 45520
rect 331494 172624 331550 172680
rect 331402 172488 331458 172544
rect 331310 170040 331366 170096
rect 332690 328344 332746 328400
rect 332782 318824 332838 318880
rect 333886 133884 333942 133920
rect 333886 133864 333888 133884
rect 333888 133864 333940 133884
rect 333940 133864 333942 133884
rect 335266 40160 335322 40216
rect 335266 40024 335322 40080
rect 335266 17176 335322 17232
rect 335266 16768 335322 16824
rect 338026 170040 338082 170096
rect 338026 169632 338082 169688
rect 342442 251096 342498 251152
rect 342626 251096 342682 251152
rect 342442 231784 342498 231840
rect 342718 231784 342774 231840
rect 342718 212744 342774 212800
rect 342442 212506 342498 212562
rect 342718 191800 342774 191856
rect 342902 191800 342958 191856
rect 342442 172488 342498 172544
rect 342718 172488 342774 172544
rect 342350 154672 342406 154728
rect 342442 154536 342498 154592
rect 342350 144880 342406 144936
rect 342534 144880 342590 144936
rect 342534 116048 342590 116104
rect 342442 115932 342498 115968
rect 342442 115912 342444 115932
rect 342444 115912 342496 115932
rect 342496 115912 342498 115932
rect 342258 4800 342314 4856
rect 344926 40296 344982 40352
rect 344926 40024 344982 40080
rect 346214 16632 346270 16688
rect 346214 16496 346270 16552
rect 346582 241440 346638 241496
rect 346766 241440 346822 241496
rect 346582 222128 346638 222184
rect 346766 222128 346822 222184
rect 346582 202816 346638 202872
rect 346766 202816 346822 202872
rect 346582 183504 346638 183560
rect 346766 183504 346822 183560
rect 346582 154536 346638 154592
rect 346766 154536 346822 154592
rect 346582 135224 346638 135280
rect 346766 135224 346822 135280
rect 347686 16668 347688 16688
rect 347688 16668 347740 16688
rect 347740 16668 347742 16688
rect 347686 16632 347742 16668
rect 347870 277344 347926 277400
rect 348054 277344 348110 277400
rect 347962 193196 347964 193216
rect 347964 193196 348016 193216
rect 348016 193196 348018 193216
rect 347962 193160 348018 193196
rect 348146 193196 348148 193216
rect 348148 193196 348200 193216
rect 348200 193196 348202 193216
rect 348146 193160 348202 193196
rect 348422 133592 348478 133648
rect 348054 116048 348110 116104
rect 347962 115932 348018 115968
rect 347962 115912 347964 115932
rect 347964 115912 348016 115932
rect 348016 115912 348018 115932
rect 347962 87080 348018 87136
rect 347870 86944 347926 87000
rect 351826 144880 351882 144936
rect 352102 269048 352158 269104
rect 352286 269048 352342 269104
rect 352010 202852 352012 202872
rect 352012 202852 352064 202872
rect 352064 202852 352066 202872
rect 352010 202816 352066 202852
rect 352102 202680 352158 202736
rect 352102 164192 352158 164248
rect 352010 164056 352066 164112
rect 352010 144900 352066 144936
rect 352010 144880 352012 144900
rect 352012 144880 352064 144900
rect 352064 144880 352066 144900
rect 352010 125588 352066 125624
rect 352010 125568 352012 125588
rect 352012 125568 352064 125588
rect 352064 125568 352066 125588
rect 352194 125588 352250 125624
rect 352194 125568 352196 125588
rect 352196 125568 352248 125588
rect 352248 125568 352250 125588
rect 352102 87080 352158 87136
rect 352010 86964 352066 87000
rect 352010 86944 352012 86964
rect 352012 86944 352064 86964
rect 352064 86944 352066 86964
rect 353482 193196 353484 193216
rect 353484 193196 353536 193216
rect 353536 193196 353538 193216
rect 353482 193160 353538 193196
rect 353666 193196 353668 193216
rect 353668 193196 353720 193216
rect 353720 193196 353722 193216
rect 353666 193160 353722 193196
rect 353482 173884 353484 173904
rect 353484 173884 353536 173904
rect 353536 173884 353538 173904
rect 353482 173848 353538 173884
rect 353574 173712 353630 173768
rect 354586 133592 354642 133648
rect 355966 170176 356022 170232
rect 355966 169496 356022 169552
rect 355966 16904 356022 16960
rect 356426 173884 356428 173904
rect 356428 173884 356480 173904
rect 356480 173884 356482 173904
rect 356426 173848 356482 173884
rect 356518 173712 356574 173768
rect 356426 135244 356482 135280
rect 356426 135224 356428 135244
rect 356428 135224 356480 135244
rect 356480 135224 356482 135244
rect 356610 135224 356666 135280
rect 356150 3304 356206 3360
rect 357622 325624 357678 325680
rect 357806 325624 357862 325680
rect 357714 298288 357770 298344
rect 357622 298152 357678 298208
rect 357622 296656 357678 296712
rect 357806 296656 357862 296712
rect 357714 115912 357770 115968
rect 357806 115776 357862 115832
rect 357622 106256 357678 106312
rect 357806 106256 357862 106312
rect 357622 77288 357678 77344
rect 357806 77288 357862 77344
rect 359002 270680 359058 270736
rect 358910 270408 358966 270464
rect 358910 200096 358966 200152
rect 359094 200096 359150 200152
rect 358910 190440 358966 190496
rect 359186 190440 359242 190496
rect 364246 251232 364302 251288
rect 364246 251096 364302 251152
rect 364246 40432 364302 40488
rect 364246 40160 364302 40216
rect 365810 337456 365866 337512
rect 365810 315968 365866 316024
rect 365994 315968 366050 316024
rect 364430 217912 364486 217968
rect 364614 217912 364670 217968
rect 364430 200096 364486 200152
rect 364614 200096 364670 200152
rect 364614 190440 364670 190496
rect 364798 190440 364854 190496
rect 364522 172488 364578 172544
rect 364706 172488 364762 172544
rect 364522 135224 364578 135280
rect 364706 135224 364762 135280
rect 367006 170176 367062 170232
rect 367006 169768 367062 169824
rect 369766 182144 369822 182200
rect 369950 278704 370006 278760
rect 370318 278704 370374 278760
rect 370042 201456 370098 201512
rect 370226 201456 370282 201512
rect 369950 182164 370006 182200
rect 369950 182144 369952 182164
rect 369952 182144 370004 182164
rect 370004 182144 370006 182164
rect 370226 172488 370282 172544
rect 370410 172488 370466 172544
rect 370042 164192 370098 164248
rect 370226 164192 370282 164248
rect 370042 157528 370098 157584
rect 371882 170040 371938 170096
rect 371882 169768 371938 169824
rect 370042 154556 370098 154592
rect 370042 154536 370044 154556
rect 370044 154536 370096 154556
rect 370096 154536 370098 154556
rect 370134 138216 370190 138272
rect 370042 135244 370098 135280
rect 370042 135224 370044 135244
rect 370044 135224 370096 135244
rect 370096 135224 370098 135244
rect 370042 96600 370098 96656
rect 370226 96600 370282 96656
rect 370502 16768 370558 16824
rect 370502 16360 370558 16416
rect 373906 40568 373962 40624
rect 373906 40160 373962 40216
rect 375194 154536 375250 154592
rect 375562 251096 375618 251152
rect 375746 251096 375802 251152
rect 375562 231820 375564 231840
rect 375564 231820 375616 231840
rect 375616 231820 375618 231840
rect 375562 231784 375618 231820
rect 375838 231820 375840 231840
rect 375840 231820 375892 231840
rect 375892 231820 375894 231840
rect 375838 231784 375894 231820
rect 375562 212508 375564 212528
rect 375564 212508 375616 212528
rect 375616 212508 375618 212528
rect 375562 212472 375618 212508
rect 375838 212508 375840 212528
rect 375840 212508 375892 212528
rect 375892 212508 375894 212528
rect 375838 212472 375894 212508
rect 375562 191936 375618 191992
rect 375562 191820 375618 191856
rect 375562 191800 375564 191820
rect 375564 191800 375616 191820
rect 375616 191800 375618 191820
rect 375470 182144 375526 182200
rect 375746 182144 375802 182200
rect 375562 172488 375618 172544
rect 375746 172488 375802 172544
rect 375562 154556 375618 154592
rect 375562 154536 375564 154556
rect 375564 154536 375616 154556
rect 375616 154536 375618 154556
rect 375746 135360 375802 135416
rect 375562 135244 375618 135280
rect 375562 135224 375564 135244
rect 375564 135224 375616 135244
rect 375616 135224 375618 135244
rect 375746 96736 375802 96792
rect 375562 96600 375618 96656
rect 376758 241440 376814 241496
rect 376942 241440 376998 241496
rect 376758 222128 376814 222184
rect 376942 222128 376998 222184
rect 376758 202816 376814 202872
rect 376942 202816 376998 202872
rect 376758 183504 376814 183560
rect 376942 183504 376998 183560
rect 376758 154536 376814 154592
rect 376942 154536 376998 154592
rect 376758 135224 376814 135280
rect 376942 135224 376998 135280
rect 378506 337456 378562 337512
rect 380806 183504 380862 183560
rect 381174 260752 381230 260808
rect 381358 260752 381414 260808
rect 381082 183504 381138 183560
rect 381450 134544 381506 134600
rect 381450 134000 381506 134056
rect 381266 116048 381322 116104
rect 381082 115932 381138 115968
rect 381082 115912 381084 115932
rect 381084 115912 381136 115932
rect 381136 115912 381138 115932
rect 386326 170312 386382 170368
rect 386326 169904 386382 169960
rect 386786 270544 386842 270600
rect 386694 270408 386750 270464
rect 386602 212472 386658 212528
rect 386786 212472 386842 212528
rect 386602 193160 386658 193216
rect 386786 193160 386842 193216
rect 386602 135224 386658 135280
rect 386786 135224 386842 135280
rect 386602 115932 386658 115968
rect 386602 115912 386604 115932
rect 386604 115912 386656 115932
rect 386656 115912 386658 115932
rect 386786 115932 386842 115968
rect 386786 115912 386788 115932
rect 386788 115912 386840 115932
rect 386840 115912 386842 115932
rect 386602 96600 386658 96656
rect 386786 96600 386842 96656
rect 387982 66272 388038 66328
rect 388166 66272 388222 66328
rect 386510 16768 386566 16824
rect 386510 16496 386566 16552
rect 392122 249736 392178 249792
rect 392398 249736 392454 249792
rect 393226 231820 393228 231840
rect 393228 231820 393280 231840
rect 393280 231820 393282 231840
rect 393226 231784 393282 231820
rect 393410 231784 393466 231840
rect 392122 212472 392178 212528
rect 392306 212472 392362 212528
rect 393226 212508 393228 212528
rect 393228 212508 393280 212528
rect 393280 212508 393282 212528
rect 393226 212472 393282 212508
rect 393410 212472 393466 212528
rect 393226 193196 393228 193216
rect 393228 193196 393280 193216
rect 393280 193196 393282 193216
rect 393226 193160 393282 193196
rect 393410 193160 393466 193216
rect 392030 190440 392086 190496
rect 392214 190440 392270 190496
rect 393226 144900 393282 144936
rect 393226 144880 393228 144900
rect 393228 144880 393280 144900
rect 393280 144880 393282 144900
rect 393410 144880 393466 144936
rect 392122 115932 392178 115968
rect 392122 115912 392124 115932
rect 392124 115912 392176 115932
rect 392176 115912 392178 115932
rect 392306 115932 392362 115968
rect 392306 115912 392308 115932
rect 392308 115912 392360 115932
rect 392360 115912 392362 115932
rect 392122 96600 392178 96656
rect 392306 96600 392362 96656
rect 393226 96600 393282 96656
rect 393410 96600 393466 96656
rect 393410 67768 393466 67824
rect 393226 67632 393282 67688
rect 395986 134136 396042 134192
rect 395986 133728 396042 133784
rect 397366 279928 397422 279984
rect 397366 259392 397422 259448
rect 397366 212472 397422 212528
rect 397366 172488 397422 172544
rect 397734 280064 397790 280120
rect 397918 259392 397974 259448
rect 397550 212508 397552 212528
rect 397552 212508 397604 212528
rect 397604 212508 397606 212528
rect 397550 212472 397606 212508
rect 397550 193196 397552 193216
rect 397552 193196 397604 193216
rect 397604 193196 397606 193216
rect 397550 193160 397606 193196
rect 397734 193160 397790 193216
rect 397550 172488 397606 172544
rect 397642 40332 397644 40352
rect 397644 40332 397696 40352
rect 397696 40332 397698 40352
rect 397642 40296 397698 40332
rect 398930 16768 398986 16824
rect 398930 16496 398986 16552
rect 400310 241440 400366 241496
rect 400494 241440 400550 241496
rect 400310 222128 400366 222184
rect 400494 222128 400550 222184
rect 400310 202816 400366 202872
rect 400494 202816 400550 202872
rect 400310 154672 400366 154728
rect 400494 154536 400550 154592
rect 400310 106256 400366 106312
rect 400494 106256 400550 106312
rect 400310 96600 400366 96656
rect 400586 96600 400642 96656
rect 405646 40332 405648 40352
rect 405648 40332 405700 40352
rect 405700 40332 405702 40352
rect 405646 40296 405702 40332
rect 408406 16804 408408 16824
rect 408408 16804 408460 16824
rect 408460 16804 408462 16824
rect 408406 16768 408462 16804
rect 408774 259392 408830 259448
rect 408958 259392 409014 259448
rect 408682 193160 408738 193216
rect 408958 193160 409014 193216
rect 408406 3848 408462 3904
rect 408590 3884 408592 3904
rect 408592 3884 408644 3904
rect 408644 3884 408646 3904
rect 408590 3848 408646 3884
rect 408314 3612 408316 3632
rect 408316 3612 408368 3632
rect 408368 3612 408370 3632
rect 408314 3576 408370 3612
rect 408590 3612 408592 3632
rect 408592 3612 408644 3632
rect 408644 3612 408646 3632
rect 408590 3576 408646 3612
rect 410706 17040 410762 17096
rect 410614 3304 410670 3360
rect 415306 134272 415362 134328
rect 415306 134136 415362 134192
rect 416870 241440 416926 241496
rect 417146 241440 417202 241496
rect 416870 222128 416926 222184
rect 417146 222128 417202 222184
rect 416870 202816 416926 202872
rect 417146 202816 417202 202872
rect 416870 183504 416926 183560
rect 417146 183504 417202 183560
rect 416962 154536 417018 154592
rect 417146 154536 417202 154592
rect 416778 135224 416834 135280
rect 416962 135224 417018 135280
rect 416778 115912 416834 115968
rect 416962 115912 417018 115968
rect 416778 96600 416834 96656
rect 416962 96600 417018 96656
rect 418066 169904 418122 169960
rect 418066 169496 418122 169552
rect 418066 40296 418122 40352
rect 418158 40160 418214 40216
rect 418066 17040 418122 17096
rect 418250 16904 418306 16960
rect 422114 27512 422170 27568
rect 422390 183504 422446 183560
rect 422666 183504 422722 183560
rect 422298 27512 422354 27568
rect 425058 169804 425060 169824
rect 425060 169804 425112 169824
rect 425112 169804 425114 169824
rect 425058 169768 425114 169804
rect 428370 328616 428426 328672
rect 428002 328480 428058 328536
rect 427542 134136 427598 134192
rect 427726 134136 427782 134192
rect 427910 24792 427966 24848
rect 428094 24792 428150 24848
rect 433246 154536 433302 154592
rect 433430 241440 433486 241496
rect 433614 241440 433670 241496
rect 433430 222128 433486 222184
rect 433614 222128 433670 222184
rect 433430 202816 433486 202872
rect 433614 202816 433670 202872
rect 434534 170040 434590 170096
rect 433706 154536 433762 154592
rect 433614 135224 433670 135280
rect 433798 135224 433854 135280
rect 433430 96600 433486 96656
rect 433706 96600 433762 96656
rect 451554 325624 451610 325680
rect 451738 325624 451794 325680
rect 451278 288360 451334 288416
rect 451462 288360 451518 288416
rect 451278 231784 451334 231840
rect 451462 231784 451518 231840
rect 451278 212472 451334 212528
rect 451462 212472 451518 212528
rect 456798 40296 456854 40352
rect 456706 40160 456762 40216
rect 456798 16904 456854 16960
rect 456706 16768 456762 16824
rect 458822 134000 458878 134056
rect 458822 133728 458878 133784
rect 466458 96600 466514 96656
rect 466642 96600 466698 96656
rect 472070 241440 472126 241496
rect 472346 241440 472402 241496
rect 472070 222128 472126 222184
rect 472346 222128 472402 222184
rect 472070 202816 472126 202872
rect 472346 202816 472402 202872
rect 472070 183504 472126 183560
rect 472346 183504 472402 183560
rect 472162 154536 472218 154592
rect 472346 154536 472402 154592
rect 471978 115912 472034 115968
rect 472162 115912 472218 115968
rect 471978 96600 472034 96656
rect 472162 96600 472218 96656
rect 475934 169924 475990 169960
rect 475934 169904 475936 169924
rect 475936 169904 475988 169924
rect 475988 169904 475990 169924
rect 475934 40196 475936 40216
rect 475936 40196 475988 40216
rect 475988 40196 475990 40216
rect 475934 40160 475990 40196
rect 475934 16804 475936 16824
rect 475936 16804 475988 16824
rect 475988 16804 475990 16824
rect 475934 16768 475990 16804
rect 477498 16804 477500 16824
rect 477500 16804 477552 16824
rect 477552 16804 477554 16824
rect 477498 16768 477554 16804
rect 478142 169924 478198 169960
rect 478142 169904 478144 169924
rect 478144 169904 478196 169924
rect 478196 169904 478198 169924
rect 478234 40196 478236 40216
rect 478236 40196 478288 40216
rect 478288 40196 478290 40216
rect 478234 40160 478290 40196
rect 514574 134036 514576 134056
rect 514576 134036 514628 134056
rect 514628 134036 514630 134056
rect 514574 134000 514630 134036
rect 514574 40196 514576 40216
rect 514576 40196 514628 40216
rect 514628 40196 514630 40216
rect 514574 40160 514630 40196
rect 514574 16768 514630 16824
rect 514574 16360 514630 16416
rect 514850 134036 514852 134056
rect 514852 134036 514904 134056
rect 514904 134036 514906 134056
rect 514850 134000 514906 134036
rect 514850 40196 514852 40216
rect 514852 40196 514904 40216
rect 514904 40196 514906 40216
rect 514850 40160 514906 40196
rect 521658 170312 521714 170368
rect 521658 169768 521714 169824
rect 521658 22208 521714 22264
rect 521658 21936 521714 21992
rect 521658 16668 521660 16688
rect 521660 16668 521712 16688
rect 521712 16668 521714 16688
rect 521658 16632 521714 16668
rect 524510 16904 524566 16960
rect 528190 337320 528246 337376
rect 527454 336504 527510 336560
rect 527454 318960 527510 319016
rect 527638 309032 527694 309088
rect 527638 302096 527694 302152
rect 527638 289720 527694 289776
rect 527638 280336 527694 280392
rect 527454 270408 527510 270464
rect 527454 261024 527510 261080
rect 527454 251096 527510 251152
rect 527454 241712 527510 241768
rect 527638 231784 527694 231840
rect 527638 222264 527694 222320
rect 527454 212472 527510 212528
rect 527454 203088 527510 203144
rect 527454 193160 527510 193216
rect 527454 183776 527510 183832
rect 527270 173848 527326 173904
rect 527270 164192 527326 164248
rect 527270 154264 527326 154320
rect 527270 144880 527326 144936
rect 527822 135088 527878 135144
rect 527822 125568 527878 125624
rect 527454 96464 527510 96520
rect 527454 86944 527510 87000
rect 527270 57704 527326 57760
rect 527270 48320 527326 48376
rect 527454 38528 527510 38584
rect 527454 29144 527510 29200
rect 525706 3304 525762 3360
rect 529662 638288 529718 638344
rect 530306 638560 530362 638616
rect 531226 638424 531282 638480
rect 540886 170176 540942 170232
rect 540886 169904 540942 169960
rect 540978 133900 540980 133920
rect 540980 133900 541032 133920
rect 541032 133900 541034 133920
rect 540978 133864 541034 133900
rect 540978 40060 540980 40080
rect 540980 40060 541032 40080
rect 541032 40060 541034 40080
rect 540978 40024 541034 40060
rect 540886 17176 540942 17232
rect 540886 16768 540942 16824
rect 545854 134000 545910 134056
rect 545854 40160 545910 40216
rect 554502 134136 554558 134192
rect 554502 133728 554558 133784
rect 554502 40296 554558 40352
rect 554502 39888 554558 39944
rect 560206 170448 560262 170504
rect 560206 170040 560262 170096
rect 560206 17312 560262 17368
rect 560206 16904 560262 16960
rect 565082 337320 565138 337376
rect 580170 651072 580226 651128
rect 579802 642232 579858 642288
rect 579618 639784 579674 639840
rect 579618 639104 579674 639160
rect 579802 627680 579858 627736
rect 579802 604152 579858 604208
rect 579802 592456 579858 592512
rect 579802 557232 579858 557288
rect 579802 545536 579858 545592
rect 579802 533840 579858 533896
rect 579802 510312 579858 510368
rect 579802 498616 579858 498672
rect 579802 486784 579858 486840
rect 579802 463392 579858 463448
rect 579894 451696 579950 451752
rect 579894 439864 579950 439920
rect 579894 416472 579950 416528
rect 579894 404776 579950 404832
rect 579894 392944 579950 393000
rect 579986 369552 580042 369608
rect 580170 639376 580226 639432
rect 580078 357856 580134 357912
rect 579802 346024 579858 346080
rect 580078 322632 580134 322688
rect 580446 639240 580502 639296
rect 580262 639104 580318 639160
rect 580170 310800 580226 310856
rect 580170 263880 580226 263936
rect 579618 252184 579674 252240
rect 579618 216960 579674 217016
rect 580170 205264 580226 205320
rect 572626 169904 572682 169960
rect 572718 169768 572774 169824
rect 579710 158344 579766 158400
rect 572626 134000 572682 134056
rect 572718 133864 572774 133920
rect 580170 111424 580226 111480
rect 580170 64504 580226 64560
rect 572626 40160 572682 40216
rect 572718 40024 572774 40080
rect 580354 87896 580410 87952
rect 580906 299104 580962 299160
rect 580814 275712 580870 275768
rect 580722 228792 580778 228848
rect 580630 181872 580686 181928
rect 580538 123120 580594 123176
rect 580446 76200 580502 76256
rect 580262 29280 580318 29336
rect 572626 16768 572682 16824
rect 572718 16632 572774 16688
rect 575018 3304 575074 3360
<< metal3 >>
rect 8109 700362 8175 700365
rect 414013 700362 414079 700365
rect 8109 700360 414079 700362
rect 8109 700304 8114 700360
rect 8170 700304 414018 700360
rect 414074 700304 414079 700360
rect 8109 700302 414079 700304
rect 8109 700299 8175 700302
rect 414013 700299 414079 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 3509 643106 3575 643109
rect 520457 643106 520523 643109
rect 3509 643104 520523 643106
rect 3509 643048 3514 643104
rect 3570 643048 520462 643104
rect 520518 643048 520523 643104
rect 3509 643046 520523 643048
rect 3509 643043 3575 643046
rect 520457 643043 520523 643046
rect 233734 642908 233740 642972
rect 233804 642970 233810 642972
rect 259913 642970 259979 642973
rect 233804 642968 259979 642970
rect 233804 642912 259918 642968
rect 259974 642912 259979 642968
rect 233804 642910 259979 642912
rect 233804 642908 233810 642910
rect 259913 642907 259979 642910
rect 325693 642970 325759 642973
rect 526110 642970 526116 642972
rect 325693 642968 526116 642970
rect 325693 642912 325698 642968
rect 325754 642912 526116 642968
rect 325693 642910 526116 642912
rect 325693 642907 325759 642910
rect 526110 642908 526116 642910
rect 526180 642908 526186 642972
rect 258717 642834 258783 642837
rect 504633 642834 504699 642837
rect 258717 642832 504699 642834
rect 258717 642776 258722 642832
rect 258778 642776 504638 642832
rect 504694 642776 504699 642832
rect 258717 642774 504699 642776
rect 258717 642771 258783 642774
rect 504633 642771 504699 642774
rect 232814 642636 232820 642700
rect 232884 642698 232890 642700
rect 483657 642698 483723 642701
rect 232884 642696 483723 642698
rect 232884 642640 483662 642696
rect 483718 642640 483723 642696
rect 232884 642638 483723 642640
rect 232884 642636 232890 642638
rect 483657 642635 483723 642638
rect 232630 642500 232636 642564
rect 232700 642562 232706 642564
rect 491477 642562 491543 642565
rect 232700 642560 491543 642562
rect 232700 642504 491482 642560
rect 491538 642504 491543 642560
rect 232700 642502 491543 642504
rect 232700 642500 232706 642502
rect 491477 642499 491543 642502
rect 232446 642364 232452 642428
rect 232516 642426 232522 642428
rect 499389 642426 499455 642429
rect 232516 642424 499455 642426
rect 232516 642368 499394 642424
rect 499450 642368 499455 642424
rect 232516 642366 499455 642368
rect 232516 642364 232522 642366
rect 499389 642363 499455 642366
rect 241513 642290 241579 642293
rect 579797 642290 579863 642293
rect 241513 642288 579863 642290
rect 241513 642232 241518 642288
rect 241574 642232 579802 642288
rect 579858 642232 579863 642288
rect 241513 642230 579863 642232
rect 241513 642227 241579 642230
rect 579797 642227 579863 642230
rect 72417 642154 72483 642157
rect 429009 642154 429075 642157
rect 72417 642152 429075 642154
rect 72417 642096 72422 642152
rect 72478 642096 429014 642152
rect 429070 642096 429075 642152
rect 72417 642094 429075 642096
rect 72417 642091 72483 642094
rect 429009 642091 429075 642094
rect 434478 642092 434484 642156
rect 434548 642154 434554 642156
rect 507301 642154 507367 642157
rect 434548 642152 507367 642154
rect 434548 642096 507306 642152
rect 507362 642096 507367 642152
rect 434548 642094 507367 642096
rect 434548 642092 434554 642094
rect 507301 642091 507367 642094
rect 4889 642018 4955 642021
rect 494145 642018 494211 642021
rect 4889 642016 494211 642018
rect 4889 641960 4894 642016
rect 4950 641960 494150 642016
rect 494206 641960 494211 642016
rect 4889 641958 494211 641960
rect 4889 641955 4955 641958
rect 494145 641955 494211 641958
rect 3693 641882 3759 641885
rect 509969 641882 510035 641885
rect 3693 641880 510035 641882
rect 3693 641824 3698 641880
rect 3754 641824 509974 641880
rect 510030 641824 510035 641880
rect 3693 641822 510035 641824
rect 3693 641819 3759 641822
rect 509969 641819 510035 641822
rect 515857 641746 515923 641749
rect 525701 641746 525767 641749
rect 515857 641744 525767 641746
rect 515857 641688 515862 641744
rect 515918 641688 525706 641744
rect 525762 641688 525767 641744
rect 515857 641686 525767 641688
rect 515857 641683 515923 641686
rect 525701 641683 525767 641686
rect 7414 641548 7420 641612
rect 7484 641610 7490 641612
rect 12934 641610 12940 641612
rect 7484 641550 12940 641610
rect 7484 641548 7490 641550
rect 12934 641548 12940 641550
rect 13004 641548 13010 641612
rect 27654 641548 27660 641612
rect 27724 641610 27730 641612
rect 41597 641610 41663 641613
rect 27724 641608 41663 641610
rect 27724 641552 41602 641608
rect 41658 641552 41663 641608
rect 27724 641550 41663 641552
rect 27724 641548 27730 641550
rect 41597 641547 41663 641550
rect 53097 641610 53163 641613
rect 60917 641610 60983 641613
rect 53097 641608 60983 641610
rect 53097 641552 53102 641608
rect 53158 641552 60922 641608
rect 60978 641552 60983 641608
rect 53097 641550 60983 641552
rect 53097 641547 53163 641550
rect 60917 641547 60983 641550
rect 68461 641610 68527 641613
rect 79726 641610 79732 641612
rect 68461 641608 79732 641610
rect 68461 641552 68466 641608
rect 68522 641552 79732 641608
rect 68461 641550 79732 641552
rect 68461 641547 68527 641550
rect 79726 641548 79732 641550
rect 79796 641548 79802 641612
rect 91737 641610 91803 641613
rect 99557 641610 99623 641613
rect 91737 641608 99623 641610
rect 91737 641552 91742 641608
rect 91798 641552 99562 641608
rect 99618 641552 99623 641608
rect 91737 641550 99623 641552
rect 91737 641547 91803 641550
rect 99557 641547 99623 641550
rect 109718 641548 109724 641612
rect 109788 641610 109794 641612
rect 118877 641610 118943 641613
rect 109788 641608 118943 641610
rect 109788 641552 118882 641608
rect 118938 641552 118943 641608
rect 109788 641550 118943 641552
rect 109788 641548 109794 641550
rect 118877 641547 118943 641550
rect 130377 641610 130443 641613
rect 137318 641610 137324 641612
rect 130377 641608 137324 641610
rect 130377 641552 130382 641608
rect 130438 641552 137324 641608
rect 130377 641550 137324 641552
rect 130377 641547 130443 641550
rect 137318 641548 137324 641550
rect 137388 641548 137394 641612
rect 146109 641610 146175 641613
rect 157517 641610 157583 641613
rect 146109 641608 157583 641610
rect 146109 641552 146114 641608
rect 146170 641552 157522 641608
rect 157578 641552 157583 641608
rect 146109 641550 157583 641552
rect 146109 641547 146175 641550
rect 157517 641547 157583 641550
rect 167310 641548 167316 641612
rect 167380 641610 167386 641612
rect 176837 641610 176903 641613
rect 167380 641608 176903 641610
rect 167380 641552 176842 641608
rect 176898 641552 176903 641608
rect 167380 641550 176903 641552
rect 167380 641548 167386 641550
rect 176837 641547 176903 641550
rect 188337 641610 188403 641613
rect 193949 641610 194015 641613
rect 188337 641608 194015 641610
rect 188337 641552 188342 641608
rect 188398 641552 193954 641608
rect 194010 641552 194015 641608
rect 188337 641550 194015 641552
rect 188337 641547 188403 641550
rect 193949 641547 194015 641550
rect 207657 641610 207723 641613
rect 215150 641610 215156 641612
rect 207657 641608 215156 641610
rect 207657 641552 207662 641608
rect 207718 641552 215156 641608
rect 207657 641550 215156 641552
rect 207657 641547 207723 641550
rect 215150 641548 215156 641550
rect 215220 641548 215226 641612
rect 222142 641548 222148 641612
rect 222212 641610 222218 641612
rect 226006 641610 226012 641612
rect 222212 641550 226012 641610
rect 222212 641548 222218 641550
rect 226006 641548 226012 641550
rect 226076 641548 226082 641612
rect 231894 641548 231900 641612
rect 231964 641610 231970 641612
rect 243537 641610 243603 641613
rect 231964 641608 243603 641610
rect 231964 641552 243542 641608
rect 243598 641552 243603 641608
rect 231964 641550 243603 641552
rect 231964 641548 231970 641550
rect 243537 641547 243603 641550
rect 275277 641610 275343 641613
rect 282678 641610 282684 641612
rect 275277 641608 282684 641610
rect 275277 641552 275282 641608
rect 275338 641552 282684 641608
rect 275277 641550 282684 641552
rect 275277 641547 275343 641550
rect 282678 641548 282684 641550
rect 282748 641548 282754 641612
rect 301630 641548 301636 641612
rect 301700 641610 301706 641612
rect 302918 641610 302924 641612
rect 301700 641550 302924 641610
rect 301700 641548 301706 641550
rect 302918 641548 302924 641550
rect 302988 641548 302994 641612
rect 309358 641548 309364 641612
rect 309428 641610 309434 641612
rect 318374 641610 318380 641612
rect 309428 641550 318380 641610
rect 309428 641548 309434 641550
rect 318374 641548 318380 641550
rect 318444 641548 318450 641612
rect 327022 641548 327028 641612
rect 327092 641610 327098 641612
rect 336590 641610 336596 641612
rect 327092 641550 336596 641610
rect 327092 641548 327098 641550
rect 336590 641548 336596 641550
rect 336660 641548 336666 641612
rect 348366 641548 348372 641612
rect 348436 641610 348442 641612
rect 351126 641610 351132 641612
rect 348436 641550 351132 641610
rect 348436 641548 348442 641550
rect 351126 641548 351132 641550
rect 351196 641548 351202 641612
rect 376702 641548 376708 641612
rect 376772 641610 376778 641612
rect 379646 641610 379652 641612
rect 376772 641550 379652 641610
rect 376772 641548 376778 641550
rect 379646 641548 379652 641550
rect 379716 641548 379722 641612
rect 423622 641548 423628 641612
rect 423692 641610 423698 641612
rect 432454 641610 432460 641612
rect 423692 641550 432460 641610
rect 423692 641548 423698 641550
rect 432454 641548 432460 641550
rect 432524 641548 432530 641612
rect 453982 641548 453988 641612
rect 454052 641610 454058 641612
rect 463550 641610 463556 641612
rect 454052 641550 463556 641610
rect 454052 641548 454058 641550
rect 463550 641548 463556 641550
rect 463620 641548 463626 641612
rect 41597 640930 41663 640933
rect 53097 640930 53163 640933
rect 41597 640928 53163 640930
rect 41597 640872 41602 640928
rect 41658 640872 53102 640928
rect 53158 640872 53163 640928
rect 41597 640870 53163 640872
rect 41597 640867 41663 640870
rect 53097 640867 53163 640870
rect 60917 640930 60983 640933
rect 68461 640930 68527 640933
rect 60917 640928 68527 640930
rect 60917 640872 60922 640928
rect 60978 640872 68466 640928
rect 68522 640872 68527 640928
rect 60917 640870 68527 640872
rect 60917 640867 60983 640870
rect 68461 640867 68527 640870
rect 80830 640868 80836 640932
rect 80900 640930 80906 640932
rect 91737 640930 91803 640933
rect 80900 640928 91803 640930
rect 80900 640872 91742 640928
rect 91798 640872 91803 640928
rect 80900 640870 91803 640872
rect 80900 640868 80906 640870
rect 91737 640867 91803 640870
rect 99557 640930 99623 640933
rect 108430 640930 108436 640932
rect 99557 640928 108436 640930
rect 99557 640872 99562 640928
rect 99618 640872 108436 640928
rect 99557 640870 108436 640872
rect 99557 640867 99623 640870
rect 108430 640868 108436 640870
rect 108500 640868 108506 640932
rect 118877 640930 118943 640933
rect 130377 640930 130443 640933
rect 118877 640928 130443 640930
rect 118877 640872 118882 640928
rect 118938 640872 130382 640928
rect 130438 640872 130443 640928
rect 118877 640870 130443 640872
rect 118877 640867 118943 640870
rect 130377 640867 130443 640870
rect 138422 640868 138428 640932
rect 138492 640930 138498 640932
rect 146109 640930 146175 640933
rect 138492 640928 146175 640930
rect 138492 640872 146114 640928
rect 146170 640872 146175 640928
rect 138492 640870 146175 640872
rect 138492 640868 138498 640870
rect 146109 640867 146175 640870
rect 157517 640930 157583 640933
rect 166022 640930 166028 640932
rect 157517 640928 166028 640930
rect 157517 640872 157522 640928
rect 157578 640872 166028 640928
rect 157517 640870 166028 640872
rect 157517 640867 157583 640870
rect 166022 640868 166028 640870
rect 166092 640868 166098 640932
rect 176837 640930 176903 640933
rect 188337 640930 188403 640933
rect 176837 640928 188403 640930
rect 176837 640872 176842 640928
rect 176898 640872 188342 640928
rect 188398 640872 188403 640928
rect 176837 640870 188403 640872
rect 176837 640867 176903 640870
rect 188337 640867 188403 640870
rect 193949 640930 194015 640933
rect 207657 640930 207723 640933
rect 193949 640928 207723 640930
rect 193949 640872 193954 640928
rect 194010 640872 207662 640928
rect 207718 640872 207723 640928
rect 193949 640870 207723 640872
rect 193949 640867 194015 640870
rect 207657 640867 207723 640870
rect 243537 640930 243603 640933
rect 251766 640930 251772 640932
rect 243537 640928 251772 640930
rect 243537 640872 243542 640928
rect 243598 640872 251772 640928
rect 243537 640870 251772 640872
rect 243537 640867 243603 640870
rect 251766 640868 251772 640870
rect 251836 640868 251842 640932
rect 264462 640868 264468 640932
rect 264532 640930 264538 640932
rect 275277 640930 275343 640933
rect 264532 640928 275343 640930
rect 264532 640872 275282 640928
rect 275338 640872 275343 640928
rect 264532 640870 275343 640872
rect 264532 640868 264538 640870
rect 275277 640867 275343 640870
rect 289854 640868 289860 640932
rect 289924 640930 289930 640932
rect 299238 640930 299244 640932
rect 289924 640870 299244 640930
rect 289924 640868 289930 640870
rect 299238 640868 299244 640870
rect 299308 640868 299314 640932
rect 318742 640868 318748 640932
rect 318812 640930 318818 640932
rect 322054 640930 322060 640932
rect 318812 640870 322060 640930
rect 318812 640868 318818 640870
rect 322054 640868 322060 640870
rect 322124 640868 322130 640932
rect 357382 640868 357388 640932
rect 357452 640930 357458 640932
rect 366950 640930 366956 640932
rect 357452 640870 366956 640930
rect 357452 640868 357458 640870
rect 366950 640868 366956 640870
rect 367020 640868 367026 640932
rect 367134 640868 367140 640932
rect 367204 640930 367210 640932
rect 376518 640930 376524 640932
rect 367204 640870 376524 640930
rect 367204 640868 367210 640870
rect 376518 640868 376524 640870
rect 376588 640868 376594 640932
rect 389030 640868 389036 640932
rect 389100 640930 389106 640932
rect 395654 640930 395660 640932
rect 389100 640870 395660 640930
rect 389100 640868 389106 640870
rect 395654 640868 395660 640870
rect 395724 640868 395730 640932
rect 396022 640868 396028 640932
rect 396092 640930 396098 640932
rect 399334 640930 399340 640932
rect 396092 640870 399340 640930
rect 396092 640868 396098 640870
rect 399334 640868 399340 640870
rect 399404 640868 399410 640932
rect 436134 640868 436140 640932
rect 436204 640930 436210 640932
rect 438526 640930 438532 640932
rect 436204 640870 438532 640930
rect 436204 640868 436210 640870
rect 438526 640868 438532 640870
rect 438596 640868 438602 640932
rect 463918 640188 463924 640252
rect 463988 640250 463994 640252
rect 480846 640250 480852 640252
rect 463988 640190 480852 640250
rect 463988 640188 463994 640190
rect 480846 640188 480852 640190
rect 480916 640188 480922 640252
rect 509182 640188 509188 640252
rect 509252 640250 509258 640252
rect 515857 640250 515923 640253
rect 509252 640248 515923 640250
rect 509252 640192 515862 640248
rect 515918 640192 515923 640248
rect 509252 640190 515923 640192
rect 509252 640188 509258 640190
rect 515857 640187 515923 640190
rect 244181 640114 244247 640117
rect 302049 640116 302115 640117
rect 252134 640114 252140 640116
rect 244181 640112 252140 640114
rect 244181 640056 244186 640112
rect 244242 640056 252140 640112
rect 244181 640054 252140 640056
rect 244181 640051 244247 640054
rect 252134 640052 252140 640054
rect 252204 640052 252210 640116
rect 301998 640114 302004 640116
rect 301958 640054 302004 640114
rect 302068 640112 302115 640116
rect 302110 640056 302115 640112
rect 301998 640052 302004 640054
rect 302068 640052 302115 640056
rect 326286 640052 326292 640116
rect 326356 640114 326362 640116
rect 336406 640114 336412 640116
rect 326356 640054 336412 640114
rect 326356 640052 326362 640054
rect 336406 640052 336412 640054
rect 336476 640052 336482 640116
rect 345790 640114 345796 640116
rect 340646 640054 345796 640114
rect 302049 640051 302115 640052
rect 231393 639978 231459 639981
rect 328177 639980 328243 639981
rect 231710 639978 231716 639980
rect 231393 639976 231716 639978
rect 231393 639920 231398 639976
rect 231454 639920 231716 639976
rect 231393 639918 231716 639920
rect 231393 639915 231459 639918
rect 231710 639916 231716 639918
rect 231780 639916 231786 639980
rect 232998 639916 233004 639980
rect 233068 639978 233074 639980
rect 239438 639978 239444 639980
rect 233068 639918 239444 639978
rect 233068 639916 233074 639918
rect 239438 639916 239444 639918
rect 239508 639916 239514 639980
rect 251766 639916 251772 639980
rect 251836 639978 251842 639980
rect 257838 639978 257844 639980
rect 251836 639918 257844 639978
rect 251836 639916 251842 639918
rect 257838 639916 257844 639918
rect 257908 639916 257914 639980
rect 287094 639916 287100 639980
rect 287164 639978 287170 639980
rect 297398 639978 297404 639980
rect 287164 639918 297404 639978
rect 287164 639916 287170 639918
rect 297398 639916 297404 639918
rect 297468 639916 297474 639980
rect 306598 639916 306604 639980
rect 306668 639978 306674 639980
rect 316718 639978 316724 639980
rect 306668 639918 316724 639978
rect 306668 639916 306674 639918
rect 316718 639916 316724 639918
rect 316788 639916 316794 639980
rect 328126 639978 328132 639980
rect 328086 639918 328132 639978
rect 328196 639976 328243 639980
rect 328238 639920 328243 639976
rect 328126 639916 328132 639918
rect 328196 639916 328243 639920
rect 335302 639916 335308 639980
rect 335372 639978 335378 639980
rect 340646 639978 340706 640054
rect 345790 640052 345796 640054
rect 345860 640052 345866 640116
rect 403566 640052 403572 640116
rect 403636 640114 403642 640116
rect 413318 640114 413324 640116
rect 403636 640054 413324 640114
rect 403636 640052 403642 640054
rect 413318 640052 413324 640054
rect 413388 640052 413394 640116
rect 456742 640052 456748 640116
rect 456812 640114 456818 640116
rect 463417 640114 463483 640117
rect 456812 640112 463483 640114
rect 456812 640056 463422 640112
rect 463478 640056 463483 640112
rect 456812 640054 463483 640056
rect 456812 640052 456818 640054
rect 463417 640051 463483 640054
rect 335372 639918 340706 639978
rect 335372 639916 335378 639918
rect 345606 639916 345612 639980
rect 345676 639978 345682 639980
rect 372286 639978 372292 639980
rect 345676 639918 372292 639978
rect 345676 639916 345682 639918
rect 372286 639916 372292 639918
rect 372356 639916 372362 639980
rect 384246 639916 384252 639980
rect 384316 639978 384322 639980
rect 393078 639978 393084 639980
rect 384316 639918 393084 639978
rect 384316 639916 384322 639918
rect 393078 639916 393084 639918
rect 393148 639916 393154 639980
rect 441654 639916 441660 639980
rect 441724 639978 441730 639980
rect 451958 639978 451964 639980
rect 441724 639918 451964 639978
rect 441724 639916 441730 639918
rect 451958 639916 451964 639918
rect 452028 639916 452034 639980
rect 463233 639978 463299 639981
rect 471053 639978 471119 639981
rect 463233 639976 471119 639978
rect 463233 639920 463238 639976
rect 463294 639920 471058 639976
rect 471114 639920 471119 639976
rect 463233 639918 471119 639920
rect 328177 639915 328243 639916
rect 463233 639915 463299 639918
rect 471053 639915 471119 639918
rect 4153 639842 4219 639845
rect 5390 639842 5396 639844
rect 4153 639840 5396 639842
rect 4153 639784 4158 639840
rect 4214 639784 5396 639840
rect 4153 639782 5396 639784
rect 4153 639779 4219 639782
rect 5390 639780 5396 639782
rect 5460 639780 5466 639844
rect 109677 639842 109743 639845
rect 119337 639842 119403 639845
rect 109677 639840 119403 639842
rect 109677 639784 109682 639840
rect 109738 639784 119342 639840
rect 119398 639784 119403 639840
rect 109677 639782 119403 639784
rect 109677 639779 109743 639782
rect 119337 639779 119403 639782
rect 162853 639842 162919 639845
rect 177297 639842 177363 639845
rect 162853 639840 177363 639842
rect 162853 639784 162858 639840
rect 162914 639784 177302 639840
rect 177358 639784 177363 639840
rect 162853 639782 177363 639784
rect 162853 639779 162919 639782
rect 177297 639779 177363 639782
rect 233969 639842 234035 639845
rect 234470 639842 234476 639844
rect 233969 639840 234476 639842
rect 233969 639784 233974 639840
rect 234030 639784 234476 639840
rect 233969 639782 234476 639784
rect 233969 639779 234035 639782
rect 234470 639780 234476 639782
rect 234540 639780 234546 639844
rect 235257 639842 235323 639845
rect 235574 639842 235580 639844
rect 235257 639840 235580 639842
rect 235257 639784 235262 639840
rect 235318 639784 235580 639840
rect 235257 639782 235580 639784
rect 235257 639779 235323 639782
rect 235574 639780 235580 639782
rect 235644 639780 235650 639844
rect 249374 639780 249380 639844
rect 249444 639842 249450 639844
rect 249517 639842 249583 639845
rect 249444 639840 249583 639842
rect 249444 639784 249522 639840
rect 249578 639784 249583 639840
rect 249444 639782 249583 639784
rect 249444 639780 249450 639782
rect 249517 639779 249583 639782
rect 254945 639842 255011 639845
rect 255630 639842 255636 639844
rect 254945 639840 255636 639842
rect 254945 639784 254950 639840
rect 255006 639784 255636 639840
rect 254945 639782 255636 639784
rect 254945 639779 255011 639782
rect 255630 639780 255636 639782
rect 255700 639780 255706 639844
rect 267774 639780 267780 639844
rect 267844 639842 267850 639844
rect 282310 639842 282316 639844
rect 267844 639782 282316 639842
rect 267844 639780 267850 639782
rect 282310 639780 282316 639782
rect 282380 639780 282386 639844
rect 289997 639842 290063 639845
rect 340781 639842 340847 639845
rect 289997 639840 340847 639842
rect 289997 639784 290002 639840
rect 290058 639784 340786 639840
rect 340842 639784 340847 639840
rect 289997 639782 340847 639784
rect 289997 639779 290063 639782
rect 340781 639779 340847 639782
rect 340965 639842 341031 639845
rect 579613 639842 579679 639845
rect 340965 639840 579679 639842
rect 340965 639784 340970 639840
rect 341026 639784 579618 639840
rect 579674 639784 579679 639840
rect 340965 639782 579679 639784
rect 340965 639779 341031 639782
rect 579613 639779 579679 639782
rect 3877 639706 3943 639709
rect 340781 639706 340847 639709
rect 3877 639704 340847 639706
rect 3877 639648 3882 639704
rect 3938 639648 340786 639704
rect 340842 639648 340847 639704
rect 3877 639646 340847 639648
rect 3877 639643 3943 639646
rect 340781 639643 340847 639646
rect 340965 639706 341031 639709
rect 462957 639706 463023 639709
rect 463233 639706 463299 639709
rect 340965 639704 463023 639706
rect 340965 639648 340970 639704
rect 341026 639648 462962 639704
rect 463018 639648 463023 639704
rect 340965 639646 463023 639648
rect 340965 639643 341031 639646
rect 462957 639643 463023 639646
rect 463190 639704 463299 639706
rect 463190 639648 463238 639704
rect 463294 639648 463299 639704
rect 463190 639643 463299 639648
rect 463417 639706 463483 639709
rect 470133 639706 470199 639709
rect 463417 639704 470199 639706
rect 463417 639648 463422 639704
rect 463478 639648 470138 639704
rect 470194 639648 470199 639704
rect 463417 639646 470199 639648
rect 463417 639643 463483 639646
rect 470133 639643 470199 639646
rect 471053 639706 471119 639709
rect 485129 639706 485195 639709
rect 471053 639704 471162 639706
rect 471053 639648 471058 639704
rect 471114 639648 471162 639704
rect 471053 639643 471162 639648
rect 3417 639570 3483 639573
rect 5533 639570 5599 639573
rect 3417 639568 5599 639570
rect 3417 639512 3422 639568
rect 3478 639512 5538 639568
rect 5594 639512 5599 639568
rect 3417 639510 5599 639512
rect 3417 639507 3483 639510
rect 5533 639507 5599 639510
rect 23381 639570 23447 639573
rect 23381 639568 23490 639570
rect 23381 639512 23386 639568
rect 23442 639512 23490 639568
rect 23381 639507 23490 639512
rect 32990 639508 32996 639572
rect 33060 639570 33066 639572
rect 33174 639570 33180 639572
rect 33060 639510 33180 639570
rect 33060 639508 33066 639510
rect 33174 639508 33180 639510
rect 33244 639508 33250 639572
rect 147765 639570 147831 639573
rect 156321 639570 156387 639573
rect 147765 639568 156387 639570
rect 147765 639512 147770 639568
rect 147826 639512 156326 639568
rect 156382 639512 156387 639568
rect 147765 639510 156387 639512
rect 147765 639507 147831 639510
rect 156321 639507 156387 639510
rect 186313 639570 186379 639573
rect 220813 639570 220879 639573
rect 186313 639568 198106 639570
rect 186313 639512 186318 639568
rect 186374 639512 198106 639568
rect 186313 639510 198106 639512
rect 186313 639507 186379 639510
rect 23430 639298 23490 639507
rect 33174 639372 33180 639436
rect 33244 639434 33250 639436
rect 50797 639434 50863 639437
rect 33244 639432 50863 639434
rect 33244 639376 50802 639432
rect 50858 639376 50863 639432
rect 33244 639374 50863 639376
rect 33244 639372 33250 639374
rect 50797 639371 50863 639374
rect 51073 639434 51139 639437
rect 60641 639434 60707 639437
rect 70117 639434 70183 639437
rect 51073 639432 60707 639434
rect 51073 639376 51078 639432
rect 51134 639376 60646 639432
rect 60702 639376 60707 639432
rect 51073 639374 60707 639376
rect 51073 639371 51139 639374
rect 60641 639371 60707 639374
rect 66118 639432 70183 639434
rect 66118 639376 70122 639432
rect 70178 639376 70183 639432
rect 66118 639374 70183 639376
rect 66118 639301 66178 639374
rect 70117 639371 70183 639374
rect 70393 639434 70459 639437
rect 79961 639434 80027 639437
rect 70393 639432 80027 639434
rect 70393 639376 70398 639432
rect 70454 639376 79966 639432
rect 80022 639376 80027 639432
rect 70393 639374 80027 639376
rect 70393 639371 70459 639374
rect 79961 639371 80027 639374
rect 80145 639434 80211 639437
rect 89437 639434 89503 639437
rect 80145 639432 89503 639434
rect 80145 639376 80150 639432
rect 80206 639376 89442 639432
rect 89498 639376 89503 639432
rect 80145 639374 89503 639376
rect 80145 639371 80211 639374
rect 89437 639371 89503 639374
rect 89713 639434 89779 639437
rect 119337 639434 119403 639437
rect 147581 639434 147647 639437
rect 89713 639432 99298 639434
rect 89713 639376 89718 639432
rect 89774 639376 99298 639432
rect 89713 639374 99298 639376
rect 89713 639371 89779 639374
rect 32990 639298 32996 639300
rect -960 639012 480 639252
rect 23430 639238 32996 639298
rect 32990 639236 32996 639238
rect 33060 639236 33066 639300
rect 66118 639296 66227 639301
rect 66118 639240 66166 639296
rect 66222 639240 66227 639296
rect 66118 639238 66227 639240
rect 99238 639298 99298 639374
rect 119337 639432 147647 639434
rect 119337 639376 119342 639432
rect 119398 639376 147586 639432
rect 147642 639376 147647 639432
rect 119337 639374 147647 639376
rect 119337 639371 119403 639374
rect 147581 639371 147647 639374
rect 177297 639434 177363 639437
rect 186037 639434 186103 639437
rect 177297 639432 186103 639434
rect 177297 639376 177302 639432
rect 177358 639376 186042 639432
rect 186098 639376 186103 639432
rect 177297 639374 186103 639376
rect 198046 639434 198106 639510
rect 212398 639568 220879 639570
rect 212398 639512 220818 639568
rect 220874 639512 220879 639568
rect 212398 639510 220879 639512
rect 201493 639434 201559 639437
rect 198046 639432 201559 639434
rect 198046 639376 201498 639432
rect 201554 639376 201559 639432
rect 198046 639374 201559 639376
rect 177297 639371 177363 639374
rect 186037 639371 186103 639374
rect 201493 639371 201559 639374
rect 109677 639298 109743 639301
rect 99238 639296 109743 639298
rect 99238 639240 109682 639296
rect 109738 639240 109743 639296
rect 99238 639238 109743 639240
rect 66161 639235 66227 639238
rect 109677 639235 109743 639238
rect 211061 639298 211127 639301
rect 212398 639298 212458 639510
rect 220813 639507 220879 639510
rect 235574 639508 235580 639572
rect 235644 639570 235650 639572
rect 249006 639570 249012 639572
rect 235644 639510 249012 639570
rect 235644 639508 235650 639510
rect 249006 639508 249012 639510
rect 249076 639508 249082 639572
rect 463190 639570 463250 639643
rect 257662 639510 268026 639570
rect 239438 639372 239444 639436
rect 239508 639434 239514 639436
rect 251766 639434 251772 639436
rect 239508 639374 251772 639434
rect 239508 639372 239514 639374
rect 251766 639372 251772 639374
rect 251836 639372 251842 639436
rect 257662 639434 257722 639510
rect 251958 639374 257722 639434
rect 211061 639296 212458 639298
rect 211061 639240 211066 639296
rect 211122 639240 212458 639296
rect 211061 639238 212458 639240
rect 211061 639235 211127 639238
rect 249006 639236 249012 639300
rect 249076 639298 249082 639300
rect 251958 639298 252018 639374
rect 257838 639372 257844 639436
rect 257908 639434 257914 639436
rect 267774 639434 267780 639436
rect 257908 639374 267780 639434
rect 257908 639372 257914 639374
rect 267774 639372 267780 639374
rect 267844 639372 267850 639436
rect 267966 639434 268026 639510
rect 277166 639510 287346 639570
rect 277166 639434 277226 639510
rect 267966 639374 277226 639434
rect 282310 639372 282316 639436
rect 282380 639434 282386 639436
rect 287094 639434 287100 639436
rect 282380 639374 287100 639434
rect 282380 639372 282386 639374
rect 287094 639372 287100 639374
rect 287164 639372 287170 639436
rect 287286 639434 287346 639510
rect 297222 639510 307034 639570
rect 297222 639434 297282 639510
rect 287286 639374 297282 639434
rect 297398 639372 297404 639436
rect 297468 639434 297474 639436
rect 306598 639434 306604 639436
rect 297468 639374 306604 639434
rect 297468 639372 297474 639374
rect 306598 639372 306604 639374
rect 306668 639372 306674 639436
rect 306974 639434 307034 639510
rect 316542 639510 326538 639570
rect 316542 639434 316602 639510
rect 306974 639374 316602 639434
rect 316718 639372 316724 639436
rect 316788 639434 316794 639436
rect 326286 639434 326292 639436
rect 316788 639374 326292 639434
rect 316788 639372 316794 639374
rect 326286 639372 326292 639374
rect 326356 639372 326362 639436
rect 326478 639434 326538 639510
rect 371926 639510 384498 639570
rect 335302 639434 335308 639436
rect 326478 639374 335308 639434
rect 335302 639372 335308 639374
rect 335372 639372 335378 639436
rect 336406 639372 336412 639436
rect 336476 639434 336482 639436
rect 345606 639434 345612 639436
rect 336476 639374 345612 639434
rect 336476 639372 336482 639374
rect 345606 639372 345612 639374
rect 345676 639372 345682 639436
rect 345790 639372 345796 639436
rect 345860 639434 345866 639436
rect 371926 639434 371986 639510
rect 345860 639374 371986 639434
rect 345860 639372 345866 639374
rect 372286 639372 372292 639436
rect 372356 639434 372362 639436
rect 384246 639434 384252 639436
rect 372356 639374 384252 639434
rect 372356 639372 372362 639374
rect 384246 639372 384252 639374
rect 384316 639372 384322 639436
rect 384438 639434 384498 639510
rect 392902 639510 441906 639570
rect 392902 639434 392962 639510
rect 384438 639374 392962 639434
rect 393078 639372 393084 639436
rect 393148 639434 393154 639436
rect 403566 639434 403572 639436
rect 393148 639374 403572 639434
rect 393148 639372 393154 639374
rect 403566 639372 403572 639374
rect 403636 639372 403642 639436
rect 413318 639372 413324 639436
rect 413388 639434 413394 639436
rect 441654 639434 441660 639436
rect 413388 639374 441660 639434
rect 413388 639372 413394 639374
rect 441654 639372 441660 639374
rect 441724 639372 441730 639436
rect 441846 639434 441906 639510
rect 451782 639510 463250 639570
rect 471102 639570 471162 639643
rect 480670 639704 485195 639706
rect 480670 639648 485134 639704
rect 485190 639648 485195 639704
rect 480670 639646 485195 639648
rect 480670 639570 480730 639646
rect 485129 639643 485195 639646
rect 493358 639644 493364 639708
rect 493428 639706 493434 639708
rect 496629 639706 496695 639709
rect 493428 639704 496695 639706
rect 493428 639648 496634 639704
rect 496690 639648 496695 639704
rect 493428 639646 496695 639648
rect 493428 639644 493434 639646
rect 496629 639643 496695 639646
rect 509182 639644 509188 639708
rect 509252 639706 509258 639708
rect 512269 639706 512335 639709
rect 509252 639704 512335 639706
rect 509252 639648 512274 639704
rect 512330 639648 512335 639704
rect 509252 639646 512335 639648
rect 509252 639644 509258 639646
rect 512269 639643 512335 639646
rect 527398 639644 527404 639708
rect 527468 639706 527474 639708
rect 528093 639706 528159 639709
rect 527468 639704 528159 639706
rect 527468 639648 528098 639704
rect 528154 639648 528159 639704
rect 527468 639646 528159 639648
rect 527468 639644 527474 639646
rect 528093 639643 528159 639646
rect 471102 639510 480730 639570
rect 451782 639434 451842 639510
rect 441846 639374 451842 639434
rect 451958 639372 451964 639436
rect 452028 639434 452034 639436
rect 456742 639434 456748 639436
rect 452028 639374 456748 639434
rect 452028 639372 452034 639374
rect 456742 639372 456748 639374
rect 456812 639372 456818 639436
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 249076 639238 252018 639298
rect 249076 639236 249082 639238
rect 252134 639236 252140 639300
rect 252204 639298 252210 639300
rect 580441 639298 580507 639301
rect 252204 639296 580507 639298
rect 252204 639240 580446 639296
rect 580502 639240 580507 639296
rect 583520 639284 584960 639374
rect 252204 639238 580507 639240
rect 252204 639236 252210 639238
rect 580441 639235 580507 639238
rect 6177 639162 6243 639165
rect 493358 639162 493364 639164
rect 6177 639160 493364 639162
rect 6177 639104 6182 639160
rect 6238 639104 493364 639160
rect 6177 639102 493364 639104
rect 6177 639099 6243 639102
rect 493358 639100 493364 639102
rect 493428 639100 493434 639164
rect 579613 639162 579679 639165
rect 580257 639162 580323 639165
rect 579613 639160 580323 639162
rect 579613 639104 579618 639160
rect 579674 639104 580262 639160
rect 580318 639104 580323 639160
rect 579613 639102 580323 639104
rect 579613 639099 579679 639102
rect 580257 639099 580323 639102
rect 3601 639026 3667 639029
rect 509182 639026 509188 639028
rect 3601 639024 509188 639026
rect 3601 638968 3606 639024
rect 3662 638968 509188 639024
rect 3601 638966 509188 638968
rect 3601 638963 3667 638966
rect 509182 638964 509188 638966
rect 509252 638964 509258 639028
rect 328126 638556 328132 638620
rect 328196 638618 328202 638620
rect 530301 638618 530367 638621
rect 328196 638616 530367 638618
rect 328196 638560 530306 638616
rect 530362 638560 530367 638616
rect 328196 638558 530367 638560
rect 328196 638556 328202 638558
rect 530301 638555 530367 638558
rect 301998 638420 302004 638484
rect 302068 638482 302074 638484
rect 531221 638482 531287 638485
rect 302068 638480 531287 638482
rect 302068 638424 531226 638480
rect 531282 638424 531287 638480
rect 302068 638422 531287 638424
rect 302068 638420 302074 638422
rect 531221 638419 531287 638422
rect 255630 638284 255636 638348
rect 255700 638346 255706 638348
rect 529657 638346 529723 638349
rect 255700 638344 529723 638346
rect 255700 638288 529662 638344
rect 529718 638288 529723 638344
rect 255700 638286 529723 638288
rect 255700 638284 255706 638286
rect 529657 638283 529723 638286
rect 3785 638210 3851 638213
rect 434478 638210 434484 638212
rect 3785 638208 434484 638210
rect 3785 638152 3790 638208
rect 3846 638152 434484 638208
rect 3785 638150 434484 638152
rect 3785 638147 3851 638150
rect 434478 638148 434484 638150
rect 434548 638148 434554 638212
rect 526110 637740 526116 637804
rect 526180 637802 526186 637804
rect 527214 637802 527220 637804
rect 526180 637742 527220 637802
rect 526180 637740 526186 637742
rect 527214 637740 527220 637742
rect 527284 637740 527290 637804
rect 527214 634340 527220 634404
rect 527284 634402 527290 634404
rect 527582 634402 527588 634404
rect 527284 634342 527588 634402
rect 527284 634340 527290 634342
rect 527582 634340 527588 634342
rect 527652 634340 527658 634404
rect 527398 634266 527404 634268
rect 527222 634206 527404 634266
rect 527222 633996 527282 634206
rect 527398 634204 527404 634206
rect 527468 634204 527474 634268
rect 527214 633932 527220 633996
rect 527284 633932 527290 633996
rect 527582 630730 527588 630732
rect 527406 630670 527588 630730
rect 527406 630596 527466 630670
rect 527582 630668 527588 630670
rect 527652 630668 527658 630732
rect 527398 630532 527404 630596
rect 527468 630532 527474 630596
rect 527766 627812 527772 627876
rect 527836 627874 527842 627876
rect 528502 627874 528508 627876
rect 527836 627814 528508 627874
rect 527836 627812 527842 627814
rect 528502 627812 528508 627814
rect 528572 627812 528578 627876
rect 579797 627738 579863 627741
rect 583520 627738 584960 627828
rect 579797 627736 584960 627738
rect 579797 627680 579802 627736
rect 579858 627680 584960 627736
rect 579797 627678 584960 627680
rect 579797 627675 579863 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3233 624882 3299 624885
rect -960 624880 3299 624882
rect -960 624824 3238 624880
rect 3294 624824 3299 624880
rect -960 624822 3299 624824
rect -960 624732 480 624822
rect 3233 624819 3299 624822
rect 527214 623052 527220 623116
rect 527284 623114 527290 623116
rect 528134 623114 528140 623116
rect 527284 623054 528140 623114
rect 527284 623052 527290 623054
rect 528134 623052 528140 623054
rect 528204 623052 528210 623116
rect 527582 618292 527588 618356
rect 527652 618354 527658 618356
rect 528502 618354 528508 618356
rect 527652 618294 528508 618354
rect 527652 618292 527658 618294
rect 528502 618292 528508 618294
rect 528572 618292 528578 618356
rect 528134 618156 528140 618220
rect 528204 618218 528210 618220
rect 528686 618218 528692 618220
rect 528204 618158 528692 618218
rect 528204 618156 528210 618158
rect 528686 618156 528692 618158
rect 528756 618156 528762 618220
rect 527214 618020 527220 618084
rect 527284 618082 527290 618084
rect 527582 618082 527588 618084
rect 527284 618022 527588 618082
rect 527284 618020 527290 618022
rect 527582 618020 527588 618022
rect 527652 618020 527658 618084
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 2773 610466 2839 610469
rect -960 610464 2839 610466
rect -960 610408 2778 610464
rect 2834 610408 2839 610464
rect -960 610406 2839 610408
rect -960 610316 480 610406
rect 2773 610403 2839 610406
rect 527214 608636 527220 608700
rect 527284 608698 527290 608700
rect 527950 608698 527956 608700
rect 527284 608638 527956 608698
rect 527284 608636 527290 608638
rect 527950 608636 527956 608638
rect 528020 608636 528026 608700
rect 528318 608636 528324 608700
rect 528388 608698 528394 608700
rect 528686 608698 528692 608700
rect 528388 608638 528692 608698
rect 528388 608636 528394 608638
rect 528686 608636 528692 608638
rect 528756 608636 528762 608700
rect 579797 604210 579863 604213
rect 583520 604210 584960 604300
rect 579797 604208 584960 604210
rect 579797 604152 579802 604208
rect 579858 604152 584960 604208
rect 579797 604150 584960 604152
rect 579797 604147 579863 604150
rect 583520 604060 584960 604150
rect 527582 603740 527588 603804
rect 527652 603802 527658 603804
rect 528318 603802 528324 603804
rect 527652 603742 528324 603802
rect 527652 603740 527658 603742
rect 528318 603740 528324 603742
rect 528388 603740 528394 603804
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 579797 592514 579863 592517
rect 583520 592514 584960 592604
rect 579797 592512 584960 592514
rect 579797 592456 579802 592512
rect 579858 592456 584960 592512
rect 579797 592454 584960 592456
rect 579797 592451 579863 592454
rect 583520 592364 584960 592454
rect 527214 587148 527220 587212
rect 527284 587210 527290 587212
rect 527950 587210 527956 587212
rect 527284 587150 527956 587210
rect 527284 587148 527290 587150
rect 527950 587148 527956 587150
rect 528020 587148 528026 587212
rect -960 581620 480 581860
rect 583520 580818 584960 580908
rect 583342 580758 584960 580818
rect 538262 579942 547890 580002
rect 527398 579804 527404 579868
rect 527468 579866 527474 579868
rect 527468 579806 538138 579866
rect 527468 579804 527474 579806
rect 538078 579730 538138 579806
rect 538262 579730 538322 579942
rect 547830 579866 547890 579942
rect 557582 579942 567210 580002
rect 547830 579806 557458 579866
rect 538078 579670 538322 579730
rect 557398 579730 557458 579806
rect 557582 579730 557642 579942
rect 567150 579866 567210 579942
rect 567150 579806 576778 579866
rect 557398 579670 557642 579730
rect 576718 579730 576778 579806
rect 583342 579730 583402 580758
rect 583520 580668 584960 580758
rect 576718 579670 583402 579730
rect 527950 579532 527956 579596
rect 528020 579594 528026 579596
rect 528318 579594 528324 579596
rect 528020 579534 528324 579594
rect 528020 579532 528026 579534
rect 528318 579532 528324 579534
rect 528388 579532 528394 579596
rect 528318 570210 528324 570212
rect 527774 570150 528324 570210
rect 527774 570076 527834 570150
rect 528318 570148 528324 570150
rect 528388 570148 528394 570212
rect 527766 570012 527772 570076
rect 527836 570012 527842 570076
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3233 567354 3299 567357
rect -960 567352 3299 567354
rect -960 567296 3238 567352
rect 3294 567296 3299 567352
rect -960 567294 3299 567296
rect -960 567204 480 567294
rect 3233 567291 3299 567294
rect 527766 563076 527772 563140
rect 527836 563076 527842 563140
rect 527774 562866 527834 563076
rect 527950 562866 527956 562868
rect 527774 562806 527956 562866
rect 527950 562804 527956 562806
rect 528020 562804 528026 562868
rect 527398 560220 527404 560284
rect 527468 560282 527474 560284
rect 527950 560282 527956 560284
rect 527468 560222 527956 560282
rect 527468 560220 527474 560222
rect 527950 560220 527956 560222
rect 528020 560220 528026 560284
rect 579797 557290 579863 557293
rect 583520 557290 584960 557380
rect 579797 557288 584960 557290
rect 579797 557232 579802 557288
rect 579858 557232 584960 557288
rect 579797 557230 584960 557232
rect 579797 557227 579863 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 2773 553074 2839 553077
rect -960 553072 2839 553074
rect -960 553016 2778 553072
rect 2834 553016 2839 553072
rect -960 553014 2839 553016
rect -960 552924 480 553014
rect 2773 553011 2839 553014
rect 527398 550836 527404 550900
rect 527468 550898 527474 550900
rect 527468 550838 527834 550898
rect 527468 550836 527474 550838
rect 527774 550764 527834 550838
rect 527766 550700 527772 550764
rect 527836 550700 527842 550764
rect 579797 545594 579863 545597
rect 583520 545594 584960 545684
rect 579797 545592 584960 545594
rect 579797 545536 579802 545592
rect 579858 545536 584960 545592
rect 579797 545534 584960 545536
rect 579797 545531 579863 545534
rect 583520 545444 584960 545534
rect 527766 543962 527772 543964
rect 527222 543902 527772 543962
rect 527222 543556 527282 543902
rect 527766 543900 527772 543902
rect 527836 543900 527842 543964
rect 527214 543492 527220 543556
rect 527284 543492 527290 543556
rect -960 538658 480 538748
rect 3233 538658 3299 538661
rect -960 538656 3299 538658
rect -960 538600 3238 538656
rect 3294 538600 3299 538656
rect -960 538598 3299 538600
rect -960 538508 480 538598
rect 3233 538595 3299 538598
rect 527214 533972 527220 534036
rect 527284 534034 527290 534036
rect 528134 534034 528140 534036
rect 527284 533974 528140 534034
rect 527284 533972 527290 533974
rect 528134 533972 528140 533974
rect 528204 533972 528210 534036
rect 579797 533898 579863 533901
rect 583520 533898 584960 533988
rect 579797 533896 584960 533898
rect 579797 533840 579802 533896
rect 579858 533840 584960 533896
rect 579797 533838 584960 533840
rect 579797 533835 579863 533838
rect 583520 533748 584960 533838
rect 528134 524650 528140 524652
rect 527958 524590 528140 524650
rect -960 524092 480 524332
rect 527958 524244 528018 524590
rect 528134 524588 528140 524590
rect 528204 524588 528210 524652
rect 527950 524180 527956 524244
rect 528020 524180 528026 524244
rect 583520 521916 584960 522156
rect 527214 521596 527220 521660
rect 527284 521658 527290 521660
rect 527950 521658 527956 521660
rect 527284 521598 527956 521658
rect 527284 521596 527290 521598
rect 527950 521596 527956 521598
rect 528020 521596 528026 521660
rect 527214 512212 527220 512276
rect 527284 512274 527290 512276
rect 527284 512214 527650 512274
rect 527284 512212 527290 512214
rect 527590 512140 527650 512214
rect 527582 512076 527588 512140
rect 527652 512076 527658 512140
rect 579797 510370 579863 510373
rect 583520 510370 584960 510460
rect 579797 510368 584960 510370
rect 579797 510312 579802 510368
rect 579858 510312 584960 510368
rect 579797 510310 584960 510312
rect 579797 510307 579863 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3233 509962 3299 509965
rect -960 509960 3299 509962
rect -960 509904 3238 509960
rect 3294 509904 3299 509960
rect -960 509902 3299 509904
rect -960 509812 480 509902
rect 3233 509899 3299 509902
rect 527582 505140 527588 505204
rect 527652 505140 527658 505204
rect 527590 504930 527650 505140
rect 527766 504930 527772 504932
rect 527590 504870 527772 504930
rect 527766 504868 527772 504870
rect 527836 504868 527842 504932
rect 527398 502284 527404 502348
rect 527468 502346 527474 502348
rect 527766 502346 527772 502348
rect 527468 502286 527772 502346
rect 527468 502284 527474 502286
rect 527766 502284 527772 502286
rect 527836 502284 527842 502348
rect 579797 498674 579863 498677
rect 583520 498674 584960 498764
rect 579797 498672 584960 498674
rect 579797 498616 579802 498672
rect 579858 498616 584960 498672
rect 579797 498614 584960 498616
rect 579797 498611 579863 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 2773 495546 2839 495549
rect -960 495544 2839 495546
rect -960 495488 2778 495544
rect 2834 495488 2839 495544
rect -960 495486 2839 495488
rect -960 495396 480 495486
rect 2773 495483 2839 495486
rect 527398 492628 527404 492692
rect 527468 492690 527474 492692
rect 527950 492690 527956 492692
rect 527468 492630 527956 492690
rect 527468 492628 527474 492630
rect 527950 492628 527956 492630
rect 528020 492628 528026 492692
rect 579797 486842 579863 486845
rect 583520 486842 584960 486932
rect 579797 486840 584960 486842
rect 579797 486784 579802 486840
rect 579858 486784 584960 486840
rect 579797 486782 584960 486784
rect 579797 486779 579863 486782
rect 583520 486692 584960 486782
rect 527950 485890 527956 485892
rect 527774 485830 527956 485890
rect 527774 485620 527834 485830
rect 527950 485828 527956 485830
rect 528020 485828 528026 485892
rect 527766 485556 527772 485620
rect 527836 485556 527842 485620
rect 527766 482836 527772 482900
rect 527836 482898 527842 482900
rect 528134 482898 528140 482900
rect 527836 482838 528140 482898
rect 527836 482836 527842 482838
rect 528134 482836 528140 482838
rect 528204 482836 528210 482900
rect -960 481130 480 481220
rect 3233 481130 3299 481133
rect -960 481128 3299 481130
rect -960 481072 3238 481128
rect 3294 481072 3299 481128
rect -960 481070 3299 481072
rect -960 480980 480 481070
rect 3233 481067 3299 481070
rect 583520 474996 584960 475236
rect 527582 473316 527588 473380
rect 527652 473378 527658 473380
rect 528134 473378 528140 473380
rect 527652 473318 528140 473378
rect 527652 473316 527658 473318
rect 528134 473316 528140 473318
rect 528204 473316 528210 473380
rect -960 466700 480 466940
rect 527214 466244 527220 466308
rect 527284 466306 527290 466308
rect 527582 466306 527588 466308
rect 527284 466246 527588 466306
rect 527284 466244 527290 466246
rect 527582 466244 527588 466246
rect 527652 466244 527658 466308
rect 579797 463450 579863 463453
rect 583520 463450 584960 463540
rect 579797 463448 584960 463450
rect 579797 463392 579802 463448
rect 579858 463392 584960 463448
rect 579797 463390 584960 463392
rect 579797 463387 579863 463390
rect 583520 463300 584960 463390
rect 527214 456724 527220 456788
rect 527284 456786 527290 456788
rect 527766 456786 527772 456788
rect 527284 456726 527772 456786
rect 527284 456724 527290 456726
rect 527766 456724 527772 456726
rect 527836 456724 527842 456788
rect -960 452434 480 452524
rect 3141 452434 3207 452437
rect -960 452432 3207 452434
rect -960 452376 3146 452432
rect 3202 452376 3207 452432
rect -960 452374 3207 452376
rect -960 452284 480 452374
rect 3141 452371 3207 452374
rect 579889 451754 579955 451757
rect 583520 451754 584960 451844
rect 579889 451752 584960 451754
rect 579889 451696 579894 451752
rect 579950 451696 584960 451752
rect 579889 451694 584960 451696
rect 579889 451691 579955 451694
rect 583520 451604 584960 451694
rect 527214 444348 527220 444412
rect 527284 444410 527290 444412
rect 527582 444410 527588 444412
rect 527284 444350 527588 444410
rect 527284 444348 527290 444350
rect 527582 444348 527588 444350
rect 527652 444348 527658 444412
rect 579889 439922 579955 439925
rect 583520 439922 584960 440012
rect 579889 439920 584960 439922
rect 579889 439864 579894 439920
rect 579950 439864 584960 439920
rect 579889 439862 584960 439864
rect 579889 439859 579955 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 527214 437412 527220 437476
rect 527284 437474 527290 437476
rect 527950 437474 527956 437476
rect 527284 437414 527956 437474
rect 527284 437412 527290 437414
rect 527950 437412 527956 437414
rect 528020 437412 528026 437476
rect 583520 428076 584960 428316
rect 527950 427954 527956 427956
rect 527774 427894 527956 427954
rect 527774 427684 527834 427894
rect 527950 427892 527956 427894
rect 528020 427892 528026 427956
rect 527766 427620 527772 427684
rect 527836 427620 527842 427684
rect 527766 424900 527772 424964
rect 527836 424900 527842 424964
rect 527398 424764 527404 424828
rect 527468 424826 527474 424828
rect 527774 424826 527834 424900
rect 527468 424766 527834 424826
rect 527468 424764 527474 424766
rect -960 423738 480 423828
rect 3325 423738 3391 423741
rect -960 423736 3391 423738
rect -960 423680 3330 423736
rect 3386 423680 3391 423736
rect -960 423678 3391 423680
rect -960 423588 480 423678
rect 3325 423675 3391 423678
rect 579889 416530 579955 416533
rect 583520 416530 584960 416620
rect 579889 416528 584960 416530
rect 579889 416472 579894 416528
rect 579950 416472 584960 416528
rect 579889 416470 584960 416472
rect 579889 416467 579955 416470
rect 583520 416380 584960 416470
rect 527398 415380 527404 415444
rect 527468 415442 527474 415444
rect 527950 415442 527956 415444
rect 527468 415382 527956 415442
rect 527468 415380 527474 415382
rect 527950 415380 527956 415382
rect 528020 415380 528026 415444
rect -960 409172 480 409412
rect 527950 408642 527956 408644
rect 527774 408582 527956 408642
rect 527774 408372 527834 408582
rect 527950 408580 527956 408582
rect 528020 408580 528026 408644
rect 527766 408308 527772 408372
rect 527836 408308 527842 408372
rect 527214 405588 527220 405652
rect 527284 405650 527290 405652
rect 527766 405650 527772 405652
rect 527284 405590 527772 405650
rect 527284 405588 527290 405590
rect 527766 405588 527772 405590
rect 527836 405588 527842 405652
rect 579889 404834 579955 404837
rect 583520 404834 584960 404924
rect 579889 404832 584960 404834
rect 579889 404776 579894 404832
rect 579950 404776 584960 404832
rect 579889 404774 584960 404776
rect 579889 404771 579955 404774
rect 583520 404684 584960 404774
rect 527214 396068 527220 396132
rect 527284 396130 527290 396132
rect 527582 396130 527588 396132
rect 527284 396070 527588 396130
rect 527284 396068 527290 396070
rect 527582 396068 527588 396070
rect 527652 396068 527658 396132
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 579889 393002 579955 393005
rect 583520 393002 584960 393092
rect 579889 393000 584960 393002
rect 579889 392944 579894 393000
rect 579950 392944 584960 393000
rect 579889 392942 584960 392944
rect 579889 392939 579955 392942
rect 583520 392852 584960 392942
rect 527582 389330 527588 389332
rect 527406 389270 527588 389330
rect 527406 389060 527466 389270
rect 527582 389268 527588 389270
rect 527652 389268 527658 389332
rect 527398 388996 527404 389060
rect 527468 388996 527474 389060
rect 527398 386276 527404 386340
rect 527468 386276 527474 386340
rect 527406 386202 527466 386276
rect 527950 386202 527956 386204
rect 527406 386142 527956 386202
rect 527950 386140 527956 386142
rect 528020 386140 528026 386204
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 2773 380626 2839 380629
rect -960 380624 2839 380626
rect -960 380568 2778 380624
rect 2834 380568 2839 380624
rect -960 380566 2839 380568
rect -960 380476 480 380566
rect 2773 380563 2839 380566
rect 527582 376756 527588 376820
rect 527652 376818 527658 376820
rect 527950 376818 527956 376820
rect 527652 376758 527956 376818
rect 527652 376756 527658 376758
rect 527950 376756 527956 376758
rect 528020 376756 528026 376820
rect 527582 369956 527588 370020
rect 527652 369956 527658 370020
rect 527590 369746 527650 369956
rect 527766 369746 527772 369748
rect 527590 369686 527772 369746
rect 527766 369684 527772 369686
rect 527836 369684 527842 369748
rect 579981 369610 580047 369613
rect 583520 369610 584960 369700
rect 579981 369608 584960 369610
rect 579981 369552 579986 369608
rect 580042 369552 584960 369608
rect 579981 369550 584960 369552
rect 579981 369547 580047 369550
rect 583520 369460 584960 369550
rect 527766 366964 527772 367028
rect 527836 366964 527842 367028
rect 527774 366890 527834 366964
rect 528318 366890 528324 366892
rect 527774 366830 528324 366890
rect 528318 366828 528324 366830
rect 528388 366828 528394 366892
rect -960 366210 480 366300
rect 3325 366210 3391 366213
rect -960 366208 3391 366210
rect -960 366152 3330 366208
rect 3386 366152 3391 366208
rect -960 366150 3391 366152
rect -960 366060 480 366150
rect 3325 366147 3391 366150
rect 580073 357914 580139 357917
rect 583520 357914 584960 358004
rect 580073 357912 584960 357914
rect 580073 357856 580078 357912
rect 580134 357856 584960 357912
rect 580073 357854 584960 357856
rect 580073 357851 580139 357854
rect 583520 357764 584960 357854
rect 527950 357444 527956 357508
rect 528020 357506 528026 357508
rect 528318 357506 528324 357508
rect 528020 357446 528324 357506
rect 528020 357444 528026 357446
rect 528318 357444 528324 357446
rect 528388 357444 528394 357508
rect -960 351780 480 352020
rect 527950 350706 527956 350708
rect 527774 350646 527956 350706
rect 527774 350436 527834 350646
rect 527950 350644 527956 350646
rect 528020 350644 528026 350708
rect 527766 350372 527772 350436
rect 527836 350372 527842 350436
rect 527766 347652 527772 347716
rect 527836 347714 527842 347716
rect 528318 347714 528324 347716
rect 527836 347654 528324 347714
rect 527836 347652 527842 347654
rect 528318 347652 528324 347654
rect 528388 347652 528394 347716
rect 579797 346082 579863 346085
rect 583520 346082 584960 346172
rect 579797 346080 584960 346082
rect 579797 346024 579802 346080
rect 579858 346024 584960 346080
rect 579797 346022 584960 346024
rect 579797 346019 579863 346022
rect 583520 345932 584960 346022
rect 527582 340308 527588 340372
rect 527652 340370 527658 340372
rect 528318 340370 528324 340372
rect 527652 340310 528324 340370
rect 527652 340308 527658 340310
rect 528318 340308 528324 340310
rect 528388 340308 528394 340372
rect -960 337514 480 337604
rect 3233 337514 3299 337517
rect -960 337512 3299 337514
rect -960 337456 3238 337512
rect 3294 337456 3299 337512
rect -960 337454 3299 337456
rect -960 337364 480 337454
rect 3233 337451 3299 337454
rect 365805 337514 365871 337517
rect 378501 337514 378567 337517
rect 365805 337512 378567 337514
rect 365805 337456 365810 337512
rect 365866 337456 378506 337512
rect 378562 337456 378567 337512
rect 365805 337454 378567 337456
rect 365805 337451 365871 337454
rect 378501 337451 378567 337454
rect 10317 337378 10383 337381
rect 232405 337378 232471 337381
rect 10317 337376 232471 337378
rect 10317 337320 10322 337376
rect 10378 337320 232410 337376
rect 232466 337320 232471 337376
rect 10317 337318 232471 337320
rect 10317 337315 10383 337318
rect 232405 337315 232471 337318
rect 528185 337378 528251 337381
rect 565077 337378 565143 337381
rect 528185 337376 565143 337378
rect 528185 337320 528190 337376
rect 528246 337320 565082 337376
rect 565138 337320 565143 337376
rect 528185 337318 565143 337320
rect 528185 337315 528251 337318
rect 565077 337315 565143 337318
rect 527582 336636 527588 336700
rect 527652 336636 527658 336700
rect 527449 336562 527515 336565
rect 527590 336562 527650 336636
rect 527449 336560 527650 336562
rect 527449 336504 527454 336560
rect 527510 336504 527650 336560
rect 527449 336502 527650 336504
rect 527449 336499 527515 336502
rect 277669 335338 277735 335341
rect 277945 335338 278011 335341
rect 277669 335336 278011 335338
rect 277669 335280 277674 335336
rect 277730 335280 277950 335336
rect 278006 335280 278011 335336
rect 277669 335278 278011 335280
rect 277669 335275 277735 335278
rect 277945 335275 278011 335278
rect 294045 335338 294111 335341
rect 294321 335338 294387 335341
rect 294045 335336 294387 335338
rect 294045 335280 294050 335336
rect 294106 335280 294326 335336
rect 294382 335280 294387 335336
rect 294045 335278 294387 335280
rect 294045 335275 294111 335278
rect 294321 335275 294387 335278
rect 583520 334236 584960 334476
rect 327441 328674 327507 328677
rect 428365 328674 428431 328677
rect 327030 328672 327507 328674
rect 327030 328616 327446 328672
rect 327502 328616 327507 328672
rect 327030 328614 327507 328616
rect 327030 328538 327090 328614
rect 327441 328611 327507 328614
rect 427862 328672 428431 328674
rect 427862 328616 428370 328672
rect 428426 328616 428431 328672
rect 427862 328614 428431 328616
rect 327165 328538 327231 328541
rect 327030 328536 327231 328538
rect 327030 328480 327170 328536
rect 327226 328480 327231 328536
rect 327030 328478 327231 328480
rect 427862 328538 427922 328614
rect 428365 328611 428431 328614
rect 427997 328538 428063 328541
rect 427862 328536 428063 328538
rect 427862 328480 428002 328536
rect 428058 328480 428063 328536
rect 427862 328478 428063 328480
rect 327165 328475 327231 328478
rect 427997 328475 428063 328478
rect 332685 328404 332751 328405
rect 332685 328402 332732 328404
rect 332640 328400 332732 328402
rect 332640 328344 332690 328400
rect 332640 328342 332732 328344
rect 332685 328340 332732 328342
rect 332796 328340 332802 328404
rect 332685 328339 332751 328340
rect 243537 327314 243603 327317
rect 242942 327312 243603 327314
rect 242942 327256 243542 327312
rect 243598 327256 243603 327312
rect 242942 327254 243603 327256
rect 242942 327178 243002 327254
rect 243537 327251 243603 327254
rect 243077 327178 243143 327181
rect 242942 327176 243143 327178
rect 242942 327120 243082 327176
rect 243138 327120 243143 327176
rect 242942 327118 243143 327120
rect 243077 327115 243143 327118
rect 277669 325682 277735 325685
rect 277853 325682 277919 325685
rect 277669 325680 277919 325682
rect 277669 325624 277674 325680
rect 277730 325624 277858 325680
rect 277914 325624 277919 325680
rect 277669 325622 277919 325624
rect 277669 325619 277735 325622
rect 277853 325619 277919 325622
rect 357617 325682 357683 325685
rect 357801 325682 357867 325685
rect 357617 325680 357867 325682
rect 357617 325624 357622 325680
rect 357678 325624 357806 325680
rect 357862 325624 357867 325680
rect 357617 325622 357867 325624
rect 357617 325619 357683 325622
rect 357801 325619 357867 325622
rect 451549 325682 451615 325685
rect 451733 325682 451799 325685
rect 451549 325680 451799 325682
rect 451549 325624 451554 325680
rect 451610 325624 451738 325680
rect 451794 325624 451799 325680
rect 451549 325622 451799 325624
rect 451549 325619 451615 325622
rect 451733 325619 451799 325622
rect -960 323098 480 323188
rect 2773 323098 2839 323101
rect -960 323096 2839 323098
rect -960 323040 2778 323096
rect 2834 323040 2839 323096
rect -960 323038 2839 323040
rect -960 322948 480 323038
rect 2773 323035 2839 323038
rect 580073 322690 580139 322693
rect 583520 322690 584960 322780
rect 580073 322688 584960 322690
rect 580073 322632 580078 322688
rect 580134 322632 584960 322688
rect 580073 322630 584960 322632
rect 580073 322627 580139 322630
rect 583520 322540 584960 322630
rect 261017 319018 261083 319021
rect 260974 319016 261083 319018
rect 260974 318960 261022 319016
rect 261078 318960 261083 319016
rect 260974 318955 261083 318960
rect 332726 318956 332732 319020
rect 332796 319018 332802 319020
rect 527449 319018 527515 319021
rect 332796 318958 332978 319018
rect 332796 318956 332802 318958
rect 260974 318885 261034 318955
rect 260974 318880 261083 318885
rect 260974 318824 261022 318880
rect 261078 318824 261083 318880
rect 260974 318822 261083 318824
rect 261017 318819 261083 318822
rect 332777 318882 332843 318885
rect 332918 318882 332978 318958
rect 527406 319016 527515 319018
rect 527406 318960 527454 319016
rect 527510 318960 527515 319016
rect 527406 318955 527515 318960
rect 527406 318884 527466 318955
rect 332777 318880 332978 318882
rect 332777 318824 332782 318880
rect 332838 318824 332978 318880
rect 332777 318822 332978 318824
rect 332777 318819 332843 318822
rect 527398 318820 527404 318884
rect 527468 318820 527474 318884
rect 324221 318746 324287 318749
rect 324405 318746 324471 318749
rect 324221 318744 324471 318746
rect 324221 318688 324226 318744
rect 324282 318688 324410 318744
rect 324466 318688 324471 318744
rect 324221 318686 324471 318688
rect 324221 318683 324287 318686
rect 324405 318683 324471 318686
rect 255589 316026 255655 316029
rect 255773 316026 255839 316029
rect 255589 316024 255839 316026
rect 255589 315968 255594 316024
rect 255650 315968 255778 316024
rect 255834 315968 255839 316024
rect 255589 315966 255839 315968
rect 255589 315963 255655 315966
rect 255773 315963 255839 315966
rect 365805 316026 365871 316029
rect 365989 316026 366055 316029
rect 365805 316024 366055 316026
rect 365805 315968 365810 316024
rect 365866 315968 365994 316024
rect 366050 315968 366055 316024
rect 365805 315966 366055 315968
rect 365805 315963 365871 315966
rect 365989 315963 366055 315966
rect 527398 312020 527404 312084
rect 527468 312020 527474 312084
rect 527406 311810 527466 312020
rect 527582 311810 527588 311812
rect 527406 311750 527588 311810
rect 527582 311748 527588 311750
rect 527652 311748 527658 311812
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect 527633 309092 527699 309093
rect 232998 309090 233004 309092
rect 614 309030 233004 309090
rect -960 308818 480 308908
rect 614 308818 674 309030
rect 232998 309028 233004 309030
rect 233068 309028 233074 309092
rect 527582 309028 527588 309092
rect 527652 309090 527699 309092
rect 527652 309088 527744 309090
rect 527694 309032 527744 309088
rect 527652 309030 527744 309032
rect 527652 309028 527699 309030
rect 527633 309027 527699 309028
rect -960 308758 674 308818
rect -960 308668 480 308758
rect 249241 307730 249307 307733
rect 249374 307730 249380 307732
rect 249241 307728 249380 307730
rect 249241 307672 249246 307728
rect 249302 307672 249380 307728
rect 249241 307670 249380 307672
rect 249241 307667 249307 307670
rect 249374 307668 249380 307670
rect 249444 307668 249450 307732
rect 261017 307730 261083 307733
rect 261201 307730 261267 307733
rect 261017 307728 261267 307730
rect 261017 307672 261022 307728
rect 261078 307672 261206 307728
rect 261262 307672 261267 307728
rect 261017 307670 261267 307672
rect 261017 307667 261083 307670
rect 261201 307667 261267 307670
rect 527398 302092 527404 302156
rect 527468 302154 527474 302156
rect 527633 302154 527699 302157
rect 527468 302152 527699 302154
rect 527468 302096 527638 302152
rect 527694 302096 527699 302152
rect 527468 302094 527699 302096
rect 527468 302092 527474 302094
rect 527633 302091 527699 302094
rect 309409 299434 309475 299437
rect 309593 299434 309659 299437
rect 309409 299432 309659 299434
rect 309409 299376 309414 299432
rect 309470 299376 309598 299432
rect 309654 299376 309659 299432
rect 309409 299374 309659 299376
rect 309409 299371 309475 299374
rect 309593 299371 309659 299374
rect 580901 299162 580967 299165
rect 583520 299162 584960 299252
rect 580901 299160 584960 299162
rect 580901 299104 580906 299160
rect 580962 299104 584960 299160
rect 580901 299102 584960 299104
rect 580901 299099 580967 299102
rect 583520 299012 584960 299102
rect 249241 298346 249307 298349
rect 249198 298344 249307 298346
rect 249198 298288 249246 298344
rect 249302 298288 249307 298344
rect 249198 298283 249307 298288
rect 357709 298346 357775 298349
rect 357709 298344 357818 298346
rect 357709 298288 357714 298344
rect 357770 298288 357818 298344
rect 357709 298283 357818 298288
rect 249198 298212 249258 298283
rect 249190 298148 249196 298212
rect 249260 298148 249266 298212
rect 357617 298210 357683 298213
rect 357758 298210 357818 298283
rect 357617 298208 357818 298210
rect 357617 298152 357622 298208
rect 357678 298152 357818 298208
rect 357617 298150 357818 298152
rect 357617 298147 357683 298150
rect 254301 296714 254367 296717
rect 254485 296714 254551 296717
rect 254301 296712 254551 296714
rect 254301 296656 254306 296712
rect 254362 296656 254490 296712
rect 254546 296656 254551 296712
rect 254301 296654 254551 296656
rect 254301 296651 254367 296654
rect 254485 296651 254551 296654
rect 357617 296714 357683 296717
rect 357801 296714 357867 296717
rect 357617 296712 357867 296714
rect 357617 296656 357622 296712
rect 357678 296656 357806 296712
rect 357862 296656 357867 296712
rect 357617 296654 357867 296656
rect 357617 296651 357683 296654
rect 357801 296651 357867 296654
rect -960 294402 480 294492
rect 3325 294402 3391 294405
rect -960 294400 3391 294402
rect -960 294344 3330 294400
rect 3386 294344 3391 294400
rect -960 294342 3391 294344
rect -960 294252 480 294342
rect 3325 294339 3391 294342
rect 249190 289852 249196 289916
rect 249260 289852 249266 289916
rect 249198 289642 249258 289852
rect 281625 289778 281691 289781
rect 281901 289778 281967 289781
rect 281625 289776 281967 289778
rect 281625 289720 281630 289776
rect 281686 289720 281906 289776
rect 281962 289720 281967 289776
rect 281625 289718 281967 289720
rect 281625 289715 281691 289718
rect 281901 289715 281967 289718
rect 324497 289778 324563 289781
rect 324681 289778 324747 289781
rect 527633 289780 527699 289781
rect 324497 289776 324747 289778
rect 324497 289720 324502 289776
rect 324558 289720 324686 289776
rect 324742 289720 324747 289776
rect 324497 289718 324747 289720
rect 324497 289715 324563 289718
rect 324681 289715 324747 289718
rect 527582 289716 527588 289780
rect 527652 289778 527699 289780
rect 527652 289776 527744 289778
rect 527694 289720 527744 289776
rect 527652 289718 527744 289720
rect 527652 289716 527699 289718
rect 527633 289715 527699 289716
rect 249558 289642 249564 289644
rect 249198 289582 249564 289642
rect 249558 289580 249564 289582
rect 249628 289580 249634 289644
rect 236453 288418 236519 288421
rect 236637 288418 236703 288421
rect 236453 288416 236703 288418
rect 236453 288360 236458 288416
rect 236514 288360 236642 288416
rect 236698 288360 236703 288416
rect 236453 288358 236703 288360
rect 236453 288355 236519 288358
rect 236637 288355 236703 288358
rect 451273 288418 451339 288421
rect 451457 288418 451523 288421
rect 451273 288416 451523 288418
rect 451273 288360 451278 288416
rect 451334 288360 451462 288416
rect 451518 288360 451523 288416
rect 451273 288358 451523 288360
rect 451273 288355 451339 288358
rect 451457 288355 451523 288358
rect 583520 287316 584960 287556
rect 527633 280394 527699 280397
rect 527406 280392 527699 280394
rect 527406 280336 527638 280392
rect 527694 280336 527699 280392
rect 527406 280334 527699 280336
rect 527406 280260 527466 280334
rect 527633 280331 527699 280334
rect -960 280122 480 280212
rect 527398 280196 527404 280260
rect 527468 280196 527474 280260
rect 3141 280122 3207 280125
rect 281717 280122 281783 280125
rect -960 280120 3207 280122
rect -960 280064 3146 280120
rect 3202 280064 3207 280120
rect -960 280062 3207 280064
rect -960 279972 480 280062
rect 3141 280059 3207 280062
rect 281582 280120 281783 280122
rect 281582 280064 281722 280120
rect 281778 280064 281783 280120
rect 281582 280062 281783 280064
rect 281582 279986 281642 280062
rect 281717 280059 281783 280062
rect 309409 280122 309475 280125
rect 309593 280122 309659 280125
rect 309409 280120 309659 280122
rect 309409 280064 309414 280120
rect 309470 280064 309598 280120
rect 309654 280064 309659 280120
rect 309409 280062 309659 280064
rect 309409 280059 309475 280062
rect 309593 280059 309659 280062
rect 397729 280122 397795 280125
rect 397729 280120 397930 280122
rect 397729 280064 397734 280120
rect 397790 280064 397930 280120
rect 397729 280062 397930 280064
rect 397729 280059 397795 280062
rect 281809 279986 281875 279989
rect 281582 279984 281875 279986
rect 281582 279928 281814 279984
rect 281870 279928 281875 279984
rect 281582 279926 281875 279928
rect 281809 279923 281875 279926
rect 397361 279986 397427 279989
rect 397870 279986 397930 280062
rect 397361 279984 397930 279986
rect 397361 279928 397366 279984
rect 397422 279928 397930 279984
rect 397361 279926 397930 279928
rect 397361 279923 397427 279926
rect 249241 279852 249307 279853
rect 249190 279850 249196 279852
rect 249150 279790 249196 279850
rect 249260 279848 249307 279852
rect 249302 279792 249307 279848
rect 249190 279788 249196 279790
rect 249260 279788 249307 279792
rect 249241 279787 249307 279788
rect 298277 278762 298343 278765
rect 298553 278762 298619 278765
rect 298277 278760 298619 278762
rect 298277 278704 298282 278760
rect 298338 278704 298558 278760
rect 298614 278704 298619 278760
rect 298277 278702 298619 278704
rect 298277 278699 298343 278702
rect 298553 278699 298619 278702
rect 369945 278762 370011 278765
rect 370313 278762 370379 278765
rect 369945 278760 370379 278762
rect 369945 278704 369950 278760
rect 370006 278704 370318 278760
rect 370374 278704 370379 278760
rect 369945 278702 370379 278704
rect 369945 278699 370011 278702
rect 370313 278699 370379 278702
rect 259361 277402 259427 277405
rect 259729 277402 259795 277405
rect 259361 277400 259795 277402
rect 259361 277344 259366 277400
rect 259422 277344 259734 277400
rect 259790 277344 259795 277400
rect 259361 277342 259795 277344
rect 259361 277339 259427 277342
rect 259729 277339 259795 277342
rect 347865 277402 347931 277405
rect 348049 277402 348115 277405
rect 347865 277400 348115 277402
rect 347865 277344 347870 277400
rect 347926 277344 348054 277400
rect 348110 277344 348115 277400
rect 347865 277342 348115 277344
rect 347865 277339 347931 277342
rect 348049 277339 348115 277342
rect 580809 275770 580875 275773
rect 583520 275770 584960 275860
rect 580809 275768 584960 275770
rect 580809 275712 580814 275768
rect 580870 275712 584960 275768
rect 580809 275710 584960 275712
rect 580809 275707 580875 275710
rect 583520 275620 584960 275710
rect 527398 273396 527404 273460
rect 527468 273396 527474 273460
rect 527406 273050 527466 273396
rect 527582 273050 527588 273052
rect 527406 272990 527588 273050
rect 527582 272988 527588 272990
rect 527652 272988 527658 273052
rect 358997 270738 359063 270741
rect 358862 270736 359063 270738
rect 358862 270680 359002 270736
rect 359058 270680 359063 270736
rect 358862 270678 359063 270680
rect 242801 270602 242867 270605
rect 249241 270602 249307 270605
rect 249374 270602 249380 270604
rect 242801 270600 243002 270602
rect 242801 270544 242806 270600
rect 242862 270544 243002 270600
rect 242801 270542 243002 270544
rect 242801 270539 242867 270542
rect 242942 270466 243002 270542
rect 249241 270600 249380 270602
rect 249241 270544 249246 270600
rect 249302 270544 249380 270600
rect 249241 270542 249380 270544
rect 249241 270539 249307 270542
rect 249374 270540 249380 270542
rect 249444 270540 249450 270604
rect 331121 270602 331187 270605
rect 331121 270600 331322 270602
rect 331121 270544 331126 270600
rect 331182 270544 331322 270600
rect 331121 270542 331322 270544
rect 331121 270539 331187 270542
rect 331262 270469 331322 270542
rect 358862 270469 358922 270678
rect 358997 270675 359063 270678
rect 386781 270602 386847 270605
rect 386646 270600 386847 270602
rect 386646 270544 386786 270600
rect 386842 270544 386847 270600
rect 386646 270542 386847 270544
rect 386646 270469 386706 270542
rect 386781 270539 386847 270542
rect 243169 270466 243235 270469
rect 242942 270464 243235 270466
rect 242942 270408 243174 270464
rect 243230 270408 243235 270464
rect 242942 270406 243235 270408
rect 243169 270403 243235 270406
rect 249241 270466 249307 270469
rect 249374 270466 249380 270468
rect 249241 270464 249380 270466
rect 249241 270408 249246 270464
rect 249302 270408 249380 270464
rect 249241 270406 249380 270408
rect 249241 270403 249307 270406
rect 249374 270404 249380 270406
rect 249444 270404 249450 270468
rect 331262 270464 331371 270469
rect 331262 270408 331310 270464
rect 331366 270408 331371 270464
rect 331262 270406 331371 270408
rect 358862 270464 358971 270469
rect 358862 270408 358910 270464
rect 358966 270408 358971 270464
rect 358862 270406 358971 270408
rect 386646 270464 386755 270469
rect 386646 270408 386694 270464
rect 386750 270408 386755 270464
rect 386646 270406 386755 270408
rect 331305 270403 331371 270406
rect 358905 270403 358971 270406
rect 386689 270403 386755 270406
rect 527449 270466 527515 270469
rect 527582 270466 527588 270468
rect 527449 270464 527588 270466
rect 527449 270408 527454 270464
rect 527510 270408 527588 270464
rect 527449 270406 527588 270408
rect 527449 270403 527515 270406
rect 527582 270404 527588 270406
rect 527652 270404 527658 270468
rect 265157 269106 265223 269109
rect 265433 269106 265499 269109
rect 265157 269104 265499 269106
rect 265157 269048 265162 269104
rect 265218 269048 265438 269104
rect 265494 269048 265499 269104
rect 265157 269046 265499 269048
rect 265157 269043 265223 269046
rect 265433 269043 265499 269046
rect 352097 269106 352163 269109
rect 352281 269106 352347 269109
rect 352097 269104 352347 269106
rect 352097 269048 352102 269104
rect 352158 269048 352286 269104
rect 352342 269048 352347 269104
rect 352097 269046 352347 269048
rect 352097 269043 352163 269046
rect 352281 269043 352347 269046
rect -960 265706 480 265796
rect 3325 265706 3391 265709
rect -960 265704 3391 265706
rect -960 265648 3330 265704
rect 3386 265648 3391 265704
rect -960 265646 3391 265648
rect -960 265556 480 265646
rect 3325 265643 3391 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 527449 261082 527515 261085
rect 527406 261080 527515 261082
rect 527406 261024 527454 261080
rect 527510 261024 527515 261080
rect 527406 261019 527515 261024
rect 249241 260946 249307 260949
rect 527406 260948 527466 261019
rect 249198 260944 249307 260946
rect 249198 260888 249246 260944
rect 249302 260888 249307 260944
rect 249198 260883 249307 260888
rect 527398 260884 527404 260948
rect 527468 260884 527474 260948
rect 249198 260674 249258 260883
rect 270769 260810 270835 260813
rect 281809 260810 281875 260813
rect 281993 260810 282059 260813
rect 270769 260808 270970 260810
rect 270769 260752 270774 260808
rect 270830 260752 270970 260808
rect 270769 260750 270970 260752
rect 270769 260747 270835 260750
rect 249558 260674 249564 260676
rect 249198 260614 249564 260674
rect 249558 260612 249564 260614
rect 249628 260612 249634 260676
rect 270585 260674 270651 260677
rect 270910 260674 270970 260750
rect 281809 260808 282059 260810
rect 281809 260752 281814 260808
rect 281870 260752 281998 260808
rect 282054 260752 282059 260808
rect 281809 260750 282059 260752
rect 281809 260747 281875 260750
rect 281993 260747 282059 260750
rect 381169 260810 381235 260813
rect 381353 260810 381419 260813
rect 381169 260808 381419 260810
rect 381169 260752 381174 260808
rect 381230 260752 381358 260808
rect 381414 260752 381419 260808
rect 381169 260750 381419 260752
rect 381169 260747 381235 260750
rect 381353 260747 381419 260750
rect 270585 260672 270970 260674
rect 270585 260616 270590 260672
rect 270646 260616 270970 260672
rect 270585 260614 270970 260616
rect 270585 260611 270651 260614
rect 254025 259450 254091 259453
rect 254209 259450 254275 259453
rect 254025 259448 254275 259450
rect 254025 259392 254030 259448
rect 254086 259392 254214 259448
rect 254270 259392 254275 259448
rect 254025 259390 254275 259392
rect 254025 259387 254091 259390
rect 254209 259387 254275 259390
rect 259545 259450 259611 259453
rect 259729 259450 259795 259453
rect 259545 259448 259795 259450
rect 259545 259392 259550 259448
rect 259606 259392 259734 259448
rect 259790 259392 259795 259448
rect 259545 259390 259795 259392
rect 259545 259387 259611 259390
rect 259729 259387 259795 259390
rect 397361 259450 397427 259453
rect 397913 259450 397979 259453
rect 397361 259448 397979 259450
rect 397361 259392 397366 259448
rect 397422 259392 397918 259448
rect 397974 259392 397979 259448
rect 397361 259390 397979 259392
rect 397361 259387 397427 259390
rect 397913 259387 397979 259390
rect 408769 259450 408835 259453
rect 408953 259450 409019 259453
rect 408769 259448 409019 259450
rect 408769 259392 408774 259448
rect 408830 259392 408958 259448
rect 409014 259392 409019 259448
rect 408769 259390 409019 259392
rect 408769 259387 408835 259390
rect 408953 259387 409019 259390
rect 527398 253948 527404 254012
rect 527468 253948 527474 254012
rect 527406 253738 527466 253948
rect 527582 253738 527588 253740
rect 527406 253678 527588 253738
rect 527582 253676 527588 253678
rect 527652 253676 527658 253740
rect 3141 252514 3207 252517
rect 232814 252514 232820 252516
rect 3141 252512 232820 252514
rect 3141 252456 3146 252512
rect 3202 252456 232820 252512
rect 3141 252454 232820 252456
rect 3141 252451 3207 252454
rect 232814 252452 232820 252454
rect 232884 252452 232890 252516
rect 579613 252242 579679 252245
rect 583520 252242 584960 252332
rect 579613 252240 584960 252242
rect 579613 252184 579618 252240
rect 579674 252184 584960 252240
rect 579613 252182 584960 252184
rect 579613 252179 579679 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3141 251290 3207 251293
rect -960 251288 3207 251290
rect -960 251232 3146 251288
rect 3202 251232 3207 251288
rect -960 251230 3207 251232
rect -960 251140 480 251230
rect 3141 251227 3207 251230
rect 242801 251290 242867 251293
rect 331121 251290 331187 251293
rect 364241 251290 364307 251293
rect 242801 251288 243002 251290
rect 242801 251232 242806 251288
rect 242862 251232 243002 251288
rect 242801 251230 243002 251232
rect 242801 251227 242867 251230
rect 242942 251157 243002 251230
rect 331121 251288 331322 251290
rect 331121 251232 331126 251288
rect 331182 251232 331322 251288
rect 331121 251230 331322 251232
rect 331121 251227 331187 251230
rect 242942 251152 243051 251157
rect 242942 251096 242990 251152
rect 243046 251096 243051 251152
rect 242942 251094 243051 251096
rect 242985 251091 243051 251094
rect 249241 251154 249307 251157
rect 249374 251154 249380 251156
rect 249241 251152 249380 251154
rect 249241 251096 249246 251152
rect 249302 251096 249380 251152
rect 249241 251094 249380 251096
rect 249241 251091 249307 251094
rect 249374 251092 249380 251094
rect 249444 251092 249450 251156
rect 309317 251154 309383 251157
rect 309501 251154 309567 251157
rect 309317 251152 309567 251154
rect 309317 251096 309322 251152
rect 309378 251096 309506 251152
rect 309562 251096 309567 251152
rect 309317 251094 309567 251096
rect 309317 251091 309383 251094
rect 309501 251091 309567 251094
rect 331121 251154 331187 251157
rect 331262 251154 331322 251230
rect 364241 251288 364442 251290
rect 364241 251232 364246 251288
rect 364302 251232 364442 251288
rect 364241 251230 364442 251232
rect 364241 251227 364307 251230
rect 331121 251152 331322 251154
rect 331121 251096 331126 251152
rect 331182 251096 331322 251152
rect 331121 251094 331322 251096
rect 342437 251154 342503 251157
rect 342621 251154 342687 251157
rect 342437 251152 342687 251154
rect 342437 251096 342442 251152
rect 342498 251096 342626 251152
rect 342682 251096 342687 251152
rect 342437 251094 342687 251096
rect 331121 251091 331187 251094
rect 342437 251091 342503 251094
rect 342621 251091 342687 251094
rect 364241 251154 364307 251157
rect 364382 251154 364442 251230
rect 364241 251152 364442 251154
rect 364241 251096 364246 251152
rect 364302 251096 364442 251152
rect 364241 251094 364442 251096
rect 375557 251154 375623 251157
rect 375741 251154 375807 251157
rect 375557 251152 375807 251154
rect 375557 251096 375562 251152
rect 375618 251096 375746 251152
rect 375802 251096 375807 251152
rect 375557 251094 375807 251096
rect 364241 251091 364307 251094
rect 375557 251091 375623 251094
rect 375741 251091 375807 251094
rect 527449 251154 527515 251157
rect 527582 251154 527588 251156
rect 527449 251152 527588 251154
rect 527449 251096 527454 251152
rect 527510 251096 527588 251152
rect 527449 251094 527588 251096
rect 527449 251091 527515 251094
rect 527582 251092 527588 251094
rect 527652 251092 527658 251156
rect 392117 249794 392183 249797
rect 392393 249794 392459 249797
rect 392117 249792 392459 249794
rect 392117 249736 392122 249792
rect 392178 249736 392398 249792
rect 392454 249736 392459 249792
rect 392117 249734 392459 249736
rect 392117 249731 392183 249734
rect 392393 249731 392459 249734
rect 249241 241770 249307 241773
rect 527449 241770 527515 241773
rect 249198 241768 249307 241770
rect 249198 241712 249246 241768
rect 249302 241712 249307 241768
rect 249198 241707 249307 241712
rect 527406 241768 527515 241770
rect 527406 241712 527454 241768
rect 527510 241712 527515 241768
rect 527406 241707 527515 241712
rect 249198 241636 249258 241707
rect 527406 241636 527466 241707
rect 249190 241572 249196 241636
rect 249260 241572 249266 241636
rect 527398 241572 527404 241636
rect 527468 241572 527474 241636
rect 242985 241498 243051 241501
rect 243169 241498 243235 241501
rect 242985 241496 243235 241498
rect 242985 241440 242990 241496
rect 243046 241440 243174 241496
rect 243230 241440 243235 241496
rect 242985 241438 243235 241440
rect 242985 241435 243051 241438
rect 243169 241435 243235 241438
rect 254025 241498 254091 241501
rect 254209 241498 254275 241501
rect 254025 241496 254275 241498
rect 254025 241440 254030 241496
rect 254086 241440 254214 241496
rect 254270 241440 254275 241496
rect 254025 241438 254275 241440
rect 254025 241435 254091 241438
rect 254209 241435 254275 241438
rect 259545 241498 259611 241501
rect 259729 241498 259795 241501
rect 259545 241496 259795 241498
rect 259545 241440 259550 241496
rect 259606 241440 259734 241496
rect 259790 241440 259795 241496
rect 259545 241438 259795 241440
rect 259545 241435 259611 241438
rect 259729 241435 259795 241438
rect 282913 241498 282979 241501
rect 283097 241498 283163 241501
rect 282913 241496 283163 241498
rect 282913 241440 282918 241496
rect 282974 241440 283102 241496
rect 283158 241440 283163 241496
rect 282913 241438 283163 241440
rect 282913 241435 282979 241438
rect 283097 241435 283163 241438
rect 305177 241498 305243 241501
rect 305361 241498 305427 241501
rect 305177 241496 305427 241498
rect 305177 241440 305182 241496
rect 305238 241440 305366 241496
rect 305422 241440 305427 241496
rect 305177 241438 305427 241440
rect 305177 241435 305243 241438
rect 305361 241435 305427 241438
rect 310697 241498 310763 241501
rect 310881 241498 310947 241501
rect 310697 241496 310947 241498
rect 310697 241440 310702 241496
rect 310758 241440 310886 241496
rect 310942 241440 310947 241496
rect 310697 241438 310947 241440
rect 310697 241435 310763 241438
rect 310881 241435 310947 241438
rect 346577 241498 346643 241501
rect 346761 241498 346827 241501
rect 346577 241496 346827 241498
rect 346577 241440 346582 241496
rect 346638 241440 346766 241496
rect 346822 241440 346827 241496
rect 346577 241438 346827 241440
rect 346577 241435 346643 241438
rect 346761 241435 346827 241438
rect 376753 241498 376819 241501
rect 376937 241498 377003 241501
rect 376753 241496 377003 241498
rect 376753 241440 376758 241496
rect 376814 241440 376942 241496
rect 376998 241440 377003 241496
rect 376753 241438 377003 241440
rect 376753 241435 376819 241438
rect 376937 241435 377003 241438
rect 400305 241498 400371 241501
rect 400489 241498 400555 241501
rect 400305 241496 400555 241498
rect 400305 241440 400310 241496
rect 400366 241440 400494 241496
rect 400550 241440 400555 241496
rect 400305 241438 400555 241440
rect 400305 241435 400371 241438
rect 400489 241435 400555 241438
rect 416865 241498 416931 241501
rect 417141 241498 417207 241501
rect 416865 241496 417207 241498
rect 416865 241440 416870 241496
rect 416926 241440 417146 241496
rect 417202 241440 417207 241496
rect 416865 241438 417207 241440
rect 416865 241435 416931 241438
rect 417141 241435 417207 241438
rect 433425 241498 433491 241501
rect 433609 241498 433675 241501
rect 433425 241496 433675 241498
rect 433425 241440 433430 241496
rect 433486 241440 433614 241496
rect 433670 241440 433675 241496
rect 433425 241438 433675 241440
rect 433425 241435 433491 241438
rect 433609 241435 433675 241438
rect 472065 241498 472131 241501
rect 472341 241498 472407 241501
rect 472065 241496 472407 241498
rect 472065 241440 472070 241496
rect 472126 241440 472346 241496
rect 472402 241440 472407 241496
rect 472065 241438 472407 241440
rect 472065 241435 472131 241438
rect 472341 241435 472407 241438
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 2773 237010 2839 237013
rect -960 237008 2839 237010
rect -960 236952 2778 237008
rect 2834 236952 2839 237008
rect -960 236950 2839 236952
rect -960 236860 480 236950
rect 2773 236947 2839 236950
rect 527398 234636 527404 234700
rect 527468 234636 527474 234700
rect 527406 234426 527466 234636
rect 527582 234426 527588 234428
rect 527406 234366 527588 234426
rect 527582 234364 527588 234366
rect 527652 234364 527658 234428
rect 249190 231916 249196 231980
rect 249260 231978 249266 231980
rect 249374 231978 249380 231980
rect 249260 231918 249380 231978
rect 249260 231916 249266 231918
rect 249374 231916 249380 231918
rect 249444 231916 249450 231980
rect 230657 231842 230723 231845
rect 230841 231842 230907 231845
rect 230657 231840 230907 231842
rect 230657 231784 230662 231840
rect 230718 231784 230846 231840
rect 230902 231784 230907 231840
rect 230657 231782 230907 231784
rect 230657 231779 230723 231782
rect 230841 231779 230907 231782
rect 252737 231842 252803 231845
rect 252921 231842 252987 231845
rect 252737 231840 252987 231842
rect 252737 231784 252742 231840
rect 252798 231784 252926 231840
rect 252982 231784 252987 231840
rect 252737 231782 252987 231784
rect 252737 231779 252803 231782
rect 252921 231779 252987 231782
rect 287237 231842 287303 231845
rect 287421 231842 287487 231845
rect 287237 231840 287487 231842
rect 287237 231784 287242 231840
rect 287298 231784 287426 231840
rect 287482 231784 287487 231840
rect 287237 231782 287487 231784
rect 287237 231779 287303 231782
rect 287421 231779 287487 231782
rect 342437 231842 342503 231845
rect 342713 231842 342779 231845
rect 342437 231840 342779 231842
rect 342437 231784 342442 231840
rect 342498 231784 342718 231840
rect 342774 231784 342779 231840
rect 342437 231782 342779 231784
rect 342437 231779 342503 231782
rect 342713 231779 342779 231782
rect 375557 231842 375623 231845
rect 375833 231842 375899 231845
rect 375557 231840 375899 231842
rect 375557 231784 375562 231840
rect 375618 231784 375838 231840
rect 375894 231784 375899 231840
rect 375557 231782 375899 231784
rect 375557 231779 375623 231782
rect 375833 231779 375899 231782
rect 393221 231842 393287 231845
rect 393405 231842 393471 231845
rect 393221 231840 393471 231842
rect 393221 231784 393226 231840
rect 393282 231784 393410 231840
rect 393466 231784 393471 231840
rect 393221 231782 393471 231784
rect 393221 231779 393287 231782
rect 393405 231779 393471 231782
rect 451273 231842 451339 231845
rect 451457 231842 451523 231845
rect 527633 231844 527699 231845
rect 527582 231842 527588 231844
rect 451273 231840 451523 231842
rect 451273 231784 451278 231840
rect 451334 231784 451462 231840
rect 451518 231784 451523 231840
rect 451273 231782 451523 231784
rect 527542 231782 527588 231842
rect 527652 231840 527699 231844
rect 527694 231784 527699 231840
rect 451273 231779 451339 231782
rect 451457 231779 451523 231782
rect 527582 231780 527588 231782
rect 527652 231780 527699 231784
rect 527633 231779 527699 231780
rect 236269 230482 236335 230485
rect 236453 230482 236519 230485
rect 236269 230480 236519 230482
rect 236269 230424 236274 230480
rect 236330 230424 236458 230480
rect 236514 230424 236519 230480
rect 236269 230422 236519 230424
rect 236269 230419 236335 230422
rect 236453 230419 236519 230422
rect 265157 230482 265223 230485
rect 265341 230482 265407 230485
rect 265157 230480 265407 230482
rect 265157 230424 265162 230480
rect 265218 230424 265346 230480
rect 265402 230424 265407 230480
rect 265157 230422 265407 230424
rect 265157 230419 265223 230422
rect 265341 230419 265407 230422
rect 580717 228850 580783 228853
rect 583520 228850 584960 228940
rect 580717 228848 584960 228850
rect 580717 228792 580722 228848
rect 580778 228792 584960 228848
rect 580717 228790 584960 228792
rect 580717 228787 580783 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 4061 222594 4127 222597
rect -960 222592 4127 222594
rect -960 222536 4066 222592
rect 4122 222536 4127 222592
rect -960 222534 4127 222536
rect -960 222444 480 222534
rect 4061 222531 4127 222534
rect 249374 222260 249380 222324
rect 249444 222322 249450 222324
rect 527633 222322 527699 222325
rect 527766 222322 527772 222324
rect 249444 222262 249626 222322
rect 249444 222260 249450 222262
rect 249425 222186 249491 222189
rect 249566 222186 249626 222262
rect 527633 222320 527772 222322
rect 527633 222264 527638 222320
rect 527694 222264 527772 222320
rect 527633 222262 527772 222264
rect 527633 222259 527699 222262
rect 527766 222260 527772 222262
rect 527836 222260 527842 222324
rect 249425 222184 249626 222186
rect 249425 222128 249430 222184
rect 249486 222128 249626 222184
rect 249425 222126 249626 222128
rect 305177 222186 305243 222189
rect 305361 222186 305427 222189
rect 305177 222184 305427 222186
rect 305177 222128 305182 222184
rect 305238 222128 305366 222184
rect 305422 222128 305427 222184
rect 305177 222126 305427 222128
rect 249425 222123 249491 222126
rect 305177 222123 305243 222126
rect 305361 222123 305427 222126
rect 310697 222186 310763 222189
rect 310881 222186 310947 222189
rect 310697 222184 310947 222186
rect 310697 222128 310702 222184
rect 310758 222128 310886 222184
rect 310942 222128 310947 222184
rect 310697 222126 310947 222128
rect 310697 222123 310763 222126
rect 310881 222123 310947 222126
rect 346577 222186 346643 222189
rect 346761 222186 346827 222189
rect 346577 222184 346827 222186
rect 346577 222128 346582 222184
rect 346638 222128 346766 222184
rect 346822 222128 346827 222184
rect 346577 222126 346827 222128
rect 346577 222123 346643 222126
rect 346761 222123 346827 222126
rect 376753 222186 376819 222189
rect 376937 222186 377003 222189
rect 376753 222184 377003 222186
rect 376753 222128 376758 222184
rect 376814 222128 376942 222184
rect 376998 222128 377003 222184
rect 376753 222126 377003 222128
rect 376753 222123 376819 222126
rect 376937 222123 377003 222126
rect 400305 222186 400371 222189
rect 400489 222186 400555 222189
rect 400305 222184 400555 222186
rect 400305 222128 400310 222184
rect 400366 222128 400494 222184
rect 400550 222128 400555 222184
rect 400305 222126 400555 222128
rect 400305 222123 400371 222126
rect 400489 222123 400555 222126
rect 416865 222186 416931 222189
rect 417141 222186 417207 222189
rect 416865 222184 417207 222186
rect 416865 222128 416870 222184
rect 416926 222128 417146 222184
rect 417202 222128 417207 222184
rect 416865 222126 417207 222128
rect 416865 222123 416931 222126
rect 417141 222123 417207 222126
rect 433425 222186 433491 222189
rect 433609 222186 433675 222189
rect 433425 222184 433675 222186
rect 433425 222128 433430 222184
rect 433486 222128 433614 222184
rect 433670 222128 433675 222184
rect 433425 222126 433675 222128
rect 433425 222123 433491 222126
rect 433609 222123 433675 222126
rect 472065 222186 472131 222189
rect 472341 222186 472407 222189
rect 472065 222184 472407 222186
rect 472065 222128 472070 222184
rect 472126 222128 472346 222184
rect 472402 222128 472407 222184
rect 472065 222126 472407 222128
rect 472065 222123 472131 222126
rect 472341 222123 472407 222126
rect 231761 220826 231827 220829
rect 231945 220826 232011 220829
rect 231761 220824 232011 220826
rect 231761 220768 231766 220824
rect 231822 220768 231950 220824
rect 232006 220768 232011 220824
rect 231761 220766 232011 220768
rect 231761 220763 231827 220766
rect 231945 220763 232011 220766
rect 364425 217970 364491 217973
rect 364609 217970 364675 217973
rect 364425 217968 364675 217970
rect 364425 217912 364430 217968
rect 364486 217912 364614 217968
rect 364670 217912 364675 217968
rect 364425 217910 364675 217912
rect 364425 217907 364491 217910
rect 364609 217907 364675 217910
rect 579613 217018 579679 217021
rect 583520 217018 584960 217108
rect 579613 217016 584960 217018
rect 579613 216960 579618 217016
rect 579674 216960 584960 217016
rect 579613 216958 584960 216960
rect 579613 216955 579679 216958
rect 583520 216868 584960 216958
rect 527766 215522 527772 215524
rect 527590 215462 527772 215522
rect 527590 215252 527650 215462
rect 527766 215460 527772 215462
rect 527836 215460 527842 215524
rect 527582 215188 527588 215252
rect 527652 215188 527658 215252
rect 249425 214572 249491 214573
rect 249374 214570 249380 214572
rect 249334 214510 249380 214570
rect 249444 214568 249491 214572
rect 249486 214512 249491 214568
rect 249374 214508 249380 214510
rect 249444 214508 249491 214512
rect 249425 214507 249491 214508
rect 342713 212802 342779 212805
rect 342302 212800 342779 212802
rect 342302 212744 342718 212800
rect 342774 212744 342779 212800
rect 342302 212742 342779 212744
rect 342302 212564 342362 212742
rect 342713 212739 342779 212742
rect 342437 212564 342503 212567
rect 342302 212562 342503 212564
rect 230657 212530 230723 212533
rect 230841 212530 230907 212533
rect 230657 212528 230907 212530
rect 230657 212472 230662 212528
rect 230718 212472 230846 212528
rect 230902 212472 230907 212528
rect 230657 212470 230907 212472
rect 230657 212467 230723 212470
rect 230841 212467 230907 212470
rect 252461 212530 252527 212533
rect 252737 212530 252803 212533
rect 252461 212528 252803 212530
rect 252461 212472 252466 212528
rect 252522 212472 252742 212528
rect 252798 212472 252803 212528
rect 342302 212506 342442 212562
rect 342498 212506 342503 212562
rect 342302 212504 342503 212506
rect 342437 212501 342503 212504
rect 375557 212530 375623 212533
rect 375833 212530 375899 212533
rect 375557 212528 375899 212530
rect 252461 212470 252803 212472
rect 252461 212467 252527 212470
rect 252737 212467 252803 212470
rect 375557 212472 375562 212528
rect 375618 212472 375838 212528
rect 375894 212472 375899 212528
rect 375557 212470 375899 212472
rect 375557 212467 375623 212470
rect 375833 212467 375899 212470
rect 386597 212530 386663 212533
rect 386781 212530 386847 212533
rect 386597 212528 386847 212530
rect 386597 212472 386602 212528
rect 386658 212472 386786 212528
rect 386842 212472 386847 212528
rect 386597 212470 386847 212472
rect 386597 212467 386663 212470
rect 386781 212467 386847 212470
rect 392117 212530 392183 212533
rect 392301 212530 392367 212533
rect 392117 212528 392367 212530
rect 392117 212472 392122 212528
rect 392178 212472 392306 212528
rect 392362 212472 392367 212528
rect 392117 212470 392367 212472
rect 392117 212467 392183 212470
rect 392301 212467 392367 212470
rect 393221 212530 393287 212533
rect 393405 212530 393471 212533
rect 393221 212528 393471 212530
rect 393221 212472 393226 212528
rect 393282 212472 393410 212528
rect 393466 212472 393471 212528
rect 393221 212470 393471 212472
rect 393221 212467 393287 212470
rect 393405 212467 393471 212470
rect 397361 212530 397427 212533
rect 397545 212530 397611 212533
rect 397361 212528 397611 212530
rect 397361 212472 397366 212528
rect 397422 212472 397550 212528
rect 397606 212472 397611 212528
rect 397361 212470 397611 212472
rect 397361 212467 397427 212470
rect 397545 212467 397611 212470
rect 451273 212530 451339 212533
rect 451457 212530 451523 212533
rect 451273 212528 451523 212530
rect 451273 212472 451278 212528
rect 451334 212472 451462 212528
rect 451518 212472 451523 212528
rect 451273 212470 451523 212472
rect 451273 212467 451339 212470
rect 451457 212467 451523 212470
rect 527449 212530 527515 212533
rect 527582 212530 527588 212532
rect 527449 212528 527588 212530
rect 527449 212472 527454 212528
rect 527510 212472 527588 212528
rect 527449 212470 527588 212472
rect 527449 212467 527515 212470
rect 527582 212468 527588 212470
rect 527652 212468 527658 212532
rect 236269 211170 236335 211173
rect 236545 211170 236611 211173
rect 236269 211168 236611 211170
rect 236269 211112 236274 211168
rect 236330 211112 236550 211168
rect 236606 211112 236611 211168
rect 236269 211110 236611 211112
rect 236269 211107 236335 211110
rect 236545 211107 236611 211110
rect 281717 211170 281783 211173
rect 281901 211170 281967 211173
rect 281717 211168 281967 211170
rect 281717 211112 281722 211168
rect 281778 211112 281906 211168
rect 281962 211112 281967 211168
rect 281717 211110 281967 211112
rect 281717 211107 281783 211110
rect 281901 211107 281967 211110
rect 331121 209810 331187 209813
rect 331489 209810 331555 209813
rect 331121 209808 331555 209810
rect 331121 209752 331126 209808
rect 331182 209752 331494 209808
rect 331550 209752 331555 209808
rect 331121 209750 331555 209752
rect 331121 209747 331187 209750
rect 331489 209747 331555 209750
rect 232630 208314 232636 208316
rect -960 208178 480 208268
rect 614 208254 232636 208314
rect 614 208178 674 208254
rect 232630 208252 232636 208254
rect 232700 208252 232706 208316
rect -960 208118 674 208178
rect -960 208028 480 208118
rect 580165 205322 580231 205325
rect 583520 205322 584960 205412
rect 580165 205320 584960 205322
rect 580165 205264 580170 205320
rect 580226 205264 584960 205320
rect 580165 205262 584960 205264
rect 580165 205259 580231 205262
rect 583520 205172 584960 205262
rect 270585 203146 270651 203149
rect 527449 203146 527515 203149
rect 270585 203144 270970 203146
rect 270585 203088 270590 203144
rect 270646 203088 270970 203144
rect 270585 203086 270970 203088
rect 270585 203083 270651 203086
rect 270769 203010 270835 203013
rect 270910 203010 270970 203086
rect 527406 203144 527515 203146
rect 527406 203088 527454 203144
rect 527510 203088 527515 203144
rect 527406 203083 527515 203088
rect 527406 203012 527466 203083
rect 270769 203008 270970 203010
rect 270769 202952 270774 203008
rect 270830 202952 270970 203008
rect 270769 202950 270970 202952
rect 270769 202947 270835 202950
rect 527398 202948 527404 203012
rect 527468 202948 527474 203012
rect 266353 202874 266419 202877
rect 266537 202874 266603 202877
rect 266353 202872 266603 202874
rect 266353 202816 266358 202872
rect 266414 202816 266542 202872
rect 266598 202816 266603 202872
rect 266353 202814 266603 202816
rect 266353 202811 266419 202814
rect 266537 202811 266603 202814
rect 305177 202874 305243 202877
rect 305361 202874 305427 202877
rect 305177 202872 305427 202874
rect 305177 202816 305182 202872
rect 305238 202816 305366 202872
rect 305422 202816 305427 202872
rect 305177 202814 305427 202816
rect 305177 202811 305243 202814
rect 305361 202811 305427 202814
rect 310697 202874 310763 202877
rect 310881 202874 310947 202877
rect 310697 202872 310947 202874
rect 310697 202816 310702 202872
rect 310758 202816 310886 202872
rect 310942 202816 310947 202872
rect 310697 202814 310947 202816
rect 310697 202811 310763 202814
rect 310881 202811 310947 202814
rect 346577 202874 346643 202877
rect 346761 202874 346827 202877
rect 346577 202872 346827 202874
rect 346577 202816 346582 202872
rect 346638 202816 346766 202872
rect 346822 202816 346827 202872
rect 346577 202814 346827 202816
rect 346577 202811 346643 202814
rect 346761 202811 346827 202814
rect 352005 202874 352071 202877
rect 376753 202874 376819 202877
rect 376937 202874 377003 202877
rect 352005 202872 352114 202874
rect 352005 202816 352010 202872
rect 352066 202816 352114 202872
rect 352005 202811 352114 202816
rect 376753 202872 377003 202874
rect 376753 202816 376758 202872
rect 376814 202816 376942 202872
rect 376998 202816 377003 202872
rect 376753 202814 377003 202816
rect 376753 202811 376819 202814
rect 376937 202811 377003 202814
rect 400305 202874 400371 202877
rect 400489 202874 400555 202877
rect 400305 202872 400555 202874
rect 400305 202816 400310 202872
rect 400366 202816 400494 202872
rect 400550 202816 400555 202872
rect 400305 202814 400555 202816
rect 400305 202811 400371 202814
rect 400489 202811 400555 202814
rect 416865 202874 416931 202877
rect 417141 202874 417207 202877
rect 416865 202872 417207 202874
rect 416865 202816 416870 202872
rect 416926 202816 417146 202872
rect 417202 202816 417207 202872
rect 416865 202814 417207 202816
rect 416865 202811 416931 202814
rect 417141 202811 417207 202814
rect 433425 202874 433491 202877
rect 433609 202874 433675 202877
rect 433425 202872 433675 202874
rect 433425 202816 433430 202872
rect 433486 202816 433614 202872
rect 433670 202816 433675 202872
rect 433425 202814 433675 202816
rect 433425 202811 433491 202814
rect 433609 202811 433675 202814
rect 472065 202874 472131 202877
rect 472341 202874 472407 202877
rect 472065 202872 472407 202874
rect 472065 202816 472070 202872
rect 472126 202816 472346 202872
rect 472402 202816 472407 202872
rect 472065 202814 472407 202816
rect 472065 202811 472131 202814
rect 472341 202811 472407 202814
rect 352054 202741 352114 202811
rect 352054 202736 352163 202741
rect 352054 202680 352102 202736
rect 352158 202680 352163 202736
rect 352054 202678 352163 202680
rect 352097 202675 352163 202678
rect 294137 201650 294203 201653
rect 294137 201648 294338 201650
rect 294137 201592 294142 201648
rect 294198 201592 294338 201648
rect 294137 201590 294338 201592
rect 294137 201587 294203 201590
rect 294137 201514 294203 201517
rect 294278 201514 294338 201590
rect 294137 201512 294338 201514
rect 294137 201456 294142 201512
rect 294198 201456 294338 201512
rect 294137 201454 294338 201456
rect 370037 201514 370103 201517
rect 370221 201514 370287 201517
rect 370037 201512 370287 201514
rect 370037 201456 370042 201512
rect 370098 201456 370226 201512
rect 370282 201456 370287 201512
rect 370037 201454 370287 201456
rect 294137 201451 294203 201454
rect 370037 201451 370103 201454
rect 370221 201451 370287 201454
rect 358905 200154 358971 200157
rect 359089 200154 359155 200157
rect 358905 200152 359155 200154
rect 358905 200096 358910 200152
rect 358966 200096 359094 200152
rect 359150 200096 359155 200152
rect 358905 200094 359155 200096
rect 358905 200091 358971 200094
rect 359089 200091 359155 200094
rect 364425 200154 364491 200157
rect 364609 200154 364675 200157
rect 364425 200152 364675 200154
rect 364425 200096 364430 200152
rect 364486 200096 364614 200152
rect 364670 200096 364675 200152
rect 364425 200094 364675 200096
rect 364425 200091 364491 200094
rect 364609 200091 364675 200094
rect 249558 199956 249564 200020
rect 249628 199956 249634 200020
rect 249566 199885 249626 199956
rect 249517 199880 249626 199885
rect 249517 199824 249522 199880
rect 249578 199824 249626 199880
rect 249517 199822 249626 199824
rect 249517 199819 249583 199822
rect 527398 196012 527404 196076
rect 527468 196012 527474 196076
rect 527406 195802 527466 196012
rect 527582 195802 527588 195804
rect 527406 195742 527588 195802
rect 527582 195740 527588 195742
rect 527652 195740 527658 195804
rect -960 193898 480 193988
rect 3141 193898 3207 193901
rect -960 193896 3207 193898
rect -960 193840 3146 193896
rect 3202 193840 3207 193896
rect -960 193838 3207 193840
rect -960 193748 480 193838
rect 3141 193835 3207 193838
rect 583520 193476 584960 193716
rect 230657 193218 230723 193221
rect 230841 193218 230907 193221
rect 230657 193216 230907 193218
rect 230657 193160 230662 193216
rect 230718 193160 230846 193216
rect 230902 193160 230907 193216
rect 230657 193158 230907 193160
rect 230657 193155 230723 193158
rect 230841 193155 230907 193158
rect 254117 193218 254183 193221
rect 254301 193218 254367 193221
rect 254117 193216 254367 193218
rect 254117 193160 254122 193216
rect 254178 193160 254306 193216
rect 254362 193160 254367 193216
rect 254117 193158 254367 193160
rect 254117 193155 254183 193158
rect 254301 193155 254367 193158
rect 287237 193218 287303 193221
rect 287421 193218 287487 193221
rect 287237 193216 287487 193218
rect 287237 193160 287242 193216
rect 287298 193160 287426 193216
rect 287482 193160 287487 193216
rect 287237 193158 287487 193160
rect 287237 193155 287303 193158
rect 287421 193155 287487 193158
rect 347957 193218 348023 193221
rect 348141 193218 348207 193221
rect 347957 193216 348207 193218
rect 347957 193160 347962 193216
rect 348018 193160 348146 193216
rect 348202 193160 348207 193216
rect 347957 193158 348207 193160
rect 347957 193155 348023 193158
rect 348141 193155 348207 193158
rect 353477 193218 353543 193221
rect 353661 193218 353727 193221
rect 353477 193216 353727 193218
rect 353477 193160 353482 193216
rect 353538 193160 353666 193216
rect 353722 193160 353727 193216
rect 353477 193158 353727 193160
rect 353477 193155 353543 193158
rect 353661 193155 353727 193158
rect 386597 193218 386663 193221
rect 386781 193218 386847 193221
rect 386597 193216 386847 193218
rect 386597 193160 386602 193216
rect 386658 193160 386786 193216
rect 386842 193160 386847 193216
rect 386597 193158 386847 193160
rect 386597 193155 386663 193158
rect 386781 193155 386847 193158
rect 393221 193218 393287 193221
rect 393405 193218 393471 193221
rect 393221 193216 393471 193218
rect 393221 193160 393226 193216
rect 393282 193160 393410 193216
rect 393466 193160 393471 193216
rect 393221 193158 393471 193160
rect 393221 193155 393287 193158
rect 393405 193155 393471 193158
rect 397545 193218 397611 193221
rect 397729 193218 397795 193221
rect 397545 193216 397795 193218
rect 397545 193160 397550 193216
rect 397606 193160 397734 193216
rect 397790 193160 397795 193216
rect 397545 193158 397795 193160
rect 397545 193155 397611 193158
rect 397729 193155 397795 193158
rect 408677 193218 408743 193221
rect 408953 193218 409019 193221
rect 408677 193216 409019 193218
rect 408677 193160 408682 193216
rect 408738 193160 408958 193216
rect 409014 193160 409019 193216
rect 408677 193158 409019 193160
rect 408677 193155 408743 193158
rect 408953 193155 409019 193158
rect 527449 193218 527515 193221
rect 527582 193218 527588 193220
rect 527449 193216 527588 193218
rect 527449 193160 527454 193216
rect 527510 193160 527588 193216
rect 527449 193158 527588 193160
rect 527449 193155 527515 193158
rect 527582 193156 527588 193158
rect 527652 193156 527658 193220
rect 375557 191994 375623 191997
rect 375422 191992 375623 191994
rect 375422 191936 375562 191992
rect 375618 191936 375623 191992
rect 375422 191934 375623 191936
rect 342713 191858 342779 191861
rect 342897 191858 342963 191861
rect 342713 191856 342963 191858
rect 342713 191800 342718 191856
rect 342774 191800 342902 191856
rect 342958 191800 342963 191856
rect 342713 191798 342963 191800
rect 375422 191858 375482 191934
rect 375557 191931 375623 191934
rect 375557 191858 375623 191861
rect 375422 191856 375623 191858
rect 375422 191800 375562 191856
rect 375618 191800 375623 191856
rect 375422 191798 375623 191800
rect 342713 191795 342779 191798
rect 342897 191795 342963 191798
rect 375557 191795 375623 191798
rect 295425 190498 295491 190501
rect 295609 190498 295675 190501
rect 295425 190496 295675 190498
rect 295425 190440 295430 190496
rect 295486 190440 295614 190496
rect 295670 190440 295675 190496
rect 295425 190438 295675 190440
rect 295425 190435 295491 190438
rect 295609 190435 295675 190438
rect 358905 190498 358971 190501
rect 359181 190498 359247 190501
rect 358905 190496 359247 190498
rect 358905 190440 358910 190496
rect 358966 190440 359186 190496
rect 359242 190440 359247 190496
rect 358905 190438 359247 190440
rect 358905 190435 358971 190438
rect 359181 190435 359247 190438
rect 364609 190498 364675 190501
rect 364793 190498 364859 190501
rect 364609 190496 364859 190498
rect 364609 190440 364614 190496
rect 364670 190440 364798 190496
rect 364854 190440 364859 190496
rect 364609 190438 364859 190440
rect 364609 190435 364675 190438
rect 364793 190435 364859 190438
rect 392025 190498 392091 190501
rect 392209 190498 392275 190501
rect 392025 190496 392275 190498
rect 392025 190440 392030 190496
rect 392086 190440 392214 190496
rect 392270 190440 392275 190496
rect 392025 190438 392275 190440
rect 392025 190435 392091 190438
rect 392209 190435 392275 190438
rect 249517 185604 249583 185605
rect 249517 185602 249564 185604
rect 249472 185600 249564 185602
rect 249472 185544 249522 185600
rect 249472 185542 249564 185544
rect 249517 185540 249564 185542
rect 249628 185540 249634 185604
rect 249517 185539 249583 185540
rect 309225 183834 309291 183837
rect 527449 183834 527515 183837
rect 309225 183832 309610 183834
rect 309225 183776 309230 183832
rect 309286 183776 309610 183832
rect 309225 183774 309610 183776
rect 309225 183771 309291 183774
rect 309409 183698 309475 183701
rect 309550 183698 309610 183774
rect 527406 183832 527515 183834
rect 527406 183776 527454 183832
rect 527510 183776 527515 183832
rect 527406 183771 527515 183776
rect 527406 183700 527466 183771
rect 309409 183696 309610 183698
rect 309409 183640 309414 183696
rect 309470 183640 309610 183696
rect 309409 183638 309610 183640
rect 309409 183635 309475 183638
rect 527398 183636 527404 183700
rect 527468 183636 527474 183700
rect 241789 183562 241855 183565
rect 241973 183562 242039 183565
rect 241789 183560 242039 183562
rect 241789 183504 241794 183560
rect 241850 183504 241978 183560
rect 242034 183504 242039 183560
rect 241789 183502 242039 183504
rect 241789 183499 241855 183502
rect 241973 183499 242039 183502
rect 266997 183562 267063 183565
rect 267181 183562 267247 183565
rect 271965 183562 272031 183565
rect 266997 183560 267247 183562
rect 266997 183504 267002 183560
rect 267058 183504 267186 183560
rect 267242 183504 267247 183560
rect 266997 183502 267247 183504
rect 266997 183499 267063 183502
rect 267181 183499 267247 183502
rect 271830 183560 272031 183562
rect 271830 183504 271970 183560
rect 272026 183504 272031 183560
rect 271830 183502 272031 183504
rect 271830 183426 271890 183502
rect 271965 183499 272031 183502
rect 282913 183562 282979 183565
rect 283097 183562 283163 183565
rect 282913 183560 283163 183562
rect 282913 183504 282918 183560
rect 282974 183504 283102 183560
rect 283158 183504 283163 183560
rect 282913 183502 283163 183504
rect 282913 183499 282979 183502
rect 283097 183499 283163 183502
rect 305177 183562 305243 183565
rect 305361 183562 305427 183565
rect 305177 183560 305427 183562
rect 305177 183504 305182 183560
rect 305238 183504 305366 183560
rect 305422 183504 305427 183560
rect 305177 183502 305427 183504
rect 305177 183499 305243 183502
rect 305361 183499 305427 183502
rect 308029 183562 308095 183565
rect 308305 183562 308371 183565
rect 308029 183560 308371 183562
rect 308029 183504 308034 183560
rect 308090 183504 308310 183560
rect 308366 183504 308371 183560
rect 308029 183502 308371 183504
rect 308029 183499 308095 183502
rect 308305 183499 308371 183502
rect 346577 183562 346643 183565
rect 346761 183562 346827 183565
rect 346577 183560 346827 183562
rect 346577 183504 346582 183560
rect 346638 183504 346766 183560
rect 346822 183504 346827 183560
rect 346577 183502 346827 183504
rect 346577 183499 346643 183502
rect 346761 183499 346827 183502
rect 376753 183562 376819 183565
rect 376937 183562 377003 183565
rect 376753 183560 377003 183562
rect 376753 183504 376758 183560
rect 376814 183504 376942 183560
rect 376998 183504 377003 183560
rect 376753 183502 377003 183504
rect 376753 183499 376819 183502
rect 376937 183499 377003 183502
rect 380801 183562 380867 183565
rect 381077 183562 381143 183565
rect 380801 183560 381143 183562
rect 380801 183504 380806 183560
rect 380862 183504 381082 183560
rect 381138 183504 381143 183560
rect 380801 183502 381143 183504
rect 380801 183499 380867 183502
rect 381077 183499 381143 183502
rect 416865 183562 416931 183565
rect 417141 183562 417207 183565
rect 416865 183560 417207 183562
rect 416865 183504 416870 183560
rect 416926 183504 417146 183560
rect 417202 183504 417207 183560
rect 416865 183502 417207 183504
rect 416865 183499 416931 183502
rect 417141 183499 417207 183502
rect 422385 183562 422451 183565
rect 422661 183562 422727 183565
rect 422385 183560 422727 183562
rect 422385 183504 422390 183560
rect 422446 183504 422666 183560
rect 422722 183504 422727 183560
rect 422385 183502 422727 183504
rect 422385 183499 422451 183502
rect 422661 183499 422727 183502
rect 472065 183562 472131 183565
rect 472341 183562 472407 183565
rect 472065 183560 472407 183562
rect 472065 183504 472070 183560
rect 472126 183504 472346 183560
rect 472402 183504 472407 183560
rect 472065 183502 472407 183504
rect 472065 183499 472131 183502
rect 472341 183499 472407 183502
rect 272241 183426 272307 183429
rect 271830 183424 272307 183426
rect 271830 183368 272246 183424
rect 272302 183368 272307 183424
rect 271830 183366 272307 183368
rect 272241 183363 272307 183366
rect 259637 182338 259703 182341
rect 259637 182336 259746 182338
rect 259637 182280 259642 182336
rect 259698 182280 259746 182336
rect 259637 182275 259746 182280
rect 259686 182205 259746 182275
rect 244457 182202 244523 182205
rect 244641 182202 244707 182205
rect 244457 182200 244707 182202
rect 244457 182144 244462 182200
rect 244518 182144 244646 182200
rect 244702 182144 244707 182200
rect 244457 182142 244707 182144
rect 259686 182200 259795 182205
rect 259686 182144 259734 182200
rect 259790 182144 259795 182200
rect 259686 182142 259795 182144
rect 244457 182139 244523 182142
rect 244641 182139 244707 182142
rect 259729 182139 259795 182142
rect 270401 182202 270467 182205
rect 270585 182202 270651 182205
rect 270401 182200 270651 182202
rect 270401 182144 270406 182200
rect 270462 182144 270590 182200
rect 270646 182144 270651 182200
rect 270401 182142 270651 182144
rect 270401 182139 270467 182142
rect 270585 182139 270651 182142
rect 324221 182202 324287 182205
rect 324497 182202 324563 182205
rect 324221 182200 324563 182202
rect 324221 182144 324226 182200
rect 324282 182144 324502 182200
rect 324558 182144 324563 182200
rect 324221 182142 324563 182144
rect 324221 182139 324287 182142
rect 324497 182139 324563 182142
rect 369761 182202 369827 182205
rect 369945 182202 370011 182205
rect 369761 182200 370011 182202
rect 369761 182144 369766 182200
rect 369822 182144 369950 182200
rect 370006 182144 370011 182200
rect 369761 182142 370011 182144
rect 369761 182139 369827 182142
rect 369945 182139 370011 182142
rect 375465 182202 375531 182205
rect 375741 182202 375807 182205
rect 375465 182200 375807 182202
rect 375465 182144 375470 182200
rect 375526 182144 375746 182200
rect 375802 182144 375807 182200
rect 375465 182142 375807 182144
rect 375465 182139 375531 182142
rect 375741 182139 375807 182142
rect 580625 181930 580691 181933
rect 583520 181930 584960 182020
rect 580625 181928 584960 181930
rect 580625 181872 580630 181928
rect 580686 181872 584960 181928
rect 580625 181870 584960 181872
rect 580625 181867 580691 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 2773 179482 2839 179485
rect -960 179480 2839 179482
rect -960 179424 2778 179480
rect 2834 179424 2839 179480
rect -960 179422 2839 179424
rect -960 179332 480 179422
rect 2773 179419 2839 179422
rect 249609 179348 249675 179349
rect 249558 179284 249564 179348
rect 249628 179346 249675 179348
rect 249628 179344 249720 179346
rect 249670 179288 249720 179344
rect 249628 179286 249720 179288
rect 249628 179284 249675 179286
rect 249609 179283 249675 179284
rect 527398 176762 527404 176764
rect 527222 176702 527404 176762
rect 527222 176492 527282 176702
rect 527398 176700 527404 176702
rect 527468 176700 527474 176764
rect 527214 176428 527220 176492
rect 527284 176428 527290 176492
rect 353477 173906 353543 173909
rect 356421 173906 356487 173909
rect 527265 173908 527331 173909
rect 527214 173906 527220 173908
rect 353477 173904 353586 173906
rect 353477 173848 353482 173904
rect 353538 173848 353586 173904
rect 353477 173843 353586 173848
rect 356421 173904 356530 173906
rect 356421 173848 356426 173904
rect 356482 173848 356530 173904
rect 356421 173843 356530 173848
rect 527174 173846 527220 173906
rect 527284 173904 527331 173908
rect 527326 173848 527331 173904
rect 527214 173844 527220 173846
rect 527284 173844 527331 173848
rect 527265 173843 527331 173844
rect 353526 173773 353586 173843
rect 356470 173773 356530 173843
rect 353526 173768 353635 173773
rect 353526 173712 353574 173768
rect 353630 173712 353635 173768
rect 353526 173710 353635 173712
rect 356470 173768 356579 173773
rect 356470 173712 356518 173768
rect 356574 173712 356579 173768
rect 356470 173710 356579 173712
rect 353569 173707 353635 173710
rect 356513 173707 356579 173710
rect 331489 172682 331555 172685
rect 331262 172680 331555 172682
rect 331262 172624 331494 172680
rect 331550 172624 331555 172680
rect 331262 172622 331555 172624
rect 259637 172546 259703 172549
rect 259913 172546 259979 172549
rect 259637 172544 259979 172546
rect 259637 172488 259642 172544
rect 259698 172488 259918 172544
rect 259974 172488 259979 172544
rect 259637 172486 259979 172488
rect 259637 172483 259703 172486
rect 259913 172483 259979 172486
rect 270677 172546 270743 172549
rect 270861 172546 270927 172549
rect 270677 172544 270927 172546
rect 270677 172488 270682 172544
rect 270738 172488 270866 172544
rect 270922 172488 270927 172544
rect 270677 172486 270927 172488
rect 331262 172546 331322 172622
rect 331489 172619 331555 172622
rect 331397 172546 331463 172549
rect 331262 172544 331463 172546
rect 331262 172488 331402 172544
rect 331458 172488 331463 172544
rect 331262 172486 331463 172488
rect 270677 172483 270743 172486
rect 270861 172483 270927 172486
rect 331397 172483 331463 172486
rect 342437 172546 342503 172549
rect 342713 172546 342779 172549
rect 342437 172544 342779 172546
rect 342437 172488 342442 172544
rect 342498 172488 342718 172544
rect 342774 172488 342779 172544
rect 342437 172486 342779 172488
rect 342437 172483 342503 172486
rect 342713 172483 342779 172486
rect 364517 172546 364583 172549
rect 364701 172546 364767 172549
rect 364517 172544 364767 172546
rect 364517 172488 364522 172544
rect 364578 172488 364706 172544
rect 364762 172488 364767 172544
rect 364517 172486 364767 172488
rect 364517 172483 364583 172486
rect 364701 172483 364767 172486
rect 370221 172546 370287 172549
rect 370405 172546 370471 172549
rect 370221 172544 370471 172546
rect 370221 172488 370226 172544
rect 370282 172488 370410 172544
rect 370466 172488 370471 172544
rect 370221 172486 370471 172488
rect 370221 172483 370287 172486
rect 370405 172483 370471 172486
rect 375557 172546 375623 172549
rect 375741 172546 375807 172549
rect 375557 172544 375807 172546
rect 375557 172488 375562 172544
rect 375618 172488 375746 172544
rect 375802 172488 375807 172544
rect 375557 172486 375807 172488
rect 375557 172483 375623 172486
rect 375741 172483 375807 172486
rect 397361 172546 397427 172549
rect 397545 172546 397611 172549
rect 397361 172544 397611 172546
rect 397361 172488 397366 172544
rect 397422 172488 397550 172544
rect 397606 172488 397611 172544
rect 397361 172486 397611 172488
rect 397361 172483 397427 172486
rect 397545 172483 397611 172486
rect 243169 171186 243235 171189
rect 243353 171186 243419 171189
rect 243169 171184 243419 171186
rect 243169 171128 243174 171184
rect 243230 171128 243358 171184
rect 243414 171128 243419 171184
rect 243169 171126 243419 171128
rect 243169 171123 243235 171126
rect 243353 171123 243419 171126
rect 324221 171186 324287 171189
rect 324405 171186 324471 171189
rect 324221 171184 324471 171186
rect 324221 171128 324226 171184
rect 324282 171128 324410 171184
rect 324466 171128 324471 171184
rect 324221 171126 324471 171128
rect 324221 171123 324287 171126
rect 324405 171123 324471 171126
rect 550582 170444 550588 170508
rect 550652 170506 550658 170508
rect 560201 170506 560267 170509
rect 550652 170504 560267 170506
rect 550652 170448 560206 170504
rect 560262 170448 560267 170504
rect 550652 170446 560267 170448
rect 550652 170444 550658 170446
rect 560201 170443 560267 170446
rect 233734 170308 233740 170372
rect 233804 170370 233810 170372
rect 238753 170370 238819 170373
rect 233804 170368 238819 170370
rect 233804 170312 238758 170368
rect 238814 170312 238819 170368
rect 233804 170310 238819 170312
rect 233804 170308 233810 170310
rect 238753 170307 238819 170310
rect 248638 170308 248644 170372
rect 248708 170370 248714 170372
rect 259361 170370 259427 170373
rect 248708 170368 259427 170370
rect 248708 170312 259366 170368
rect 259422 170312 259427 170368
rect 248708 170310 259427 170312
rect 248708 170308 248714 170310
rect 259361 170307 259427 170310
rect 376702 170308 376708 170372
rect 376772 170370 376778 170372
rect 386321 170370 386387 170373
rect 376772 170368 386387 170370
rect 376772 170312 386326 170368
rect 386382 170312 386387 170368
rect 376772 170310 386387 170312
rect 376772 170308 376778 170310
rect 386321 170307 386387 170310
rect 521653 170370 521719 170373
rect 521653 170368 531330 170370
rect 521653 170312 521658 170368
rect 521714 170312 531330 170368
rect 521653 170310 531330 170312
rect 521653 170307 521719 170310
rect 355961 170234 356027 170237
rect 367001 170234 367067 170237
rect 531270 170234 531330 170310
rect 540881 170234 540947 170237
rect 550582 170234 550588 170236
rect 311758 170174 317338 170234
rect 248321 170098 248387 170101
rect 248454 170098 248460 170100
rect 248321 170096 248460 170098
rect 248321 170040 248326 170096
rect 248382 170040 248460 170096
rect 248321 170038 248460 170040
rect 248321 170035 248387 170038
rect 248454 170036 248460 170038
rect 248524 170036 248530 170100
rect 292941 170098 293007 170101
rect 298185 170098 298251 170101
rect 292941 170096 298251 170098
rect 292941 170040 292946 170096
rect 293002 170040 298190 170096
rect 298246 170040 298251 170096
rect 292941 170038 298251 170040
rect 292941 170035 293007 170038
rect 298185 170035 298251 170038
rect 249609 169962 249675 169965
rect 249566 169960 249675 169962
rect 249566 169904 249614 169960
rect 249670 169904 249675 169960
rect 249566 169899 249675 169904
rect 259361 169962 259427 169965
rect 267733 169962 267799 169965
rect 259361 169960 267799 169962
rect 259361 169904 259366 169960
rect 259422 169904 267738 169960
rect 267794 169904 267799 169960
rect 259361 169902 267799 169904
rect 259361 169899 259427 169902
rect 267733 169899 267799 169902
rect 283465 169962 283531 169965
rect 289629 169962 289695 169965
rect 283465 169960 289695 169962
rect 283465 169904 283470 169960
rect 283526 169904 289634 169960
rect 289690 169904 289695 169960
rect 283465 169902 289695 169904
rect 283465 169899 283531 169902
rect 289629 169899 289695 169902
rect 298185 169962 298251 169965
rect 311758 169962 311818 170174
rect 317278 170098 317338 170174
rect 355961 170232 367067 170234
rect 355961 170176 355966 170232
rect 356022 170176 367006 170232
rect 367062 170176 367067 170232
rect 355961 170174 367067 170176
rect 355961 170171 356027 170174
rect 367001 170171 367067 170174
rect 456566 170174 463618 170234
rect 317505 170098 317571 170101
rect 317278 170096 317571 170098
rect 317278 170040 317510 170096
rect 317566 170040 317571 170096
rect 317278 170038 317571 170040
rect 317505 170035 317571 170038
rect 331305 170098 331371 170101
rect 338021 170098 338087 170101
rect 331305 170096 338087 170098
rect 331305 170040 331310 170096
rect 331366 170040 338026 170096
rect 338082 170040 338087 170096
rect 331305 170038 338087 170040
rect 331305 170035 331371 170038
rect 338021 170035 338087 170038
rect 371877 170098 371943 170101
rect 376702 170098 376708 170100
rect 371877 170096 376708 170098
rect 371877 170040 371882 170096
rect 371938 170040 376708 170096
rect 371877 170038 376708 170040
rect 371877 170035 371943 170038
rect 376702 170036 376708 170038
rect 376772 170036 376778 170100
rect 434529 170098 434595 170101
rect 389222 170038 398850 170098
rect 298185 169960 311818 169962
rect 298185 169904 298190 169960
rect 298246 169904 311818 169960
rect 298185 169902 311818 169904
rect 386321 169962 386387 169965
rect 389222 169962 389282 170038
rect 386321 169960 389282 169962
rect 386321 169904 386326 169960
rect 386382 169904 389282 169960
rect 386321 169902 389282 169904
rect 298185 169899 298251 169902
rect 386321 169899 386387 169902
rect 249566 169828 249626 169899
rect 249558 169764 249564 169828
rect 249628 169764 249634 169828
rect 278681 169826 278747 169829
rect 317505 169826 317571 169829
rect 326061 169826 326127 169829
rect 367001 169826 367067 169829
rect 371877 169826 371943 169829
rect 278681 169824 278882 169826
rect 278681 169768 278686 169824
rect 278742 169768 278882 169824
rect 278681 169766 278882 169768
rect 278681 169763 278747 169766
rect 278822 169554 278882 169766
rect 317505 169824 326127 169826
rect 317505 169768 317510 169824
rect 317566 169768 326066 169824
rect 326122 169768 326127 169824
rect 317505 169766 326127 169768
rect 317505 169763 317571 169766
rect 326061 169763 326127 169766
rect 338254 169766 346410 169826
rect 338021 169690 338087 169693
rect 338254 169690 338314 169766
rect 338021 169688 338314 169690
rect 338021 169632 338026 169688
rect 338082 169632 338314 169688
rect 338021 169630 338314 169632
rect 338021 169627 338087 169630
rect 283465 169554 283531 169557
rect 278822 169552 283531 169554
rect 278822 169496 283470 169552
rect 283526 169496 283531 169552
rect 278822 169494 283531 169496
rect 346350 169554 346410 169766
rect 367001 169824 371943 169826
rect 367001 169768 367006 169824
rect 367062 169768 371882 169824
rect 371938 169768 371943 169824
rect 367001 169766 371943 169768
rect 398790 169826 398850 170038
rect 434529 170096 437490 170098
rect 434529 170040 434534 170096
rect 434590 170040 437490 170096
rect 434529 170038 437490 170040
rect 434529 170035 434595 170038
rect 418061 169962 418127 169965
rect 408542 169960 418127 169962
rect 408542 169904 418066 169960
rect 418122 169904 418127 169960
rect 408542 169902 418127 169904
rect 408542 169826 408602 169902
rect 418061 169899 418127 169902
rect 425053 169826 425119 169829
rect 398790 169766 408602 169826
rect 424918 169824 425119 169826
rect 424918 169768 425058 169824
rect 425114 169768 425119 169824
rect 424918 169766 425119 169768
rect 437430 169826 437490 170038
rect 456566 169962 456626 170174
rect 447182 169902 456626 169962
rect 447182 169826 447242 169902
rect 437430 169766 447242 169826
rect 463558 169826 463618 170174
rect 495206 170174 502258 170234
rect 531270 170232 540947 170234
rect 531270 170176 540886 170232
rect 540942 170176 540947 170232
rect 531270 170174 540947 170176
rect 475929 169962 475995 169965
rect 466502 169960 475995 169962
rect 466502 169904 475934 169960
rect 475990 169904 475995 169960
rect 466502 169902 475995 169904
rect 466502 169826 466562 169902
rect 475929 169899 475995 169902
rect 478137 169962 478203 169965
rect 495206 169962 495266 170174
rect 478137 169960 482938 169962
rect 478137 169904 478142 169960
rect 478198 169904 482938 169960
rect 478137 169902 482938 169904
rect 478137 169899 478203 169902
rect 463558 169766 466562 169826
rect 482878 169826 482938 169902
rect 485822 169902 495266 169962
rect 485822 169826 485882 169902
rect 482878 169766 485882 169826
rect 502198 169826 502258 170174
rect 540881 170171 540947 170174
rect 543782 170174 550588 170234
rect 540881 169962 540947 169965
rect 543782 169962 543842 170174
rect 550582 170172 550588 170174
rect 550652 170172 550658 170236
rect 560201 170098 560267 170101
rect 583520 170098 584960 170188
rect 560201 170096 563162 170098
rect 560201 170040 560206 170096
rect 560262 170040 563162 170096
rect 560201 170038 563162 170040
rect 560201 170035 560267 170038
rect 505142 169902 521578 169962
rect 505142 169826 505202 169902
rect 502198 169766 505202 169826
rect 521518 169826 521578 169902
rect 540881 169960 543842 169962
rect 540881 169904 540886 169960
rect 540942 169904 543842 169960
rect 540881 169902 543842 169904
rect 540881 169899 540947 169902
rect 521653 169826 521719 169829
rect 521518 169824 521719 169826
rect 521518 169768 521658 169824
rect 521714 169768 521719 169824
rect 521518 169766 521719 169768
rect 563102 169826 563162 170038
rect 583342 170038 584960 170098
rect 572621 169962 572687 169965
rect 583342 169962 583402 170038
rect 569910 169960 572687 169962
rect 569910 169904 572626 169960
rect 572682 169904 572687 169960
rect 569910 169902 572687 169904
rect 569910 169826 569970 169902
rect 572621 169899 572687 169902
rect 576902 169902 583402 169962
rect 583520 169948 584960 170038
rect 563102 169766 569970 169826
rect 572713 169826 572779 169829
rect 576902 169826 576962 169902
rect 572713 169824 576962 169826
rect 572713 169768 572718 169824
rect 572774 169768 576962 169824
rect 572713 169766 576962 169768
rect 367001 169763 367067 169766
rect 371877 169763 371943 169766
rect 355961 169554 356027 169557
rect 346350 169552 356027 169554
rect 346350 169496 355966 169552
rect 356022 169496 356027 169552
rect 346350 169494 356027 169496
rect 283465 169491 283531 169494
rect 355961 169491 356027 169494
rect 418061 169554 418127 169557
rect 424918 169554 424978 169766
rect 425053 169763 425119 169766
rect 521653 169763 521719 169766
rect 572713 169763 572779 169766
rect 418061 169552 424978 169554
rect 418061 169496 418066 169552
rect 418122 169496 424978 169552
rect 418061 169494 424978 169496
rect 418061 169491 418127 169494
rect 249558 167044 249564 167108
rect 249628 167044 249634 167108
rect 249566 166972 249626 167044
rect 249558 166908 249564 166972
rect 249628 166908 249634 166972
rect 232446 165610 232452 165612
rect 614 165550 232452 165610
rect -960 165066 480 165156
rect 614 165066 674 165550
rect 232446 165548 232452 165550
rect 232516 165548 232522 165612
rect -960 165006 674 165066
rect -960 164916 480 165006
rect 265157 164386 265223 164389
rect 265157 164384 265266 164386
rect 265157 164328 265162 164384
rect 265218 164328 265266 164384
rect 265157 164323 265266 164328
rect 265206 164253 265266 164323
rect 240133 164250 240199 164253
rect 240317 164250 240383 164253
rect 240133 164248 240383 164250
rect 240133 164192 240138 164248
rect 240194 164192 240322 164248
rect 240378 164192 240383 164248
rect 240133 164190 240383 164192
rect 265206 164248 265315 164253
rect 265206 164192 265254 164248
rect 265310 164192 265315 164248
rect 265206 164190 265315 164192
rect 240133 164187 240199 164190
rect 240317 164187 240383 164190
rect 265249 164187 265315 164190
rect 272057 164250 272123 164253
rect 272241 164250 272307 164253
rect 352097 164250 352163 164253
rect 272057 164248 272307 164250
rect 272057 164192 272062 164248
rect 272118 164192 272246 164248
rect 272302 164192 272307 164248
rect 272057 164190 272307 164192
rect 272057 164187 272123 164190
rect 272241 164187 272307 164190
rect 351870 164248 352163 164250
rect 351870 164192 352102 164248
rect 352158 164192 352163 164248
rect 351870 164190 352163 164192
rect 351870 164114 351930 164190
rect 352097 164187 352163 164190
rect 370037 164250 370103 164253
rect 370221 164250 370287 164253
rect 370037 164248 370287 164250
rect 370037 164192 370042 164248
rect 370098 164192 370226 164248
rect 370282 164192 370287 164248
rect 370037 164190 370287 164192
rect 370037 164187 370103 164190
rect 370221 164187 370287 164190
rect 527265 164250 527331 164253
rect 527398 164250 527404 164252
rect 527265 164248 527404 164250
rect 527265 164192 527270 164248
rect 527326 164192 527404 164248
rect 527265 164190 527404 164192
rect 527265 164187 527331 164190
rect 527398 164188 527404 164190
rect 527468 164188 527474 164252
rect 352005 164114 352071 164117
rect 351870 164112 352071 164114
rect 351870 164056 352010 164112
rect 352066 164056 352071 164112
rect 351870 164054 352071 164056
rect 352005 164051 352071 164054
rect 579705 158402 579771 158405
rect 583520 158402 584960 158492
rect 579705 158400 584960 158402
rect 579705 158344 579710 158400
rect 579766 158344 584960 158400
rect 579705 158342 584960 158344
rect 579705 158339 579771 158342
rect 583520 158252 584960 158342
rect 370037 157588 370103 157589
rect 370037 157584 370084 157588
rect 370148 157586 370154 157588
rect 370037 157528 370042 157584
rect 370037 157524 370084 157528
rect 370148 157526 370194 157586
rect 370148 157524 370154 157526
rect 370037 157523 370103 157524
rect 527398 157450 527404 157452
rect 527222 157390 527404 157450
rect 527222 157180 527282 157390
rect 527398 157388 527404 157390
rect 527468 157388 527474 157452
rect 527214 157116 527220 157180
rect 527284 157116 527290 157180
rect 270861 154730 270927 154733
rect 342345 154730 342411 154733
rect 270542 154728 270927 154730
rect 270542 154672 270866 154728
rect 270922 154672 270927 154728
rect 270542 154670 270927 154672
rect 230657 154594 230723 154597
rect 230841 154594 230907 154597
rect 230657 154592 230907 154594
rect 230657 154536 230662 154592
rect 230718 154536 230846 154592
rect 230902 154536 230907 154592
rect 230657 154534 230907 154536
rect 230657 154531 230723 154534
rect 230841 154531 230907 154534
rect 249742 154532 249748 154596
rect 249812 154532 249818 154596
rect 252553 154594 252619 154597
rect 252737 154594 252803 154597
rect 254301 154594 254367 154597
rect 252553 154592 252803 154594
rect 252553 154536 252558 154592
rect 252614 154536 252742 154592
rect 252798 154536 252803 154592
rect 252553 154534 252803 154536
rect 249750 154460 249810 154532
rect 252553 154531 252619 154534
rect 252737 154531 252803 154534
rect 254166 154592 254367 154594
rect 254166 154536 254306 154592
rect 254362 154536 254367 154592
rect 254166 154534 254367 154536
rect 270542 154594 270602 154670
rect 270861 154667 270927 154670
rect 342302 154728 342411 154730
rect 342302 154672 342350 154728
rect 342406 154672 342411 154728
rect 342302 154667 342411 154672
rect 400305 154730 400371 154733
rect 400305 154728 400690 154730
rect 400305 154672 400310 154728
rect 400366 154672 400690 154728
rect 400305 154670 400690 154672
rect 400305 154667 400371 154670
rect 270677 154594 270743 154597
rect 270542 154592 270743 154594
rect 270542 154536 270682 154592
rect 270738 154536 270743 154592
rect 270542 154534 270743 154536
rect 249742 154396 249748 154460
rect 249812 154396 249818 154460
rect 254166 154458 254226 154534
rect 254301 154531 254367 154534
rect 270677 154531 270743 154534
rect 272057 154594 272123 154597
rect 272241 154594 272307 154597
rect 272057 154592 272307 154594
rect 272057 154536 272062 154592
rect 272118 154536 272246 154592
rect 272302 154536 272307 154592
rect 272057 154534 272307 154536
rect 272057 154531 272123 154534
rect 272241 154531 272307 154534
rect 277393 154594 277459 154597
rect 277669 154594 277735 154597
rect 277393 154592 277735 154594
rect 277393 154536 277398 154592
rect 277454 154536 277674 154592
rect 277730 154536 277735 154592
rect 277393 154534 277735 154536
rect 277393 154531 277459 154534
rect 277669 154531 277735 154534
rect 287237 154594 287303 154597
rect 287421 154594 287487 154597
rect 287237 154592 287487 154594
rect 287237 154536 287242 154592
rect 287298 154536 287426 154592
rect 287482 154536 287487 154592
rect 287237 154534 287487 154536
rect 287237 154531 287303 154534
rect 287421 154531 287487 154534
rect 308029 154594 308095 154597
rect 308305 154594 308371 154597
rect 308029 154592 308371 154594
rect 308029 154536 308034 154592
rect 308090 154536 308310 154592
rect 308366 154536 308371 154592
rect 308029 154534 308371 154536
rect 308029 154531 308095 154534
rect 308305 154531 308371 154534
rect 310697 154594 310763 154597
rect 310881 154594 310947 154597
rect 310697 154592 310947 154594
rect 310697 154536 310702 154592
rect 310758 154536 310886 154592
rect 310942 154536 310947 154592
rect 310697 154534 310947 154536
rect 342302 154594 342362 154667
rect 342437 154594 342503 154597
rect 342302 154592 342503 154594
rect 342302 154536 342442 154592
rect 342498 154536 342503 154592
rect 342302 154534 342503 154536
rect 310697 154531 310763 154534
rect 310881 154531 310947 154534
rect 342437 154531 342503 154534
rect 346577 154594 346643 154597
rect 346761 154594 346827 154597
rect 370037 154596 370103 154597
rect 370037 154594 370084 154596
rect 346577 154592 346827 154594
rect 346577 154536 346582 154592
rect 346638 154536 346766 154592
rect 346822 154536 346827 154592
rect 346577 154534 346827 154536
rect 369992 154592 370084 154594
rect 369992 154536 370042 154592
rect 369992 154534 370084 154536
rect 346577 154531 346643 154534
rect 346761 154531 346827 154534
rect 370037 154532 370084 154534
rect 370148 154532 370154 154596
rect 375189 154594 375255 154597
rect 375557 154594 375623 154597
rect 375189 154592 375623 154594
rect 375189 154536 375194 154592
rect 375250 154536 375562 154592
rect 375618 154536 375623 154592
rect 375189 154534 375623 154536
rect 370037 154531 370103 154532
rect 375189 154531 375255 154534
rect 375557 154531 375623 154534
rect 376753 154594 376819 154597
rect 376937 154594 377003 154597
rect 376753 154592 377003 154594
rect 376753 154536 376758 154592
rect 376814 154536 376942 154592
rect 376998 154536 377003 154592
rect 376753 154534 377003 154536
rect 376753 154531 376819 154534
rect 376937 154531 377003 154534
rect 400489 154594 400555 154597
rect 400630 154594 400690 154670
rect 400489 154592 400690 154594
rect 400489 154536 400494 154592
rect 400550 154536 400690 154592
rect 400489 154534 400690 154536
rect 416957 154594 417023 154597
rect 417141 154594 417207 154597
rect 416957 154592 417207 154594
rect 416957 154536 416962 154592
rect 417018 154536 417146 154592
rect 417202 154536 417207 154592
rect 416957 154534 417207 154536
rect 400489 154531 400555 154534
rect 416957 154531 417023 154534
rect 417141 154531 417207 154534
rect 433241 154594 433307 154597
rect 433701 154594 433767 154597
rect 433241 154592 433767 154594
rect 433241 154536 433246 154592
rect 433302 154536 433706 154592
rect 433762 154536 433767 154592
rect 433241 154534 433767 154536
rect 433241 154531 433307 154534
rect 433701 154531 433767 154534
rect 472157 154594 472223 154597
rect 472341 154594 472407 154597
rect 472157 154592 472407 154594
rect 472157 154536 472162 154592
rect 472218 154536 472346 154592
rect 472402 154536 472407 154592
rect 472157 154534 472407 154536
rect 472157 154531 472223 154534
rect 472341 154531 472407 154534
rect 254301 154458 254367 154461
rect 254166 154456 254367 154458
rect 254166 154400 254306 154456
rect 254362 154400 254367 154456
rect 254166 154398 254367 154400
rect 254301 154395 254367 154398
rect 527214 154396 527220 154460
rect 527284 154396 527290 154460
rect 527222 154325 527282 154396
rect 527222 154320 527331 154325
rect 527222 154264 527270 154320
rect 527326 154264 527331 154320
rect 527222 154262 527331 154264
rect 527265 154259 527331 154262
rect -960 150786 480 150876
rect 3969 150786 4035 150789
rect -960 150784 4035 150786
rect -960 150728 3974 150784
rect 4030 150728 4035 150784
rect -960 150726 4035 150728
rect -960 150636 480 150726
rect 3969 150723 4035 150726
rect 583520 146556 584960 146796
rect 230749 144938 230815 144941
rect 231025 144938 231091 144941
rect 230749 144936 231091 144938
rect 230749 144880 230754 144936
rect 230810 144880 231030 144936
rect 231086 144880 231091 144936
rect 230749 144878 231091 144880
rect 230749 144875 230815 144878
rect 231025 144875 231091 144878
rect 249374 144876 249380 144940
rect 249444 144938 249450 144940
rect 249742 144938 249748 144940
rect 249444 144878 249748 144938
rect 249444 144876 249450 144878
rect 249742 144876 249748 144878
rect 249812 144876 249818 144940
rect 271781 144938 271847 144941
rect 271965 144938 272031 144941
rect 271781 144936 272031 144938
rect 271781 144880 271786 144936
rect 271842 144880 271970 144936
rect 272026 144880 272031 144936
rect 271781 144878 272031 144880
rect 271781 144875 271847 144878
rect 271965 144875 272031 144878
rect 342345 144938 342411 144941
rect 342529 144938 342595 144941
rect 342345 144936 342595 144938
rect 342345 144880 342350 144936
rect 342406 144880 342534 144936
rect 342590 144880 342595 144936
rect 342345 144878 342595 144880
rect 342345 144875 342411 144878
rect 342529 144875 342595 144878
rect 351821 144938 351887 144941
rect 352005 144938 352071 144941
rect 351821 144936 352071 144938
rect 351821 144880 351826 144936
rect 351882 144880 352010 144936
rect 352066 144880 352071 144936
rect 351821 144878 352071 144880
rect 351821 144875 351887 144878
rect 352005 144875 352071 144878
rect 393221 144938 393287 144941
rect 393405 144938 393471 144941
rect 393221 144936 393471 144938
rect 393221 144880 393226 144936
rect 393282 144880 393410 144936
rect 393466 144880 393471 144936
rect 393221 144878 393471 144880
rect 393221 144875 393287 144878
rect 393405 144875 393471 144878
rect 527265 144938 527331 144941
rect 527398 144938 527404 144940
rect 527265 144936 527404 144938
rect 527265 144880 527270 144936
rect 527326 144880 527404 144936
rect 527265 144878 527404 144880
rect 527265 144875 527331 144878
rect 527398 144876 527404 144878
rect 527468 144876 527474 144940
rect 240133 143714 240199 143717
rect 240133 143712 240242 143714
rect 240133 143656 240138 143712
rect 240194 143656 240242 143712
rect 240133 143651 240242 143656
rect 240182 143581 240242 143651
rect 231945 143578 232011 143581
rect 232221 143578 232287 143581
rect 231945 143576 232287 143578
rect 231945 143520 231950 143576
rect 232006 143520 232226 143576
rect 232282 143520 232287 143576
rect 231945 143518 232287 143520
rect 231945 143515 232011 143518
rect 232221 143515 232287 143518
rect 240133 143576 240242 143581
rect 265249 143578 265315 143581
rect 240133 143520 240138 143576
rect 240194 143520 240242 143576
rect 240133 143518 240242 143520
rect 265206 143576 265315 143578
rect 265206 143520 265254 143576
rect 265310 143520 265315 143576
rect 240133 143515 240199 143518
rect 265206 143515 265315 143520
rect 281625 143578 281691 143581
rect 281809 143578 281875 143581
rect 281625 143576 281875 143578
rect 281625 143520 281630 143576
rect 281686 143520 281814 143576
rect 281870 143520 281875 143576
rect 281625 143518 281875 143520
rect 281625 143515 281691 143518
rect 281809 143515 281875 143518
rect 265206 143442 265266 143515
rect 265433 143442 265499 143445
rect 265206 143440 265499 143442
rect 265206 143384 265438 143440
rect 265494 143384 265499 143440
rect 265206 143382 265499 143384
rect 265433 143379 265499 143382
rect 527398 139980 527404 140044
rect 527468 140042 527474 140044
rect 527766 140042 527772 140044
rect 527468 139982 527772 140042
rect 527468 139980 527474 139982
rect 527766 139980 527772 139982
rect 527836 139980 527842 140044
rect 370129 138276 370195 138277
rect 370078 138274 370084 138276
rect 370038 138214 370084 138274
rect 370148 138272 370195 138276
rect 370190 138216 370195 138272
rect 370078 138212 370084 138214
rect 370148 138212 370195 138216
rect 370129 138211 370195 138212
rect -960 136370 480 136460
rect 3877 136370 3943 136373
rect -960 136368 3943 136370
rect -960 136312 3882 136368
rect 3938 136312 3943 136368
rect -960 136310 3943 136312
rect -960 136220 480 136310
rect 3877 136307 3943 136310
rect 375741 135418 375807 135421
rect 375422 135416 375807 135418
rect 375422 135360 375746 135416
rect 375802 135360 375807 135416
rect 375422 135358 375807 135360
rect 252553 135282 252619 135285
rect 252737 135282 252803 135285
rect 252553 135280 252803 135282
rect 252553 135224 252558 135280
rect 252614 135224 252742 135280
rect 252798 135224 252803 135280
rect 252553 135222 252803 135224
rect 252553 135219 252619 135222
rect 252737 135219 252803 135222
rect 254117 135282 254183 135285
rect 254301 135282 254367 135285
rect 254117 135280 254367 135282
rect 254117 135224 254122 135280
rect 254178 135224 254306 135280
rect 254362 135224 254367 135280
rect 254117 135222 254367 135224
rect 254117 135219 254183 135222
rect 254301 135219 254367 135222
rect 259637 135282 259703 135285
rect 259821 135282 259887 135285
rect 259637 135280 259887 135282
rect 259637 135224 259642 135280
rect 259698 135224 259826 135280
rect 259882 135224 259887 135280
rect 259637 135222 259887 135224
rect 259637 135219 259703 135222
rect 259821 135219 259887 135222
rect 270677 135282 270743 135285
rect 270861 135282 270927 135285
rect 270677 135280 270927 135282
rect 270677 135224 270682 135280
rect 270738 135224 270866 135280
rect 270922 135224 270927 135280
rect 270677 135222 270927 135224
rect 270677 135219 270743 135222
rect 270861 135219 270927 135222
rect 308121 135282 308187 135285
rect 308305 135282 308371 135285
rect 308121 135280 308371 135282
rect 308121 135224 308126 135280
rect 308182 135224 308310 135280
rect 308366 135224 308371 135280
rect 308121 135222 308371 135224
rect 308121 135219 308187 135222
rect 308305 135219 308371 135222
rect 310697 135282 310763 135285
rect 310881 135282 310947 135285
rect 330201 135282 330267 135285
rect 310697 135280 310947 135282
rect 310697 135224 310702 135280
rect 310758 135224 310886 135280
rect 310942 135224 310947 135280
rect 310697 135222 310947 135224
rect 310697 135219 310763 135222
rect 310881 135219 310947 135222
rect 329974 135280 330267 135282
rect 329974 135224 330206 135280
rect 330262 135224 330267 135280
rect 329974 135222 330267 135224
rect 329974 135149 330034 135222
rect 330201 135219 330267 135222
rect 346577 135282 346643 135285
rect 346761 135282 346827 135285
rect 346577 135280 346827 135282
rect 346577 135224 346582 135280
rect 346638 135224 346766 135280
rect 346822 135224 346827 135280
rect 346577 135222 346827 135224
rect 346577 135219 346643 135222
rect 346761 135219 346827 135222
rect 356421 135282 356487 135285
rect 356605 135282 356671 135285
rect 356421 135280 356671 135282
rect 356421 135224 356426 135280
rect 356482 135224 356610 135280
rect 356666 135224 356671 135280
rect 356421 135222 356671 135224
rect 356421 135219 356487 135222
rect 356605 135219 356671 135222
rect 364517 135282 364583 135285
rect 364701 135282 364767 135285
rect 370037 135284 370103 135285
rect 370037 135282 370084 135284
rect 364517 135280 364767 135282
rect 364517 135224 364522 135280
rect 364578 135224 364706 135280
rect 364762 135224 364767 135280
rect 364517 135222 364767 135224
rect 369992 135280 370084 135282
rect 369992 135224 370042 135280
rect 369992 135222 370084 135224
rect 364517 135219 364583 135222
rect 364701 135219 364767 135222
rect 370037 135220 370084 135222
rect 370148 135220 370154 135284
rect 375422 135282 375482 135358
rect 375741 135355 375807 135358
rect 375557 135282 375623 135285
rect 375422 135280 375623 135282
rect 375422 135224 375562 135280
rect 375618 135224 375623 135280
rect 375422 135222 375623 135224
rect 370037 135219 370103 135220
rect 375557 135219 375623 135222
rect 376753 135282 376819 135285
rect 376937 135282 377003 135285
rect 376753 135280 377003 135282
rect 376753 135224 376758 135280
rect 376814 135224 376942 135280
rect 376998 135224 377003 135280
rect 376753 135222 377003 135224
rect 376753 135219 376819 135222
rect 376937 135219 377003 135222
rect 386597 135282 386663 135285
rect 386781 135282 386847 135285
rect 386597 135280 386847 135282
rect 386597 135224 386602 135280
rect 386658 135224 386786 135280
rect 386842 135224 386847 135280
rect 386597 135222 386847 135224
rect 386597 135219 386663 135222
rect 386781 135219 386847 135222
rect 416773 135282 416839 135285
rect 416957 135282 417023 135285
rect 416773 135280 417023 135282
rect 416773 135224 416778 135280
rect 416834 135224 416962 135280
rect 417018 135224 417023 135280
rect 416773 135222 417023 135224
rect 416773 135219 416839 135222
rect 416957 135219 417023 135222
rect 433609 135282 433675 135285
rect 433793 135282 433859 135285
rect 433609 135280 433859 135282
rect 433609 135224 433614 135280
rect 433670 135224 433798 135280
rect 433854 135224 433859 135280
rect 433609 135222 433859 135224
rect 433609 135219 433675 135222
rect 433793 135219 433859 135222
rect 329925 135144 330034 135149
rect 527817 135148 527883 135149
rect 329925 135088 329930 135144
rect 329986 135088 330034 135144
rect 329925 135086 330034 135088
rect 329925 135083 329991 135086
rect 527766 135084 527772 135148
rect 527836 135146 527883 135148
rect 527836 135144 527928 135146
rect 527878 135088 527928 135144
rect 527836 135086 527928 135088
rect 527836 135084 527883 135086
rect 527817 135083 527883 135084
rect 583520 134874 584960 134964
rect 583342 134814 584960 134874
rect 376702 134540 376708 134604
rect 376772 134602 376778 134604
rect 381445 134602 381511 134605
rect 376772 134600 381511 134602
rect 376772 134544 381450 134600
rect 381506 134544 381511 134600
rect 376772 134542 381511 134544
rect 376772 134540 376778 134542
rect 381445 134539 381511 134542
rect 304942 134404 304948 134468
rect 305012 134466 305018 134468
rect 314561 134466 314627 134469
rect 305012 134464 314627 134466
rect 305012 134408 314566 134464
rect 314622 134408 314627 134464
rect 305012 134406 314627 134408
rect 305012 134404 305018 134406
rect 314561 134403 314627 134406
rect 417742 134406 424978 134466
rect 293769 134330 293835 134333
rect 295241 134330 295307 134333
rect 293769 134328 295307 134330
rect 293769 134272 293774 134328
rect 293830 134272 295246 134328
rect 295302 134272 295307 134328
rect 293769 134270 295307 134272
rect 293769 134267 293835 134270
rect 295241 134267 295307 134270
rect 367134 134268 367140 134332
rect 367204 134330 367210 134332
rect 376702 134330 376708 134332
rect 367204 134270 376708 134330
rect 367204 134268 367210 134270
rect 376702 134268 376708 134270
rect 376772 134268 376778 134332
rect 415301 134330 415367 134333
rect 408358 134328 415367 134330
rect 408358 134272 415306 134328
rect 415362 134272 415367 134328
rect 408358 134270 415367 134272
rect 314561 134194 314627 134197
rect 315982 134194 315988 134196
rect 314561 134192 315988 134194
rect 314561 134136 314566 134192
rect 314622 134136 315988 134192
rect 314561 134134 315988 134136
rect 314561 134131 314627 134134
rect 315982 134132 315988 134134
rect 316052 134132 316058 134196
rect 395981 134194 396047 134197
rect 408358 134194 408418 134270
rect 415301 134267 415367 134270
rect 395981 134192 408418 134194
rect 395981 134136 395986 134192
rect 396042 134136 408418 134192
rect 395981 134134 408418 134136
rect 415301 134194 415367 134197
rect 417742 134194 417802 134406
rect 415301 134192 417802 134194
rect 415301 134136 415306 134192
rect 415362 134136 417802 134192
rect 415301 134134 417802 134136
rect 424918 134194 424978 134406
rect 492630 134270 502258 134330
rect 427537 134194 427603 134197
rect 424918 134192 427603 134194
rect 424918 134136 427542 134192
rect 427598 134136 427603 134192
rect 424918 134134 427603 134136
rect 395981 134131 396047 134134
rect 415301 134131 415367 134134
rect 427537 134131 427603 134134
rect 427721 134194 427787 134197
rect 427721 134192 437490 134194
rect 427721 134136 427726 134192
rect 427782 134136 437490 134192
rect 427721 134134 437490 134136
rect 427721 134131 427787 134134
rect 284293 134058 284359 134061
rect 259502 134056 284359 134058
rect 259502 134000 284298 134056
rect 284354 134000 284359 134056
rect 259502 133998 284359 134000
rect 249374 133860 249380 133924
rect 249444 133922 249450 133924
rect 259502 133922 259562 133998
rect 284293 133995 284359 133998
rect 357382 133996 357388 134060
rect 357452 134058 357458 134060
rect 367134 134058 367140 134060
rect 357452 133998 367140 134058
rect 357452 133996 357458 133998
rect 367134 133996 367140 133998
rect 367204 133996 367210 134060
rect 381445 134058 381511 134061
rect 381445 134056 386522 134058
rect 381445 134000 381450 134056
rect 381506 134000 386522 134056
rect 381445 133998 386522 134000
rect 381445 133995 381511 133998
rect 249444 133862 259562 133922
rect 295241 133922 295307 133925
rect 295241 133920 295442 133922
rect 295241 133864 295246 133920
rect 295302 133864 295442 133920
rect 295241 133862 295442 133864
rect 249444 133860 249450 133862
rect 295241 133859 295307 133862
rect 295382 133786 295442 133862
rect 299614 133862 305010 133922
rect 299614 133786 299674 133862
rect 304950 133788 305010 133862
rect 315982 133860 315988 133924
rect 316052 133922 316058 133924
rect 325601 133922 325667 133925
rect 316052 133920 325667 133922
rect 316052 133864 325606 133920
rect 325662 133864 325667 133920
rect 316052 133862 325667 133864
rect 316052 133860 316058 133862
rect 325601 133859 325667 133862
rect 333881 133922 333947 133925
rect 343582 133922 343588 133924
rect 333881 133920 343588 133922
rect 333881 133864 333886 133920
rect 333942 133864 343588 133920
rect 333881 133862 343588 133864
rect 333881 133859 333947 133862
rect 343582 133860 343588 133862
rect 343652 133860 343658 133924
rect 295382 133726 299674 133786
rect 304942 133724 304948 133788
rect 305012 133724 305018 133788
rect 386462 133786 386522 133998
rect 437430 133922 437490 134134
rect 453982 134058 453988 134060
rect 447182 133998 453988 134058
rect 447182 133922 447242 133998
rect 453982 133996 453988 133998
rect 454052 133996 454058 134060
rect 458817 134058 458883 134061
rect 473302 134058 473308 134060
rect 458817 134056 466378 134058
rect 458817 134000 458822 134056
rect 458878 134000 466378 134056
rect 458817 133998 466378 134000
rect 458817 133995 458883 133998
rect 437430 133862 447242 133922
rect 466318 133922 466378 133998
rect 466502 133998 473308 134058
rect 466502 133922 466562 133998
rect 473302 133996 473308 133998
rect 473372 133996 473378 134060
rect 492630 134058 492690 134270
rect 502198 134196 502258 134270
rect 502190 134132 502196 134196
rect 502260 134132 502266 134196
rect 554497 134194 554563 134197
rect 554497 134192 563162 134194
rect 554497 134136 554502 134192
rect 554558 134136 563162 134192
rect 554497 134134 563162 134136
rect 554497 134131 554563 134134
rect 514569 134058 514635 134061
rect 485822 133998 492690 134058
rect 505142 134056 514635 134058
rect 505142 134000 514574 134056
rect 514630 134000 514635 134056
rect 505142 133998 514635 134000
rect 485822 133922 485882 133998
rect 466318 133862 466562 133922
rect 482878 133862 485882 133922
rect 395981 133786 396047 133789
rect 386462 133784 396047 133786
rect 386462 133728 395986 133784
rect 396042 133728 396047 133784
rect 386462 133726 396047 133728
rect 395981 133723 396047 133726
rect 453982 133724 453988 133788
rect 454052 133786 454058 133788
rect 458817 133786 458883 133789
rect 454052 133784 458883 133786
rect 454052 133728 458822 133784
rect 458878 133728 458883 133784
rect 454052 133726 458883 133728
rect 454052 133724 454058 133726
rect 458817 133723 458883 133726
rect 343582 133588 343588 133652
rect 343652 133650 343658 133652
rect 348417 133650 348483 133653
rect 343652 133648 348483 133650
rect 343652 133592 348422 133648
rect 348478 133592 348483 133648
rect 343652 133590 348483 133592
rect 343652 133588 343658 133590
rect 348417 133587 348483 133590
rect 354581 133650 354647 133653
rect 357198 133650 357204 133652
rect 354581 133648 357204 133650
rect 354581 133592 354586 133648
rect 354642 133592 357204 133648
rect 354581 133590 357204 133592
rect 354581 133587 354647 133590
rect 357198 133588 357204 133590
rect 357268 133588 357274 133652
rect 473302 133588 473308 133652
rect 473372 133650 473378 133652
rect 482878 133650 482938 133862
rect 502190 133860 502196 133924
rect 502260 133922 502266 133924
rect 505142 133922 505202 133998
rect 514569 133995 514635 133998
rect 514845 134058 514911 134061
rect 531262 134058 531268 134060
rect 514845 134056 524338 134058
rect 514845 134000 514850 134056
rect 514906 134000 524338 134056
rect 514845 133998 524338 134000
rect 514845 133995 514911 133998
rect 502260 133862 505202 133922
rect 524278 133922 524338 133998
rect 524462 133998 531268 134058
rect 524462 133922 524522 133998
rect 531262 133996 531268 133998
rect 531332 133996 531338 134060
rect 545849 134058 545915 134061
rect 550582 134058 550588 134060
rect 545849 134056 550588 134058
rect 545849 134000 545854 134056
rect 545910 134000 550588 134056
rect 545849 133998 550588 134000
rect 545849 133995 545915 133998
rect 550582 133996 550588 133998
rect 550652 133996 550658 134060
rect 540973 133922 541039 133925
rect 524278 133862 524522 133922
rect 540838 133920 541039 133922
rect 540838 133864 540978 133920
rect 541034 133864 541039 133920
rect 540838 133862 541039 133864
rect 563102 133922 563162 134134
rect 572621 134058 572687 134061
rect 583342 134058 583402 134814
rect 583520 134724 584960 134814
rect 569910 134056 572687 134058
rect 569910 134000 572626 134056
rect 572682 134000 572687 134056
rect 569910 133998 572687 134000
rect 569910 133922 569970 133998
rect 572621 133995 572687 133998
rect 576902 133998 583402 134058
rect 563102 133862 569970 133922
rect 572713 133922 572779 133925
rect 576902 133922 576962 133998
rect 572713 133920 576962 133922
rect 572713 133864 572718 133920
rect 572774 133864 576962 133920
rect 572713 133862 576962 133864
rect 502260 133860 502266 133862
rect 473372 133590 482938 133650
rect 473372 133588 473378 133590
rect 531262 133588 531268 133652
rect 531332 133650 531338 133652
rect 540838 133650 540898 133862
rect 540973 133859 541039 133862
rect 572713 133859 572779 133862
rect 550582 133724 550588 133788
rect 550652 133786 550658 133788
rect 554497 133786 554563 133789
rect 550652 133784 554563 133786
rect 550652 133728 554502 133784
rect 554558 133728 554563 133784
rect 550652 133726 554563 133728
rect 550652 133724 550658 133726
rect 554497 133723 554563 133726
rect 531332 133590 540898 133650
rect 531332 133588 531338 133590
rect 295701 131338 295767 131341
rect 295382 131336 295767 131338
rect 295382 131280 295706 131336
rect 295762 131280 295767 131336
rect 295382 131278 295767 131280
rect 295382 131202 295442 131278
rect 295701 131275 295767 131278
rect 295517 131202 295583 131205
rect 295382 131200 295583 131202
rect 295382 131144 295522 131200
rect 295578 131144 295583 131200
rect 295382 131142 295583 131144
rect 295517 131139 295583 131142
rect 230749 125626 230815 125629
rect 231025 125626 231091 125629
rect 230749 125624 231091 125626
rect 230749 125568 230754 125624
rect 230810 125568 231030 125624
rect 231086 125568 231091 125624
rect 230749 125566 231091 125568
rect 230749 125563 230815 125566
rect 231025 125563 231091 125566
rect 352005 125626 352071 125629
rect 352189 125626 352255 125629
rect 352005 125624 352255 125626
rect 352005 125568 352010 125624
rect 352066 125568 352194 125624
rect 352250 125568 352255 125624
rect 352005 125566 352255 125568
rect 352005 125563 352071 125566
rect 352189 125563 352255 125566
rect 527398 125564 527404 125628
rect 527468 125626 527474 125628
rect 527817 125626 527883 125629
rect 527468 125624 527883 125626
rect 527468 125568 527822 125624
rect 527878 125568 527883 125624
rect 527468 125566 527883 125568
rect 527468 125564 527474 125566
rect 527817 125563 527883 125566
rect 327165 124266 327231 124269
rect 327165 124264 327458 124266
rect 327165 124208 327170 124264
rect 327226 124208 327458 124264
rect 327165 124206 327458 124208
rect 327165 124203 327231 124206
rect 327165 123994 327231 123997
rect 327398 123994 327458 124206
rect 327165 123992 327458 123994
rect 327165 123936 327170 123992
rect 327226 123936 327458 123992
rect 327165 123934 327458 123936
rect 327165 123931 327231 123934
rect 580533 123178 580599 123181
rect 583520 123178 584960 123268
rect 580533 123176 584960 123178
rect 580533 123120 580538 123176
rect 580594 123120 584960 123176
rect 580533 123118 584960 123120
rect 580533 123115 580599 123118
rect 583520 123028 584960 123118
rect 324221 122770 324287 122773
rect 324405 122770 324471 122773
rect 324221 122768 324471 122770
rect 324221 122712 324226 122768
rect 324282 122712 324410 122768
rect 324466 122712 324471 122768
rect 324221 122710 324471 122712
rect 324221 122707 324287 122710
rect 324405 122707 324471 122710
rect -960 122090 480 122180
rect 3785 122090 3851 122093
rect -960 122088 3851 122090
rect -960 122032 3790 122088
rect 3846 122032 3851 122088
rect -960 122030 3851 122032
rect -960 121940 480 122030
rect 3785 122027 3851 122030
rect 527398 118764 527404 118828
rect 527468 118764 527474 118828
rect 527406 118554 527466 118764
rect 527582 118554 527588 118556
rect 527406 118494 527588 118554
rect 527582 118492 527588 118494
rect 527652 118492 527658 118556
rect 342529 116106 342595 116109
rect 348049 116106 348115 116109
rect 381261 116106 381327 116109
rect 342486 116104 342595 116106
rect 342486 116048 342534 116104
rect 342590 116048 342595 116104
rect 342486 116043 342595 116048
rect 348006 116104 348115 116106
rect 348006 116048 348054 116104
rect 348110 116048 348115 116104
rect 348006 116043 348115 116048
rect 381126 116104 381327 116106
rect 381126 116048 381266 116104
rect 381322 116048 381327 116104
rect 381126 116046 381327 116048
rect 342486 115973 342546 116043
rect 348006 115973 348066 116043
rect 381126 115973 381186 116046
rect 381261 116043 381327 116046
rect 241789 115970 241855 115973
rect 241973 115970 242039 115973
rect 241789 115968 242039 115970
rect 241789 115912 241794 115968
rect 241850 115912 241978 115968
rect 242034 115912 242039 115968
rect 241789 115910 242039 115912
rect 241789 115907 241855 115910
rect 241973 115907 242039 115910
rect 252737 115970 252803 115973
rect 252921 115970 252987 115973
rect 252737 115968 252987 115970
rect 252737 115912 252742 115968
rect 252798 115912 252926 115968
rect 252982 115912 252987 115968
rect 252737 115910 252987 115912
rect 252737 115907 252803 115910
rect 252921 115907 252987 115910
rect 254117 115970 254183 115973
rect 254301 115970 254367 115973
rect 254117 115968 254367 115970
rect 254117 115912 254122 115968
rect 254178 115912 254306 115968
rect 254362 115912 254367 115968
rect 254117 115910 254367 115912
rect 254117 115907 254183 115910
rect 254301 115907 254367 115910
rect 259637 115970 259703 115973
rect 259821 115970 259887 115973
rect 259637 115968 259887 115970
rect 259637 115912 259642 115968
rect 259698 115912 259826 115968
rect 259882 115912 259887 115968
rect 259637 115910 259887 115912
rect 259637 115907 259703 115910
rect 259821 115907 259887 115910
rect 265157 115970 265223 115973
rect 265341 115970 265407 115973
rect 266721 115970 266787 115973
rect 265157 115968 265407 115970
rect 265157 115912 265162 115968
rect 265218 115912 265346 115968
rect 265402 115912 265407 115968
rect 265157 115910 265407 115912
rect 265157 115907 265223 115910
rect 265341 115907 265407 115910
rect 266494 115968 266787 115970
rect 266494 115912 266726 115968
rect 266782 115912 266787 115968
rect 266494 115910 266787 115912
rect 266494 115837 266554 115910
rect 266721 115907 266787 115910
rect 267089 115970 267155 115973
rect 267273 115970 267339 115973
rect 267089 115968 267339 115970
rect 267089 115912 267094 115968
rect 267150 115912 267278 115968
rect 267334 115912 267339 115968
rect 267089 115910 267339 115912
rect 267089 115907 267155 115910
rect 267273 115907 267339 115910
rect 308029 115970 308095 115973
rect 308305 115970 308371 115973
rect 308029 115968 308371 115970
rect 308029 115912 308034 115968
rect 308090 115912 308310 115968
rect 308366 115912 308371 115968
rect 308029 115910 308371 115912
rect 308029 115907 308095 115910
rect 308305 115907 308371 115910
rect 342437 115968 342546 115973
rect 342437 115912 342442 115968
rect 342498 115912 342546 115968
rect 342437 115910 342546 115912
rect 347957 115968 348066 115973
rect 357709 115970 357775 115973
rect 347957 115912 347962 115968
rect 348018 115912 348066 115968
rect 347957 115910 348066 115912
rect 357574 115968 357775 115970
rect 357574 115912 357714 115968
rect 357770 115912 357775 115968
rect 357574 115910 357775 115912
rect 342437 115907 342503 115910
rect 347957 115907 348023 115910
rect 266494 115832 266603 115837
rect 266494 115776 266542 115832
rect 266598 115776 266603 115832
rect 266494 115774 266603 115776
rect 357574 115834 357634 115910
rect 357709 115907 357775 115910
rect 381077 115968 381186 115973
rect 381077 115912 381082 115968
rect 381138 115912 381186 115968
rect 381077 115910 381186 115912
rect 386597 115970 386663 115973
rect 386781 115970 386847 115973
rect 386597 115968 386847 115970
rect 386597 115912 386602 115968
rect 386658 115912 386786 115968
rect 386842 115912 386847 115968
rect 386597 115910 386847 115912
rect 381077 115907 381143 115910
rect 386597 115907 386663 115910
rect 386781 115907 386847 115910
rect 392117 115970 392183 115973
rect 392301 115970 392367 115973
rect 392117 115968 392367 115970
rect 392117 115912 392122 115968
rect 392178 115912 392306 115968
rect 392362 115912 392367 115968
rect 392117 115910 392367 115912
rect 392117 115907 392183 115910
rect 392301 115907 392367 115910
rect 416773 115970 416839 115973
rect 416957 115970 417023 115973
rect 416773 115968 417023 115970
rect 416773 115912 416778 115968
rect 416834 115912 416962 115968
rect 417018 115912 417023 115968
rect 416773 115910 417023 115912
rect 416773 115907 416839 115910
rect 416957 115907 417023 115910
rect 471973 115970 472039 115973
rect 472157 115970 472223 115973
rect 471973 115968 472223 115970
rect 471973 115912 471978 115968
rect 472034 115912 472162 115968
rect 472218 115912 472223 115968
rect 471973 115910 472223 115912
rect 471973 115907 472039 115910
rect 472157 115907 472223 115910
rect 357801 115834 357867 115837
rect 357574 115832 357867 115834
rect 357574 115776 357806 115832
rect 357862 115776 357867 115832
rect 357574 115774 357867 115776
rect 266537 115771 266603 115774
rect 357801 115771 357867 115774
rect 580165 111482 580231 111485
rect 583520 111482 584960 111572
rect 580165 111480 584960 111482
rect 580165 111424 580170 111480
rect 580226 111424 584960 111480
rect 580165 111422 584960 111424
rect 580165 111419 580231 111422
rect 583520 111332 584960 111422
rect 527214 108972 527220 109036
rect 527284 109034 527290 109036
rect 527766 109034 527772 109036
rect 527284 108974 527772 109034
rect 527284 108972 527290 108974
rect 527766 108972 527772 108974
rect 527836 108972 527842 109036
rect -960 107674 480 107764
rect 3601 107674 3667 107677
rect -960 107672 3667 107674
rect -960 107616 3606 107672
rect 3662 107616 3667 107672
rect -960 107614 3667 107616
rect -960 107524 480 107614
rect 3601 107611 3667 107614
rect 230749 106314 230815 106317
rect 231025 106314 231091 106317
rect 230749 106312 231091 106314
rect 230749 106256 230754 106312
rect 230810 106256 231030 106312
rect 231086 106256 231091 106312
rect 230749 106254 231091 106256
rect 230749 106251 230815 106254
rect 231025 106251 231091 106254
rect 236269 106314 236335 106317
rect 236453 106314 236519 106317
rect 236269 106312 236519 106314
rect 236269 106256 236274 106312
rect 236330 106256 236458 106312
rect 236514 106256 236519 106312
rect 236269 106254 236519 106256
rect 236269 106251 236335 106254
rect 236453 106251 236519 106254
rect 357617 106314 357683 106317
rect 357801 106314 357867 106317
rect 357617 106312 357867 106314
rect 357617 106256 357622 106312
rect 357678 106256 357806 106312
rect 357862 106256 357867 106312
rect 357617 106254 357867 106256
rect 357617 106251 357683 106254
rect 357801 106251 357867 106254
rect 400305 106314 400371 106317
rect 400489 106314 400555 106317
rect 400305 106312 400555 106314
rect 400305 106256 400310 106312
rect 400366 106256 400494 106312
rect 400550 106256 400555 106312
rect 400305 106254 400555 106256
rect 400305 106251 400371 106254
rect 400489 106251 400555 106254
rect 583520 99636 584960 99876
rect 527766 99514 527772 99516
rect 527590 99454 527772 99514
rect 527590 99244 527650 99454
rect 527766 99452 527772 99454
rect 527836 99452 527842 99516
rect 527582 99180 527588 99244
rect 527652 99180 527658 99244
rect 375741 96794 375807 96797
rect 375422 96792 375807 96794
rect 375422 96736 375746 96792
rect 375802 96736 375807 96792
rect 375422 96734 375807 96736
rect 236361 96658 236427 96661
rect 236545 96658 236611 96661
rect 236361 96656 236611 96658
rect 236361 96600 236366 96656
rect 236422 96600 236550 96656
rect 236606 96600 236611 96656
rect 236361 96598 236611 96600
rect 236361 96595 236427 96598
rect 236545 96595 236611 96598
rect 241789 96658 241855 96661
rect 241973 96658 242039 96661
rect 241789 96656 242039 96658
rect 241789 96600 241794 96656
rect 241850 96600 241978 96656
rect 242034 96600 242039 96656
rect 241789 96598 242039 96600
rect 241789 96595 241855 96598
rect 241973 96595 242039 96598
rect 259637 96658 259703 96661
rect 259821 96658 259887 96661
rect 259637 96656 259887 96658
rect 259637 96600 259642 96656
rect 259698 96600 259826 96656
rect 259882 96600 259887 96656
rect 259637 96598 259887 96600
rect 259637 96595 259703 96598
rect 259821 96595 259887 96598
rect 308029 96658 308095 96661
rect 308213 96658 308279 96661
rect 308029 96656 308279 96658
rect 308029 96600 308034 96656
rect 308090 96600 308218 96656
rect 308274 96600 308279 96656
rect 308029 96598 308279 96600
rect 308029 96595 308095 96598
rect 308213 96595 308279 96598
rect 370037 96658 370103 96661
rect 370221 96658 370287 96661
rect 370037 96656 370287 96658
rect 370037 96600 370042 96656
rect 370098 96600 370226 96656
rect 370282 96600 370287 96656
rect 370037 96598 370287 96600
rect 375422 96658 375482 96734
rect 375741 96731 375807 96734
rect 375557 96658 375623 96661
rect 375422 96656 375623 96658
rect 375422 96600 375562 96656
rect 375618 96600 375623 96656
rect 375422 96598 375623 96600
rect 370037 96595 370103 96598
rect 370221 96595 370287 96598
rect 375557 96595 375623 96598
rect 386597 96658 386663 96661
rect 386781 96658 386847 96661
rect 386597 96656 386847 96658
rect 386597 96600 386602 96656
rect 386658 96600 386786 96656
rect 386842 96600 386847 96656
rect 386597 96598 386847 96600
rect 386597 96595 386663 96598
rect 386781 96595 386847 96598
rect 392117 96658 392183 96661
rect 392301 96658 392367 96661
rect 392117 96656 392367 96658
rect 392117 96600 392122 96656
rect 392178 96600 392306 96656
rect 392362 96600 392367 96656
rect 392117 96598 392367 96600
rect 392117 96595 392183 96598
rect 392301 96595 392367 96598
rect 393221 96658 393287 96661
rect 393405 96658 393471 96661
rect 393221 96656 393471 96658
rect 393221 96600 393226 96656
rect 393282 96600 393410 96656
rect 393466 96600 393471 96656
rect 393221 96598 393471 96600
rect 393221 96595 393287 96598
rect 393405 96595 393471 96598
rect 400305 96658 400371 96661
rect 400581 96658 400647 96661
rect 400305 96656 400647 96658
rect 400305 96600 400310 96656
rect 400366 96600 400586 96656
rect 400642 96600 400647 96656
rect 400305 96598 400647 96600
rect 400305 96595 400371 96598
rect 400581 96595 400647 96598
rect 416773 96658 416839 96661
rect 416957 96658 417023 96661
rect 416773 96656 417023 96658
rect 416773 96600 416778 96656
rect 416834 96600 416962 96656
rect 417018 96600 417023 96656
rect 416773 96598 417023 96600
rect 416773 96595 416839 96598
rect 416957 96595 417023 96598
rect 433425 96658 433491 96661
rect 433701 96658 433767 96661
rect 433425 96656 433767 96658
rect 433425 96600 433430 96656
rect 433486 96600 433706 96656
rect 433762 96600 433767 96656
rect 433425 96598 433767 96600
rect 433425 96595 433491 96598
rect 433701 96595 433767 96598
rect 466453 96658 466519 96661
rect 466637 96658 466703 96661
rect 466453 96656 466703 96658
rect 466453 96600 466458 96656
rect 466514 96600 466642 96656
rect 466698 96600 466703 96656
rect 466453 96598 466703 96600
rect 466453 96595 466519 96598
rect 466637 96595 466703 96598
rect 471973 96658 472039 96661
rect 472157 96658 472223 96661
rect 471973 96656 472223 96658
rect 471973 96600 471978 96656
rect 472034 96600 472162 96656
rect 472218 96600 472223 96656
rect 471973 96598 472223 96600
rect 471973 96595 472039 96598
rect 472157 96595 472223 96598
rect 527449 96522 527515 96525
rect 527582 96522 527588 96524
rect 527449 96520 527588 96522
rect 527449 96464 527454 96520
rect 527510 96464 527588 96520
rect 527449 96462 527588 96464
rect 527449 96459 527515 96462
rect 527582 96460 527588 96462
rect 527652 96460 527658 96524
rect 324497 95298 324563 95301
rect 324681 95298 324747 95301
rect 324497 95296 324747 95298
rect 324497 95240 324502 95296
rect 324558 95240 324686 95296
rect 324742 95240 324747 95296
rect 324497 95238 324747 95240
rect 324497 95235 324563 95238
rect 324681 95235 324747 95238
rect -960 93258 480 93348
rect 3693 93258 3759 93261
rect -960 93256 3759 93258
rect -960 93200 3698 93256
rect 3754 93200 3759 93256
rect -960 93198 3759 93200
rect -960 93108 480 93198
rect 3693 93195 3759 93198
rect 580349 87954 580415 87957
rect 583520 87954 584960 88044
rect 580349 87952 584960 87954
rect 580349 87896 580354 87952
rect 580410 87896 584960 87952
rect 580349 87894 584960 87896
rect 580349 87891 580415 87894
rect 583520 87804 584960 87894
rect 236361 87138 236427 87141
rect 347957 87138 348023 87141
rect 352097 87138 352163 87141
rect 236134 87136 236427 87138
rect 236134 87080 236366 87136
rect 236422 87080 236427 87136
rect 236134 87078 236427 87080
rect 231945 87002 232011 87005
rect 232221 87002 232287 87005
rect 231945 87000 232287 87002
rect 231945 86944 231950 87000
rect 232006 86944 232226 87000
rect 232282 86944 232287 87000
rect 231945 86942 232287 86944
rect 236134 87002 236194 87078
rect 236361 87075 236427 87078
rect 347822 87136 348023 87138
rect 347822 87080 347962 87136
rect 348018 87080 348023 87136
rect 347822 87078 348023 87080
rect 347822 87005 347882 87078
rect 347957 87075 348023 87078
rect 352054 87136 352163 87138
rect 352054 87080 352102 87136
rect 352158 87080 352163 87136
rect 352054 87075 352163 87080
rect 352054 87005 352114 87075
rect 236269 87002 236335 87005
rect 236134 87000 236335 87002
rect 236134 86944 236274 87000
rect 236330 86944 236335 87000
rect 236134 86942 236335 86944
rect 347822 87000 347931 87005
rect 347822 86944 347870 87000
rect 347926 86944 347931 87000
rect 347822 86942 347931 86944
rect 231945 86939 232011 86942
rect 232221 86939 232287 86942
rect 236269 86939 236335 86942
rect 347865 86939 347931 86942
rect 352005 87000 352114 87005
rect 527449 87004 527515 87005
rect 527398 87002 527404 87004
rect 352005 86944 352010 87000
rect 352066 86944 352114 87000
rect 352005 86942 352114 86944
rect 527358 86942 527404 87002
rect 527468 87000 527515 87004
rect 527510 86944 527515 87000
rect 352005 86939 352071 86942
rect 527398 86940 527404 86942
rect 527468 86940 527515 86944
rect 527449 86939 527515 86940
rect 527398 80202 527404 80204
rect 527222 80142 527404 80202
rect 527222 79932 527282 80142
rect 527398 80140 527404 80142
rect 527468 80140 527474 80204
rect 527214 79868 527220 79932
rect 527284 79868 527290 79932
rect -960 78978 480 79068
rect 2773 78978 2839 78981
rect -960 78976 2839 78978
rect -960 78920 2778 78976
rect 2834 78920 2839 78976
rect -960 78918 2839 78920
rect -960 78828 480 78918
rect 2773 78915 2839 78918
rect 243118 77420 243124 77484
rect 243188 77482 243194 77484
rect 243261 77482 243327 77485
rect 243188 77480 243327 77482
rect 243188 77424 243266 77480
rect 243322 77424 243327 77480
rect 243188 77422 243327 77424
rect 243188 77420 243194 77422
rect 243261 77419 243327 77422
rect 357617 77346 357683 77349
rect 357801 77346 357867 77349
rect 357617 77344 357867 77346
rect 357617 77288 357622 77344
rect 357678 77288 357806 77344
rect 357862 77288 357867 77344
rect 357617 77286 357867 77288
rect 357617 77283 357683 77286
rect 357801 77283 357867 77286
rect 580441 76258 580507 76261
rect 583520 76258 584960 76348
rect 580441 76256 584960 76258
rect 580441 76200 580446 76256
rect 580502 76200 584960 76256
rect 580441 76198 584960 76200
rect 580441 76195 580507 76198
rect 583520 76108 584960 76198
rect 243077 75988 243143 75989
rect 243077 75984 243124 75988
rect 243188 75986 243194 75988
rect 243077 75928 243082 75984
rect 243077 75924 243124 75928
rect 243188 75926 243234 75986
rect 243188 75924 243194 75926
rect 243077 75923 243143 75924
rect 527214 70484 527220 70548
rect 527284 70484 527290 70548
rect 527222 70274 527282 70484
rect 527582 70274 527588 70276
rect 527222 70214 527588 70274
rect 527582 70212 527588 70214
rect 527652 70212 527658 70276
rect 393405 67826 393471 67829
rect 393086 67824 393471 67826
rect 393086 67768 393410 67824
rect 393466 67768 393471 67824
rect 393086 67766 393471 67768
rect 281809 67690 281875 67693
rect 281993 67690 282059 67693
rect 281809 67688 282059 67690
rect 281809 67632 281814 67688
rect 281870 67632 281998 67688
rect 282054 67632 282059 67688
rect 281809 67630 282059 67632
rect 393086 67690 393146 67766
rect 393405 67763 393471 67766
rect 393221 67690 393287 67693
rect 393086 67688 393287 67690
rect 393086 67632 393226 67688
rect 393282 67632 393287 67688
rect 393086 67630 393287 67632
rect 281809 67627 281875 67630
rect 281993 67627 282059 67630
rect 393221 67627 393287 67630
rect 387977 66330 388043 66333
rect 388161 66330 388227 66333
rect 387977 66328 388227 66330
rect 387977 66272 387982 66328
rect 388038 66272 388166 66328
rect 388222 66272 388227 66328
rect 387977 66270 388227 66272
rect 387977 66267 388043 66270
rect 388161 66267 388227 66270
rect -960 64562 480 64652
rect 3509 64562 3575 64565
rect -960 64560 3575 64562
rect -960 64504 3514 64560
rect 3570 64504 3575 64560
rect -960 64502 3575 64504
rect -960 64412 480 64502
rect 3509 64499 3575 64502
rect 580165 64562 580231 64565
rect 583520 64562 584960 64652
rect 580165 64560 584960 64562
rect 580165 64504 580170 64560
rect 580226 64504 584960 64560
rect 580165 64502 584960 64504
rect 580165 64499 580231 64502
rect 583520 64412 584960 64502
rect 527214 62732 527220 62796
rect 527284 62794 527290 62796
rect 527766 62794 527772 62796
rect 527284 62734 527772 62794
rect 527284 62732 527290 62734
rect 527766 62732 527772 62734
rect 527836 62732 527842 62796
rect 527214 57836 527220 57900
rect 527284 57836 527290 57900
rect 527222 57765 527282 57836
rect 527222 57760 527331 57765
rect 527222 57704 527270 57760
rect 527326 57704 527331 57760
rect 527222 57702 527331 57704
rect 527265 57699 527331 57702
rect 292481 55314 292547 55317
rect 292757 55314 292823 55317
rect 292481 55312 292823 55314
rect 292481 55256 292486 55312
rect 292542 55256 292762 55312
rect 292818 55256 292823 55312
rect 292481 55254 292823 55256
rect 292481 55251 292547 55254
rect 292757 55251 292823 55254
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 310697 48514 310763 48517
rect 310470 48512 310763 48514
rect 310470 48456 310702 48512
rect 310758 48456 310763 48512
rect 310470 48454 310763 48456
rect 310470 48378 310530 48454
rect 310697 48451 310763 48454
rect 310605 48378 310671 48381
rect 310470 48376 310671 48378
rect 310470 48320 310610 48376
rect 310666 48320 310671 48376
rect 310470 48318 310671 48320
rect 310605 48315 310671 48318
rect 527265 48378 527331 48381
rect 527398 48378 527404 48380
rect 527265 48376 527404 48378
rect 527265 48320 527270 48376
rect 527326 48320 527404 48376
rect 527265 48318 527404 48320
rect 527265 48315 527331 48318
rect 527398 48316 527404 48318
rect 527468 48316 527474 48380
rect 329925 45658 329991 45661
rect 329925 45656 330034 45658
rect 329925 45600 329930 45656
rect 329986 45600 330034 45656
rect 329925 45595 330034 45600
rect 329974 45522 330034 45595
rect 330109 45522 330175 45525
rect 329974 45520 330175 45522
rect 329974 45464 330114 45520
rect 330170 45464 330175 45520
rect 329974 45462 330175 45464
rect 330109 45459 330175 45462
rect 527398 41516 527404 41580
rect 527468 41516 527474 41580
rect 527406 41306 527466 41516
rect 527582 41306 527588 41308
rect 527406 41246 527588 41306
rect 527582 41244 527588 41246
rect 527652 41244 527658 41308
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 373901 40628 373967 40629
rect 373901 40624 373948 40628
rect 374012 40626 374018 40628
rect 373901 40568 373906 40624
rect 373901 40564 373948 40568
rect 374012 40566 374094 40626
rect 374012 40564 374018 40566
rect 373901 40563 373967 40564
rect 253798 40430 254042 40490
rect 253798 40218 253858 40430
rect 253982 40354 254042 40430
rect 354622 40428 354628 40492
rect 354692 40490 354698 40492
rect 364241 40490 364307 40493
rect 354692 40488 364307 40490
rect 354692 40432 364246 40488
rect 364302 40432 364307 40488
rect 354692 40430 364307 40432
rect 354692 40428 354698 40430
rect 364241 40427 364307 40430
rect 492630 40430 502258 40490
rect 273069 40354 273135 40357
rect 253982 40352 273135 40354
rect 253982 40296 273074 40352
rect 273130 40296 273135 40352
rect 253982 40294 273135 40296
rect 273069 40291 273135 40294
rect 273253 40354 273319 40357
rect 273253 40352 284954 40354
rect 273253 40296 273258 40352
rect 273314 40296 284954 40352
rect 273253 40294 284954 40296
rect 273253 40291 273319 40294
rect 234662 40158 253858 40218
rect 284894 40218 284954 40294
rect 335302 40292 335308 40356
rect 335372 40354 335378 40356
rect 344921 40354 344987 40357
rect 335372 40352 344987 40354
rect 335372 40296 344926 40352
rect 344982 40296 344987 40352
rect 335372 40294 344987 40296
rect 335372 40292 335378 40294
rect 344921 40291 344987 40294
rect 373942 40292 373948 40356
rect 374012 40354 374018 40356
rect 397637 40354 397703 40357
rect 374012 40294 374194 40354
rect 374012 40292 374018 40294
rect 289813 40218 289879 40221
rect 284894 40216 289879 40218
rect 284894 40160 289818 40216
rect 289874 40160 289879 40216
rect 284894 40158 289879 40160
rect 234470 40020 234476 40084
rect 234540 40082 234546 40084
rect 234662 40082 234722 40158
rect 289813 40155 289879 40158
rect 307293 40218 307359 40221
rect 335261 40218 335327 40221
rect 354622 40218 354628 40220
rect 307293 40216 335327 40218
rect 307293 40160 307298 40216
rect 307354 40160 335266 40216
rect 335322 40160 335327 40216
rect 307293 40158 335327 40160
rect 307293 40155 307359 40158
rect 335261 40155 335327 40158
rect 345062 40158 354628 40218
rect 234540 40022 234722 40082
rect 289813 40082 289879 40085
rect 302141 40082 302207 40085
rect 289813 40080 302207 40082
rect 289813 40024 289818 40080
rect 289874 40024 302146 40080
rect 302202 40024 302207 40080
rect 289813 40022 302207 40024
rect 234540 40020 234546 40022
rect 289813 40019 289879 40022
rect 302141 40019 302207 40022
rect 335261 40084 335327 40085
rect 335261 40080 335308 40084
rect 335372 40082 335378 40084
rect 344921 40082 344987 40085
rect 345062 40082 345122 40158
rect 354622 40156 354628 40158
rect 354692 40156 354698 40220
rect 364241 40218 364307 40221
rect 373901 40218 373967 40221
rect 364241 40216 373967 40218
rect 364241 40160 364246 40216
rect 364302 40160 373906 40216
rect 373962 40160 373967 40216
rect 364241 40158 373967 40160
rect 374134 40218 374194 40294
rect 389222 40352 397703 40354
rect 389222 40296 397642 40352
rect 397698 40296 397703 40352
rect 389222 40294 397703 40296
rect 389222 40218 389282 40294
rect 397637 40291 397703 40294
rect 405641 40354 405707 40357
rect 418061 40354 418127 40357
rect 456793 40354 456859 40357
rect 405641 40352 408418 40354
rect 405641 40296 405646 40352
rect 405702 40296 408418 40352
rect 405641 40294 408418 40296
rect 405641 40291 405707 40294
rect 374134 40158 389282 40218
rect 364241 40155 364307 40158
rect 373901 40155 373967 40158
rect 335261 40024 335266 40080
rect 335261 40020 335308 40024
rect 335372 40022 335454 40082
rect 344921 40080 345122 40082
rect 344921 40024 344926 40080
rect 344982 40024 345122 40080
rect 344921 40022 345122 40024
rect 408358 40082 408418 40294
rect 415350 40352 418127 40354
rect 415350 40296 418066 40352
rect 418122 40296 418127 40352
rect 415350 40294 418127 40296
rect 415350 40218 415410 40294
rect 418061 40291 418127 40294
rect 424918 40294 427738 40354
rect 408542 40158 415410 40218
rect 418153 40218 418219 40221
rect 424918 40218 424978 40294
rect 418153 40216 424978 40218
rect 418153 40160 418158 40216
rect 418214 40160 424978 40216
rect 418153 40158 424978 40160
rect 408542 40082 408602 40158
rect 418153 40155 418219 40158
rect 408358 40022 408602 40082
rect 427678 40082 427738 40294
rect 427862 40294 437490 40354
rect 427862 40082 427922 40294
rect 427678 40022 427922 40082
rect 437430 40082 437490 40294
rect 456793 40352 456994 40354
rect 456793 40296 456798 40352
rect 456854 40296 456994 40352
rect 456793 40294 456994 40296
rect 456793 40291 456859 40294
rect 456701 40218 456767 40221
rect 447182 40216 456767 40218
rect 447182 40160 456706 40216
rect 456762 40160 456767 40216
rect 447182 40158 456767 40160
rect 456934 40218 456994 40294
rect 475929 40218 475995 40221
rect 456934 40158 466378 40218
rect 447182 40082 447242 40158
rect 456701 40155 456767 40158
rect 437430 40022 447242 40082
rect 466318 40082 466378 40158
rect 466502 40216 475995 40218
rect 466502 40160 475934 40216
rect 475990 40160 475995 40216
rect 466502 40158 475995 40160
rect 466502 40082 466562 40158
rect 475929 40155 475995 40158
rect 478229 40218 478295 40221
rect 492630 40218 492690 40430
rect 502198 40356 502258 40430
rect 502190 40292 502196 40356
rect 502260 40292 502266 40356
rect 554497 40354 554563 40357
rect 554497 40352 563162 40354
rect 554497 40296 554502 40352
rect 554558 40296 563162 40352
rect 554497 40294 563162 40296
rect 554497 40291 554563 40294
rect 514569 40218 514635 40221
rect 478229 40216 482938 40218
rect 478229 40160 478234 40216
rect 478290 40160 482938 40216
rect 478229 40158 482938 40160
rect 478229 40155 478295 40158
rect 466318 40022 466562 40082
rect 482878 40082 482938 40158
rect 485822 40158 492690 40218
rect 505142 40216 514635 40218
rect 505142 40160 514574 40216
rect 514630 40160 514635 40216
rect 505142 40158 514635 40160
rect 485822 40082 485882 40158
rect 482878 40022 485882 40082
rect 335372 40020 335378 40022
rect 335261 40019 335327 40020
rect 344921 40019 344987 40022
rect 502190 40020 502196 40084
rect 502260 40082 502266 40084
rect 505142 40082 505202 40158
rect 514569 40155 514635 40158
rect 514845 40218 514911 40221
rect 531262 40218 531268 40220
rect 514845 40216 524338 40218
rect 514845 40160 514850 40216
rect 514906 40160 524338 40216
rect 514845 40158 524338 40160
rect 514845 40155 514911 40158
rect 502260 40022 505202 40082
rect 524278 40082 524338 40158
rect 524462 40158 531268 40218
rect 524462 40082 524522 40158
rect 531262 40156 531268 40158
rect 531332 40156 531338 40220
rect 545849 40218 545915 40221
rect 550582 40218 550588 40220
rect 545849 40216 550588 40218
rect 545849 40160 545854 40216
rect 545910 40160 550588 40216
rect 545849 40158 550588 40160
rect 545849 40155 545915 40158
rect 550582 40156 550588 40158
rect 550652 40156 550658 40220
rect 540973 40082 541039 40085
rect 524278 40022 524522 40082
rect 540838 40080 541039 40082
rect 540838 40024 540978 40080
rect 541034 40024 541039 40080
rect 540838 40022 541039 40024
rect 563102 40082 563162 40294
rect 572621 40218 572687 40221
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 569910 40216 572687 40218
rect 569910 40160 572626 40216
rect 572682 40160 572687 40216
rect 569910 40158 572687 40160
rect 569910 40082 569970 40158
rect 572621 40155 572687 40158
rect 576902 40158 583402 40218
rect 563102 40022 569970 40082
rect 572713 40082 572779 40085
rect 576902 40082 576962 40158
rect 572713 40080 576962 40082
rect 572713 40024 572718 40080
rect 572774 40024 576962 40080
rect 572713 40022 576962 40024
rect 502260 40020 502266 40022
rect 531262 39748 531268 39812
rect 531332 39810 531338 39812
rect 540838 39810 540898 40022
rect 540973 40019 541039 40022
rect 572713 40019 572779 40022
rect 550582 39884 550588 39948
rect 550652 39946 550658 39948
rect 554497 39946 554563 39949
rect 550652 39944 554563 39946
rect 550652 39888 554502 39944
rect 554558 39888 554563 39944
rect 550652 39886 554563 39888
rect 550652 39884 550658 39886
rect 554497 39883 554563 39886
rect 531332 39750 540898 39810
rect 531332 39748 531338 39750
rect 527449 38586 527515 38589
rect 527582 38586 527588 38588
rect 527449 38584 527588 38586
rect 527449 38528 527454 38584
rect 527510 38528 527588 38584
rect 527449 38526 527588 38528
rect 527449 38523 527515 38526
rect 527582 38524 527588 38526
rect 527652 38524 527658 38588
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580257 29338 580323 29341
rect 583520 29338 584960 29428
rect 580257 29336 584960 29338
rect 580257 29280 580262 29336
rect 580318 29280 584960 29336
rect 580257 29278 584960 29280
rect 580257 29275 580323 29278
rect 527449 29202 527515 29205
rect 527406 29200 527515 29202
rect 527406 29144 527454 29200
rect 527510 29144 527515 29200
rect 583520 29188 584960 29278
rect 527406 29139 527515 29144
rect 527406 29068 527466 29139
rect 527398 29004 527404 29068
rect 527468 29004 527474 29068
rect 310421 28930 310487 28933
rect 310605 28930 310671 28933
rect 310421 28928 310671 28930
rect 310421 28872 310426 28928
rect 310482 28872 310610 28928
rect 310666 28872 310671 28928
rect 310421 28870 310671 28872
rect 310421 28867 310487 28870
rect 310605 28867 310671 28870
rect 422109 27570 422175 27573
rect 422293 27570 422359 27573
rect 422109 27568 422359 27570
rect 422109 27512 422114 27568
rect 422170 27512 422298 27568
rect 422354 27512 422359 27568
rect 422109 27510 422359 27512
rect 422109 27507 422175 27510
rect 422293 27507 422359 27510
rect 427905 24850 427971 24853
rect 428089 24850 428155 24853
rect 427905 24848 428155 24850
rect 427905 24792 427910 24848
rect 427966 24792 428094 24848
rect 428150 24792 428155 24848
rect 427905 24790 428155 24792
rect 427905 24787 427971 24790
rect 428089 24787 428155 24790
rect 521653 22266 521719 22269
rect 527398 22266 527404 22268
rect 521653 22264 527404 22266
rect 521653 22208 521658 22264
rect 521714 22208 527404 22264
rect 521653 22206 527404 22208
rect 521653 22203 521719 22206
rect 527398 22204 527404 22206
rect 527468 22204 527474 22268
rect 521653 21994 521719 21997
rect 614 21992 521719 21994
rect 614 21936 521658 21992
rect 521714 21936 521719 21992
rect 614 21934 521719 21936
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 521653 21931 521719 21934
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 583520 17642 584960 17732
rect 583342 17582 584960 17642
rect 550582 17308 550588 17372
rect 550652 17370 550658 17372
rect 560201 17370 560267 17373
rect 550652 17368 560267 17370
rect 550652 17312 560206 17368
rect 560262 17312 560267 17368
rect 550652 17310 560267 17312
rect 550652 17308 550658 17310
rect 560201 17307 560267 17310
rect 259494 17172 259500 17236
rect 259564 17234 259570 17236
rect 269021 17234 269087 17237
rect 259564 17232 269087 17234
rect 259564 17176 269026 17232
rect 269082 17176 269087 17232
rect 259564 17174 269087 17176
rect 259564 17172 259570 17174
rect 269021 17171 269087 17174
rect 325734 17172 325740 17236
rect 325804 17234 325810 17236
rect 335261 17234 335327 17237
rect 325804 17232 335327 17234
rect 325804 17176 335266 17232
rect 335322 17176 335327 17232
rect 325804 17174 335327 17176
rect 325804 17172 325810 17174
rect 335261 17171 335327 17174
rect 531262 17172 531268 17236
rect 531332 17234 531338 17236
rect 540881 17234 540947 17237
rect 531332 17232 540947 17234
rect 531332 17176 540886 17232
rect 540942 17176 540947 17232
rect 531332 17174 540947 17176
rect 531332 17172 531338 17174
rect 540881 17171 540947 17174
rect 410701 17098 410767 17101
rect 418061 17098 418127 17101
rect 502006 17098 502012 17100
rect 410701 17096 418127 17098
rect 410701 17040 410706 17096
rect 410762 17040 418066 17096
rect 418122 17040 418127 17096
rect 410701 17038 418127 17040
rect 410701 17035 410767 17038
rect 418061 17035 418127 17038
rect 495206 17038 502012 17098
rect 259494 16962 259500 16964
rect 251038 16902 259500 16962
rect 231710 16764 231716 16828
rect 231780 16826 231786 16828
rect 244181 16826 244247 16829
rect 231780 16824 244247 16826
rect 231780 16768 244186 16824
rect 244242 16768 244247 16824
rect 231780 16766 244247 16768
rect 231780 16764 231786 16766
rect 244181 16763 244247 16766
rect 244365 16826 244431 16829
rect 251038 16826 251098 16902
rect 259494 16900 259500 16902
rect 259564 16900 259570 16964
rect 278773 16962 278839 16965
rect 270358 16960 278839 16962
rect 270358 16904 278778 16960
rect 278834 16904 278839 16960
rect 270358 16902 278839 16904
rect 244365 16824 251098 16826
rect 244365 16768 244370 16824
rect 244426 16768 251098 16824
rect 244365 16766 251098 16768
rect 269021 16826 269087 16829
rect 270358 16826 270418 16902
rect 278773 16899 278839 16902
rect 323577 16962 323643 16965
rect 325734 16962 325740 16964
rect 323577 16960 325740 16962
rect 323577 16904 323582 16960
rect 323638 16904 325740 16960
rect 323577 16902 325740 16904
rect 323577 16899 323643 16902
rect 325734 16900 325740 16902
rect 325804 16900 325810 16964
rect 355961 16962 356027 16965
rect 357382 16962 357388 16964
rect 355961 16960 357388 16962
rect 355961 16904 355966 16960
rect 356022 16904 357388 16960
rect 355961 16902 357388 16904
rect 355961 16899 356027 16902
rect 357382 16900 357388 16902
rect 357452 16900 357458 16964
rect 418245 16962 418311 16965
rect 456793 16962 456859 16965
rect 375238 16902 381554 16962
rect 269021 16824 270418 16826
rect 269021 16768 269026 16824
rect 269082 16768 270418 16824
rect 269021 16766 270418 16768
rect 309041 16826 309107 16829
rect 323485 16826 323551 16829
rect 309041 16824 311818 16826
rect 309041 16768 309046 16824
rect 309102 16768 311818 16824
rect 309041 16766 311818 16768
rect 244365 16763 244431 16766
rect 269021 16763 269087 16766
rect 309041 16763 309107 16766
rect 288341 16690 288407 16693
rect 299289 16690 299355 16693
rect 299422 16690 299428 16692
rect 288341 16688 289922 16690
rect 288341 16632 288346 16688
rect 288402 16632 289922 16688
rect 288341 16630 289922 16632
rect 288341 16627 288407 16630
rect 289862 16554 289922 16630
rect 299289 16688 299428 16690
rect 299289 16632 299294 16688
rect 299350 16632 299428 16688
rect 299289 16630 299428 16632
rect 299289 16627 299355 16630
rect 299422 16628 299428 16630
rect 299492 16628 299498 16692
rect 311758 16690 311818 16766
rect 317462 16824 323551 16826
rect 317462 16768 323490 16824
rect 323546 16768 323551 16824
rect 317462 16766 323551 16768
rect 317462 16690 317522 16766
rect 323485 16763 323551 16766
rect 335261 16826 335327 16829
rect 370497 16826 370563 16829
rect 375238 16826 375298 16902
rect 335261 16824 337946 16826
rect 335261 16768 335266 16824
rect 335322 16768 337946 16824
rect 335261 16766 337946 16768
rect 335261 16763 335327 16766
rect 311758 16630 317522 16690
rect 337886 16690 337946 16766
rect 370497 16824 375298 16826
rect 370497 16768 370502 16824
rect 370558 16768 375298 16824
rect 370497 16766 375298 16768
rect 381494 16826 381554 16902
rect 418245 16960 427738 16962
rect 418245 16904 418250 16960
rect 418306 16904 427738 16960
rect 418245 16902 427738 16904
rect 418245 16899 418311 16902
rect 386505 16826 386571 16829
rect 381494 16824 386571 16826
rect 381494 16768 386510 16824
rect 386566 16768 386571 16824
rect 381494 16766 386571 16768
rect 370497 16763 370563 16766
rect 386505 16763 386571 16766
rect 398925 16826 398991 16829
rect 408401 16826 408467 16829
rect 398925 16824 408467 16826
rect 398925 16768 398930 16824
rect 398986 16768 408406 16824
rect 408462 16768 408467 16824
rect 398925 16766 408467 16768
rect 398925 16763 398991 16766
rect 408401 16763 408467 16766
rect 346209 16690 346275 16693
rect 347681 16690 347747 16693
rect 337886 16688 346275 16690
rect 337886 16632 346214 16688
rect 346270 16632 346275 16688
rect 337886 16630 346275 16632
rect 346209 16627 346275 16630
rect 346350 16688 347747 16690
rect 346350 16632 347686 16688
rect 347742 16632 347747 16688
rect 346350 16630 347747 16632
rect 299289 16554 299355 16557
rect 289862 16552 299355 16554
rect 289862 16496 299294 16552
rect 299350 16496 299355 16552
rect 289862 16494 299355 16496
rect 299289 16491 299355 16494
rect 346209 16554 346275 16557
rect 346350 16554 346410 16630
rect 347681 16627 347747 16630
rect 357566 16628 357572 16692
rect 357636 16690 357642 16692
rect 365662 16690 365668 16692
rect 357636 16630 365668 16690
rect 357636 16628 357642 16630
rect 365662 16628 365668 16630
rect 365732 16628 365738 16692
rect 427678 16690 427738 16902
rect 427862 16902 437490 16962
rect 427862 16690 427922 16902
rect 427678 16630 427922 16690
rect 437430 16690 437490 16902
rect 456793 16960 456994 16962
rect 456793 16904 456798 16960
rect 456854 16904 456994 16960
rect 456793 16902 456994 16904
rect 456793 16899 456859 16902
rect 456701 16826 456767 16829
rect 447182 16824 456767 16826
rect 447182 16768 456706 16824
rect 456762 16768 456767 16824
rect 447182 16766 456767 16768
rect 456934 16826 456994 16902
rect 475929 16826 475995 16829
rect 456934 16766 466378 16826
rect 447182 16690 447242 16766
rect 456701 16763 456767 16766
rect 437430 16630 447242 16690
rect 466318 16690 466378 16766
rect 466502 16824 475995 16826
rect 466502 16768 475934 16824
rect 475990 16768 475995 16824
rect 466502 16766 475995 16768
rect 466502 16690 466562 16766
rect 475929 16763 475995 16766
rect 477493 16826 477559 16829
rect 495206 16826 495266 17038
rect 502006 17036 502012 17038
rect 502076 17036 502082 17100
rect 550582 17098 550588 17100
rect 543782 17038 550588 17098
rect 524505 16962 524571 16965
rect 531262 16962 531268 16964
rect 524505 16960 531268 16962
rect 524505 16904 524510 16960
rect 524566 16904 531268 16960
rect 524505 16902 531268 16904
rect 524505 16899 524571 16902
rect 531262 16900 531268 16902
rect 531332 16900 531338 16964
rect 514569 16826 514635 16829
rect 477493 16824 482938 16826
rect 477493 16768 477498 16824
rect 477554 16768 482938 16824
rect 477493 16766 482938 16768
rect 477493 16763 477559 16766
rect 466318 16630 466562 16690
rect 482878 16690 482938 16766
rect 485822 16766 495266 16826
rect 505142 16824 514635 16826
rect 505142 16768 514574 16824
rect 514630 16768 514635 16824
rect 505142 16766 514635 16768
rect 485822 16690 485882 16766
rect 482878 16630 485882 16690
rect 502190 16628 502196 16692
rect 502260 16690 502266 16692
rect 505142 16690 505202 16766
rect 514569 16763 514635 16766
rect 540881 16826 540947 16829
rect 543782 16826 543842 17038
rect 550582 17036 550588 17038
rect 550652 17036 550658 17100
rect 560201 16962 560267 16965
rect 560201 16960 563162 16962
rect 560201 16904 560206 16960
rect 560262 16904 563162 16960
rect 560201 16902 563162 16904
rect 560201 16899 560267 16902
rect 540881 16824 543842 16826
rect 540881 16768 540886 16824
rect 540942 16768 543842 16824
rect 540881 16766 543842 16768
rect 540881 16763 540947 16766
rect 521653 16690 521719 16693
rect 502260 16630 505202 16690
rect 521518 16688 521719 16690
rect 521518 16632 521658 16688
rect 521714 16632 521719 16688
rect 521518 16630 521719 16632
rect 563102 16690 563162 16902
rect 572621 16826 572687 16829
rect 583342 16826 583402 17582
rect 583520 17492 584960 17582
rect 569910 16824 572687 16826
rect 569910 16768 572626 16824
rect 572682 16768 572687 16824
rect 569910 16766 572687 16768
rect 569910 16690 569970 16766
rect 572621 16763 572687 16766
rect 576902 16766 583402 16826
rect 563102 16630 569970 16690
rect 572713 16690 572779 16693
rect 576902 16690 576962 16766
rect 572713 16688 576962 16690
rect 572713 16632 572718 16688
rect 572774 16632 576962 16688
rect 572713 16630 576962 16632
rect 502260 16628 502266 16630
rect 346209 16552 346410 16554
rect 346209 16496 346214 16552
rect 346270 16496 346410 16552
rect 346209 16494 346410 16496
rect 386505 16554 386571 16557
rect 395838 16554 395844 16556
rect 386505 16552 395844 16554
rect 386505 16496 386510 16552
rect 386566 16496 395844 16552
rect 386505 16494 395844 16496
rect 346209 16491 346275 16494
rect 386505 16491 386571 16494
rect 395838 16492 395844 16494
rect 395908 16492 395914 16556
rect 396022 16492 396028 16556
rect 396092 16554 396098 16556
rect 398925 16554 398991 16557
rect 396092 16552 398991 16554
rect 396092 16496 398930 16552
rect 398986 16496 398991 16552
rect 396092 16494 398991 16496
rect 396092 16492 396098 16494
rect 398925 16491 398991 16494
rect 299422 16356 299428 16420
rect 299492 16418 299498 16420
rect 309041 16418 309107 16421
rect 299492 16416 309107 16418
rect 299492 16360 309046 16416
rect 309102 16360 309107 16416
rect 299492 16358 309107 16360
rect 299492 16356 299498 16358
rect 309041 16355 309107 16358
rect 365662 16356 365668 16420
rect 365732 16418 365738 16420
rect 370497 16418 370563 16421
rect 365732 16416 370563 16418
rect 365732 16360 370502 16416
rect 370558 16360 370563 16416
rect 365732 16358 370563 16360
rect 365732 16356 365738 16358
rect 370497 16355 370563 16358
rect 514569 16418 514635 16421
rect 521518 16418 521578 16630
rect 521653 16627 521719 16630
rect 572713 16627 572779 16630
rect 514569 16416 521578 16418
rect 514569 16360 514574 16416
rect 514630 16360 521578 16416
rect 514569 16358 521578 16360
rect 514569 16355 514635 16358
rect 60641 10298 60707 10301
rect 259821 10298 259887 10301
rect 60641 10296 259887 10298
rect 60641 10240 60646 10296
rect 60702 10240 259826 10296
rect 259882 10240 259887 10296
rect 60641 10238 259887 10240
rect 60641 10235 60707 10238
rect 259821 10235 259887 10238
rect 136081 8938 136147 8941
rect 299565 8938 299631 8941
rect 136081 8936 299631 8938
rect 136081 8880 136086 8936
rect 136142 8880 299570 8936
rect 299626 8880 299631 8936
rect 136081 8878 299631 8880
rect 136081 8875 136147 8878
rect 299565 8875 299631 8878
rect 277485 8530 277551 8533
rect 277485 8528 277778 8530
rect 277485 8472 277490 8528
rect 277546 8472 277778 8528
rect 277485 8470 277778 8472
rect 277485 8467 277551 8470
rect 277577 8394 277643 8397
rect 277718 8394 277778 8470
rect 277577 8392 277778 8394
rect 277577 8336 277582 8392
rect 277638 8336 277778 8392
rect 277577 8334 277778 8336
rect 277577 8331 277643 8334
rect 134885 7578 134951 7581
rect 298277 7578 298343 7581
rect 134885 7576 298343 7578
rect 134885 7520 134890 7576
rect 134946 7520 298282 7576
rect 298338 7520 298343 7576
rect 134885 7518 298343 7520
rect 134885 7515 134951 7518
rect 298277 7515 298343 7518
rect -960 7170 480 7260
rect 4061 7170 4127 7173
rect -960 7168 4127 7170
rect -960 7112 4066 7168
rect 4122 7112 4127 7168
rect -960 7110 4127 7112
rect -960 7020 480 7110
rect 4061 7107 4127 7110
rect 48129 6218 48195 6221
rect 253933 6218 253999 6221
rect 48129 6216 253999 6218
rect 48129 6160 48134 6216
rect 48190 6160 253938 6216
rect 253994 6160 253999 6216
rect 48129 6158 253999 6160
rect 48129 6155 48195 6158
rect 253933 6155 253999 6158
rect 583520 5796 584960 6036
rect 219341 4858 219407 4861
rect 342253 4858 342319 4861
rect 219341 4856 342319 4858
rect 219341 4800 219346 4856
rect 219402 4800 342258 4856
rect 342314 4800 342319 4856
rect 219341 4798 342319 4800
rect 219341 4795 219407 4798
rect 342253 4795 342319 4798
rect 408401 3906 408467 3909
rect 408585 3906 408651 3909
rect 408401 3904 408651 3906
rect 408401 3848 408406 3904
rect 408462 3848 408590 3904
rect 408646 3848 408651 3904
rect 408401 3846 408651 3848
rect 408401 3843 408467 3846
rect 408585 3843 408651 3846
rect 408309 3634 408375 3637
rect 408585 3634 408651 3637
rect 408309 3632 408651 3634
rect 408309 3576 408314 3632
rect 408370 3576 408590 3632
rect 408646 3576 408651 3632
rect 408309 3574 408651 3576
rect 408309 3571 408375 3574
rect 408585 3571 408651 3574
rect 6453 3362 6519 3365
rect 231945 3362 232011 3365
rect 6453 3360 232011 3362
rect 6453 3304 6458 3360
rect 6514 3304 231950 3360
rect 232006 3304 232011 3360
rect 6453 3302 232011 3304
rect 6453 3299 6519 3302
rect 231945 3299 232011 3302
rect 356145 3362 356211 3365
rect 410609 3362 410675 3365
rect 356145 3360 410675 3362
rect 356145 3304 356150 3360
rect 356206 3304 410614 3360
rect 410670 3304 410675 3360
rect 356145 3302 410675 3304
rect 356145 3299 356211 3302
rect 410609 3299 410675 3302
rect 525701 3362 525767 3365
rect 575013 3362 575079 3365
rect 525701 3360 575079 3362
rect 525701 3304 525706 3360
rect 525762 3304 575018 3360
rect 575074 3304 575079 3360
rect 525701 3302 575079 3304
rect 525701 3299 525767 3302
rect 575013 3299 575079 3302
<< via3 >>
rect 233740 642908 233804 642972
rect 526116 642908 526180 642972
rect 232820 642636 232884 642700
rect 232636 642500 232700 642564
rect 232452 642364 232516 642428
rect 434484 642092 434548 642156
rect 7420 641548 7484 641612
rect 12940 641548 13004 641612
rect 27660 641548 27724 641612
rect 79732 641548 79796 641612
rect 109724 641548 109788 641612
rect 137324 641548 137388 641612
rect 167316 641548 167380 641612
rect 215156 641548 215220 641612
rect 222148 641548 222212 641612
rect 226012 641548 226076 641612
rect 231900 641548 231964 641612
rect 282684 641548 282748 641612
rect 301636 641548 301700 641612
rect 302924 641548 302988 641612
rect 309364 641548 309428 641612
rect 318380 641548 318444 641612
rect 327028 641548 327092 641612
rect 336596 641548 336660 641612
rect 348372 641548 348436 641612
rect 351132 641548 351196 641612
rect 376708 641548 376772 641612
rect 379652 641548 379716 641612
rect 423628 641548 423692 641612
rect 432460 641548 432524 641612
rect 453988 641548 454052 641612
rect 463556 641548 463620 641612
rect 80836 640868 80900 640932
rect 108436 640868 108500 640932
rect 138428 640868 138492 640932
rect 166028 640868 166092 640932
rect 251772 640868 251836 640932
rect 264468 640868 264532 640932
rect 289860 640868 289924 640932
rect 299244 640868 299308 640932
rect 318748 640868 318812 640932
rect 322060 640868 322124 640932
rect 357388 640868 357452 640932
rect 366956 640868 367020 640932
rect 367140 640868 367204 640932
rect 376524 640868 376588 640932
rect 389036 640868 389100 640932
rect 395660 640868 395724 640932
rect 396028 640868 396092 640932
rect 399340 640868 399404 640932
rect 436140 640868 436204 640932
rect 438532 640868 438596 640932
rect 463924 640188 463988 640252
rect 480852 640188 480916 640252
rect 509188 640188 509252 640252
rect 252140 640052 252204 640116
rect 302004 640112 302068 640116
rect 302004 640056 302054 640112
rect 302054 640056 302068 640112
rect 302004 640052 302068 640056
rect 326292 640052 326356 640116
rect 336412 640052 336476 640116
rect 231716 639916 231780 639980
rect 233004 639916 233068 639980
rect 239444 639916 239508 639980
rect 251772 639916 251836 639980
rect 257844 639916 257908 639980
rect 287100 639916 287164 639980
rect 297404 639916 297468 639980
rect 306604 639916 306668 639980
rect 316724 639916 316788 639980
rect 328132 639976 328196 639980
rect 328132 639920 328182 639976
rect 328182 639920 328196 639976
rect 328132 639916 328196 639920
rect 335308 639916 335372 639980
rect 345796 640052 345860 640116
rect 403572 640052 403636 640116
rect 413324 640052 413388 640116
rect 456748 640052 456812 640116
rect 345612 639916 345676 639980
rect 372292 639916 372356 639980
rect 384252 639916 384316 639980
rect 393084 639916 393148 639980
rect 441660 639916 441724 639980
rect 451964 639916 452028 639980
rect 5396 639780 5460 639844
rect 234476 639780 234540 639844
rect 235580 639780 235644 639844
rect 249380 639780 249444 639844
rect 255636 639780 255700 639844
rect 267780 639780 267844 639844
rect 282316 639780 282380 639844
rect 32996 639508 33060 639572
rect 33180 639508 33244 639572
rect 33180 639372 33244 639436
rect 32996 639236 33060 639300
rect 235580 639508 235644 639572
rect 249012 639508 249076 639572
rect 239444 639372 239508 639436
rect 251772 639372 251836 639436
rect 249012 639236 249076 639300
rect 257844 639372 257908 639436
rect 267780 639372 267844 639436
rect 282316 639372 282380 639436
rect 287100 639372 287164 639436
rect 297404 639372 297468 639436
rect 306604 639372 306668 639436
rect 316724 639372 316788 639436
rect 326292 639372 326356 639436
rect 335308 639372 335372 639436
rect 336412 639372 336476 639436
rect 345612 639372 345676 639436
rect 345796 639372 345860 639436
rect 372292 639372 372356 639436
rect 384252 639372 384316 639436
rect 393084 639372 393148 639436
rect 403572 639372 403636 639436
rect 413324 639372 413388 639436
rect 441660 639372 441724 639436
rect 493364 639644 493428 639708
rect 509188 639644 509252 639708
rect 527404 639644 527468 639708
rect 451964 639372 452028 639436
rect 456748 639372 456812 639436
rect 252140 639236 252204 639300
rect 493364 639100 493428 639164
rect 509188 638964 509252 639028
rect 328132 638556 328196 638620
rect 302004 638420 302068 638484
rect 255636 638284 255700 638348
rect 434484 638148 434548 638212
rect 526116 637740 526180 637804
rect 527220 637740 527284 637804
rect 527220 634340 527284 634404
rect 527588 634340 527652 634404
rect 527404 634204 527468 634268
rect 527220 633932 527284 633996
rect 527588 630668 527652 630732
rect 527404 630532 527468 630596
rect 527772 627812 527836 627876
rect 528508 627812 528572 627876
rect 527220 623052 527284 623116
rect 528140 623052 528204 623116
rect 527588 618292 527652 618356
rect 528508 618292 528572 618356
rect 528140 618156 528204 618220
rect 528692 618156 528756 618220
rect 527220 618020 527284 618084
rect 527588 618020 527652 618084
rect 527220 608636 527284 608700
rect 527956 608636 528020 608700
rect 528324 608636 528388 608700
rect 528692 608636 528756 608700
rect 527588 603740 527652 603804
rect 528324 603740 528388 603804
rect 527220 587148 527284 587212
rect 527956 587148 528020 587212
rect 527404 579804 527468 579868
rect 527956 579532 528020 579596
rect 528324 579532 528388 579596
rect 528324 570148 528388 570212
rect 527772 570012 527836 570076
rect 527772 563076 527836 563140
rect 527956 562804 528020 562868
rect 527404 560220 527468 560284
rect 527956 560220 528020 560284
rect 527404 550836 527468 550900
rect 527772 550700 527836 550764
rect 527772 543900 527836 543964
rect 527220 543492 527284 543556
rect 527220 533972 527284 534036
rect 528140 533972 528204 534036
rect 528140 524588 528204 524652
rect 527956 524180 528020 524244
rect 527220 521596 527284 521660
rect 527956 521596 528020 521660
rect 527220 512212 527284 512276
rect 527588 512076 527652 512140
rect 527588 505140 527652 505204
rect 527772 504868 527836 504932
rect 527404 502284 527468 502348
rect 527772 502284 527836 502348
rect 527404 492628 527468 492692
rect 527956 492628 528020 492692
rect 527956 485828 528020 485892
rect 527772 485556 527836 485620
rect 527772 482836 527836 482900
rect 528140 482836 528204 482900
rect 527588 473316 527652 473380
rect 528140 473316 528204 473380
rect 527220 466244 527284 466308
rect 527588 466244 527652 466308
rect 527220 456724 527284 456788
rect 527772 456724 527836 456788
rect 527220 444348 527284 444412
rect 527588 444348 527652 444412
rect 527220 437412 527284 437476
rect 527956 437412 528020 437476
rect 527956 427892 528020 427956
rect 527772 427620 527836 427684
rect 527772 424900 527836 424964
rect 527404 424764 527468 424828
rect 527404 415380 527468 415444
rect 527956 415380 528020 415444
rect 527956 408580 528020 408644
rect 527772 408308 527836 408372
rect 527220 405588 527284 405652
rect 527772 405588 527836 405652
rect 527220 396068 527284 396132
rect 527588 396068 527652 396132
rect 527588 389268 527652 389332
rect 527404 388996 527468 389060
rect 527404 386276 527468 386340
rect 527956 386140 528020 386204
rect 527588 376756 527652 376820
rect 527956 376756 528020 376820
rect 527588 369956 527652 370020
rect 527772 369684 527836 369748
rect 527772 366964 527836 367028
rect 528324 366828 528388 366892
rect 527956 357444 528020 357508
rect 528324 357444 528388 357508
rect 527956 350644 528020 350708
rect 527772 350372 527836 350436
rect 527772 347652 527836 347716
rect 528324 347652 528388 347716
rect 527588 340308 527652 340372
rect 528324 340308 528388 340372
rect 527588 336636 527652 336700
rect 332732 328400 332796 328404
rect 332732 328344 332746 328400
rect 332746 328344 332796 328400
rect 332732 328340 332796 328344
rect 332732 318956 332796 319020
rect 527404 318820 527468 318884
rect 527404 312020 527468 312084
rect 527588 311748 527652 311812
rect 233004 309028 233068 309092
rect 527588 309088 527652 309092
rect 527588 309032 527638 309088
rect 527638 309032 527652 309088
rect 527588 309028 527652 309032
rect 249380 307668 249444 307732
rect 527404 302092 527468 302156
rect 249196 298148 249260 298212
rect 249196 289852 249260 289916
rect 527588 289776 527652 289780
rect 527588 289720 527638 289776
rect 527638 289720 527652 289776
rect 527588 289716 527652 289720
rect 249564 289580 249628 289644
rect 527404 280196 527468 280260
rect 249196 279848 249260 279852
rect 249196 279792 249246 279848
rect 249246 279792 249260 279848
rect 249196 279788 249260 279792
rect 527404 273396 527468 273460
rect 527588 272988 527652 273052
rect 249380 270540 249444 270604
rect 249380 270404 249444 270468
rect 527588 270404 527652 270468
rect 527404 260884 527468 260948
rect 249564 260612 249628 260676
rect 527404 253948 527468 254012
rect 527588 253676 527652 253740
rect 232820 252452 232884 252516
rect 249380 251092 249444 251156
rect 527588 251092 527652 251156
rect 249196 241572 249260 241636
rect 527404 241572 527468 241636
rect 527404 234636 527468 234700
rect 527588 234364 527652 234428
rect 249196 231916 249260 231980
rect 249380 231916 249444 231980
rect 527588 231840 527652 231844
rect 527588 231784 527638 231840
rect 527638 231784 527652 231840
rect 527588 231780 527652 231784
rect 249380 222260 249444 222324
rect 527772 222260 527836 222324
rect 527772 215460 527836 215524
rect 527588 215188 527652 215252
rect 249380 214568 249444 214572
rect 249380 214512 249430 214568
rect 249430 214512 249444 214568
rect 249380 214508 249444 214512
rect 527588 212468 527652 212532
rect 232636 208252 232700 208316
rect 527404 202948 527468 203012
rect 249564 199956 249628 200020
rect 527404 196012 527468 196076
rect 527588 195740 527652 195804
rect 527588 193156 527652 193220
rect 249564 185600 249628 185604
rect 249564 185544 249578 185600
rect 249578 185544 249628 185600
rect 249564 185540 249628 185544
rect 527404 183636 527468 183700
rect 249564 179344 249628 179348
rect 249564 179288 249614 179344
rect 249614 179288 249628 179344
rect 249564 179284 249628 179288
rect 527404 176700 527468 176764
rect 527220 176428 527284 176492
rect 527220 173904 527284 173908
rect 527220 173848 527270 173904
rect 527270 173848 527284 173904
rect 527220 173844 527284 173848
rect 550588 170444 550652 170508
rect 233740 170308 233804 170372
rect 248644 170308 248708 170372
rect 376708 170308 376772 170372
rect 248460 170036 248524 170100
rect 376708 170036 376772 170100
rect 249564 169764 249628 169828
rect 550588 170172 550652 170236
rect 249564 167044 249628 167108
rect 249564 166908 249628 166972
rect 232452 165548 232516 165612
rect 527404 164188 527468 164252
rect 370084 157584 370148 157588
rect 370084 157528 370098 157584
rect 370098 157528 370148 157584
rect 370084 157524 370148 157528
rect 527404 157388 527468 157452
rect 527220 157116 527284 157180
rect 249748 154532 249812 154596
rect 249748 154396 249812 154460
rect 370084 154592 370148 154596
rect 370084 154536 370098 154592
rect 370098 154536 370148 154592
rect 370084 154532 370148 154536
rect 527220 154396 527284 154460
rect 249380 144876 249444 144940
rect 249748 144876 249812 144940
rect 527404 144876 527468 144940
rect 527404 139980 527468 140044
rect 527772 139980 527836 140044
rect 370084 138272 370148 138276
rect 370084 138216 370134 138272
rect 370134 138216 370148 138272
rect 370084 138212 370148 138216
rect 370084 135280 370148 135284
rect 370084 135224 370098 135280
rect 370098 135224 370148 135280
rect 370084 135220 370148 135224
rect 527772 135144 527836 135148
rect 527772 135088 527822 135144
rect 527822 135088 527836 135144
rect 527772 135084 527836 135088
rect 376708 134540 376772 134604
rect 304948 134404 305012 134468
rect 367140 134268 367204 134332
rect 376708 134268 376772 134332
rect 315988 134132 316052 134196
rect 249380 133860 249444 133924
rect 357388 133996 357452 134060
rect 367140 133996 367204 134060
rect 315988 133860 316052 133924
rect 343588 133860 343652 133924
rect 304948 133724 305012 133788
rect 453988 133996 454052 134060
rect 473308 133996 473372 134060
rect 502196 134132 502260 134196
rect 453988 133724 454052 133788
rect 343588 133588 343652 133652
rect 357204 133588 357268 133652
rect 473308 133588 473372 133652
rect 502196 133860 502260 133924
rect 531268 133996 531332 134060
rect 550588 133996 550652 134060
rect 531268 133588 531332 133652
rect 550588 133724 550652 133788
rect 527404 125564 527468 125628
rect 527404 118764 527468 118828
rect 527588 118492 527652 118556
rect 527220 108972 527284 109036
rect 527772 108972 527836 109036
rect 527772 99452 527836 99516
rect 527588 99180 527652 99244
rect 527588 96460 527652 96524
rect 527404 87000 527468 87004
rect 527404 86944 527454 87000
rect 527454 86944 527468 87000
rect 527404 86940 527468 86944
rect 527404 80140 527468 80204
rect 527220 79868 527284 79932
rect 243124 77420 243188 77484
rect 243124 75984 243188 75988
rect 243124 75928 243138 75984
rect 243138 75928 243188 75984
rect 243124 75924 243188 75928
rect 527220 70484 527284 70548
rect 527588 70212 527652 70276
rect 527220 62732 527284 62796
rect 527772 62732 527836 62796
rect 527220 57836 527284 57900
rect 527404 48316 527468 48380
rect 527404 41516 527468 41580
rect 527588 41244 527652 41308
rect 373948 40624 374012 40628
rect 373948 40568 373962 40624
rect 373962 40568 374012 40624
rect 373948 40564 374012 40568
rect 354628 40428 354692 40492
rect 335308 40292 335372 40356
rect 373948 40292 374012 40356
rect 234476 40020 234540 40084
rect 335308 40080 335372 40084
rect 354628 40156 354692 40220
rect 335308 40024 335322 40080
rect 335322 40024 335372 40080
rect 335308 40020 335372 40024
rect 502196 40292 502260 40356
rect 502196 40020 502260 40084
rect 531268 40156 531332 40220
rect 550588 40156 550652 40220
rect 531268 39748 531332 39812
rect 550588 39884 550652 39948
rect 527588 38524 527652 38588
rect 527404 29004 527468 29068
rect 527404 22204 527468 22268
rect 550588 17308 550652 17372
rect 259500 17172 259564 17236
rect 325740 17172 325804 17236
rect 531268 17172 531332 17236
rect 231716 16764 231780 16828
rect 259500 16900 259564 16964
rect 325740 16900 325804 16964
rect 357388 16900 357452 16964
rect 299428 16628 299492 16692
rect 357572 16628 357636 16692
rect 365668 16628 365732 16692
rect 502012 17036 502076 17100
rect 531268 16900 531332 16964
rect 502196 16628 502260 16692
rect 550588 17036 550652 17100
rect 395844 16492 395908 16556
rect 396028 16492 396092 16556
rect 299428 16356 299492 16420
rect 365668 16356 365732 16420
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 5398 639845 5458 641462
rect 5395 639844 5461 639845
rect 5395 639780 5396 639844
rect 5460 639780 5461 639844
rect 5395 639779 5461 639780
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 12939 641612 13005 641613
rect 12939 641548 12940 641612
rect 13004 641548 13005 641612
rect 12939 641547 13005 641548
rect 12942 641018 13002 641547
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 607254 30204 642698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 32995 639572 33061 639573
rect 32995 639508 32996 639572
rect 33060 639508 33061 639572
rect 32995 639507 33061 639508
rect 33179 639572 33245 639573
rect 33179 639508 33180 639572
rect 33244 639508 33245 639572
rect 33179 639507 33245 639508
rect 32998 639301 33058 639507
rect 33182 639437 33242 639507
rect 33179 639436 33245 639437
rect 33179 639372 33180 639436
rect 33244 639372 33245 639436
rect 33179 639371 33245 639372
rect 32995 639300 33061 639301
rect 32995 639236 32996 639300
rect 33060 639236 33061 639300
rect 32995 639235 33061 639236
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 621654 80604 657098
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 80838 640933 80898 641462
rect 80835 640932 80901 640933
rect 80835 640868 80836 640932
rect 80900 640868 80901 640932
rect 80835 640867 80901 640868
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 614454 109404 649898
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 109723 641612 109789 641613
rect 109723 641548 109724 641612
rect 109788 641548 109789 641612
rect 109723 641547 109789 641548
rect 109726 641018 109786 641547
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 607254 138204 642698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 138430 640933 138490 641462
rect 138427 640932 138493 640933
rect 138427 640868 138428 640932
rect 138492 640868 138493 640932
rect 138427 640867 138493 640868
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 636054 167004 671498
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 167315 641612 167381 641613
rect 167315 641548 167316 641612
rect 167380 641548 167381 641612
rect 167315 641547 167381 641548
rect 167318 641018 167378 641547
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 621654 224604 657098
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 226011 641612 226077 641613
rect 226011 641548 226012 641612
rect 226076 641548 226077 641612
rect 226011 641547 226077 641548
rect 226014 641018 226074 641547
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 625254 228204 660698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 233739 642972 233805 642973
rect 233739 642908 233740 642972
rect 233804 642908 233805 642972
rect 233739 642907 233805 642908
rect 232819 642700 232885 642701
rect 232819 642636 232820 642700
rect 232884 642636 232885 642700
rect 232819 642635 232885 642636
rect 232635 642564 232701 642565
rect 232635 642500 232636 642564
rect 232700 642500 232701 642564
rect 232635 642499 232701 642500
rect 232451 642428 232517 642429
rect 232451 642364 232452 642428
rect 232516 642364 232517 642428
rect 232451 642363 232517 642364
rect 231899 641612 231965 641613
rect 231899 641548 231900 641612
rect 231964 641548 231965 641612
rect 231899 641547 231965 641548
rect 231902 641018 231962 641547
rect 231715 639980 231781 639981
rect 231715 639916 231716 639980
rect 231780 639916 231781 639980
rect 231715 639915 231781 639916
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 231718 16829 231778 639915
rect 232454 165613 232514 642363
rect 232638 208317 232698 642499
rect 232822 252517 232882 642635
rect 233003 639980 233069 639981
rect 233003 639916 233004 639980
rect 233068 639916 233069 639980
rect 233003 639915 233069 639916
rect 233006 309093 233066 639915
rect 233003 309092 233069 309093
rect 233003 309028 233004 309092
rect 233068 309028 233069 309092
rect 233003 309027 233069 309028
rect 232819 252516 232885 252517
rect 232819 252452 232820 252516
rect 232884 252452 232885 252516
rect 232819 252451 232885 252452
rect 232635 208316 232701 208317
rect 232635 208252 232636 208316
rect 232700 208252 232701 208316
rect 232635 208251 232701 208252
rect 233742 170373 233802 642907
rect 234475 639844 234541 639845
rect 234475 639780 234476 639844
rect 234540 639780 234541 639844
rect 234475 639779 234541 639780
rect 233739 170372 233805 170373
rect 233739 170308 233740 170372
rect 233804 170308 233805 170372
rect 233739 170307 233805 170308
rect 232451 165612 232517 165613
rect 232451 165548 232452 165612
rect 232516 165548 232517 165612
rect 232451 165547 232517 165548
rect 234478 40085 234538 639779
rect 234804 632454 235404 667898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 235579 639844 235645 639845
rect 235579 639780 235580 639844
rect 235644 639780 235645 639844
rect 235579 639779 235645 639780
rect 235582 639573 235642 639779
rect 235579 639572 235645 639573
rect 235579 639508 235580 639572
rect 235644 639508 235645 639572
rect 235579 639507 235645 639508
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234475 40084 234541 40085
rect 234475 40020 234476 40084
rect 234540 40020 234541 40084
rect 234475 40019 234541 40020
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 231715 16828 231781 16829
rect 231715 16764 231716 16828
rect 231780 16764 231781 16828
rect 231715 16763 231781 16764
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 636054 239004 671498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 239443 639980 239509 639981
rect 239443 639916 239444 639980
rect 239508 639916 239509 639980
rect 239443 639915 239509 639916
rect 239446 639437 239506 639915
rect 242004 639654 242604 675098
rect 239443 639436 239509 639437
rect 239443 639372 239444 639436
rect 239508 639372 239509 639436
rect 239443 639371 239509 639372
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252139 640116 252205 640117
rect 252139 640052 252140 640116
rect 252204 640052 252205 640116
rect 252139 640051 252205 640052
rect 251771 639980 251837 639981
rect 251771 639916 251772 639980
rect 251836 639916 251837 639980
rect 251771 639915 251837 639916
rect 249379 639844 249445 639845
rect 249379 639780 249380 639844
rect 249444 639780 249445 639844
rect 249379 639779 249445 639780
rect 249011 639572 249077 639573
rect 249011 639508 249012 639572
rect 249076 639508 249077 639572
rect 249011 639507 249077 639508
rect 249014 639301 249074 639507
rect 249011 639300 249077 639301
rect 249011 639236 249012 639300
rect 249076 639236 249077 639300
rect 249011 639235 249077 639236
rect 249382 630730 249442 639779
rect 251774 639437 251834 639915
rect 251771 639436 251837 639437
rect 251771 639372 251772 639436
rect 251836 639372 251837 639436
rect 251771 639371 251837 639372
rect 252142 639301 252202 640051
rect 252139 639300 252205 639301
rect 252139 639236 252140 639300
rect 252204 639236 252205 639300
rect 252139 639235 252205 639236
rect 249382 630670 249626 630730
rect 249566 630138 249626 630670
rect 249382 625290 249442 627182
rect 249382 625230 249626 625290
rect 249566 617810 249626 625230
rect 249382 617750 249626 617810
rect 249382 615858 249442 617750
rect 249566 613050 249626 614942
rect 249530 612990 249626 613050
rect 252804 614454 253404 649898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 255635 639844 255701 639845
rect 255635 639780 255636 639844
rect 255700 639780 255701 639844
rect 255635 639779 255701 639780
rect 255638 638349 255698 639779
rect 255635 638348 255701 638349
rect 255635 638284 255636 638348
rect 255700 638284 255701 638348
rect 255635 638283 255701 638284
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 249198 608290 249258 608822
rect 249198 608230 249442 608290
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 249382 369610 249442 608230
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 249382 369550 249626 369610
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 249566 347850 249626 369550
rect 249382 347790 249626 347850
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 249382 343090 249442 347790
rect 249382 343030 249626 343090
rect 249566 342498 249626 343030
rect 249198 332210 249258 341582
rect 249198 332150 249442 332210
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 249382 307733 249442 332150
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 249379 307732 249445 307733
rect 249379 307668 249380 307732
rect 249444 307668 249445 307732
rect 249379 307667 249445 307668
rect 249195 298212 249261 298213
rect 249195 298148 249196 298212
rect 249260 298148 249261 298212
rect 249195 298147 249261 298148
rect 249198 289917 249258 298147
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 249195 289916 249261 289917
rect 249195 289852 249196 289916
rect 249260 289852 249261 289916
rect 249195 289851 249261 289852
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 249563 289644 249629 289645
rect 249563 289580 249564 289644
rect 249628 289580 249629 289644
rect 249563 289579 249629 289580
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 249566 281890 249626 289579
rect 249198 281830 249626 281890
rect 249198 279853 249258 281830
rect 249195 279852 249261 279853
rect 249195 279788 249196 279852
rect 249260 279788 249261 279852
rect 249195 279787 249261 279788
rect 249379 270604 249445 270605
rect 249379 270540 249380 270604
rect 249444 270540 249445 270604
rect 249379 270539 249445 270540
rect 249382 270469 249442 270539
rect 249379 270468 249445 270469
rect 249379 270404 249380 270468
rect 249444 270404 249445 270468
rect 249379 270403 249445 270404
rect 249563 260676 249629 260677
rect 249563 260612 249564 260676
rect 249628 260612 249629 260676
rect 249563 260611 249629 260612
rect 249566 251290 249626 260611
rect 249382 251230 249626 251290
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 249382 251157 249442 251230
rect 249379 251156 249445 251157
rect 249379 251092 249380 251156
rect 249444 251092 249445 251156
rect 249379 251091 249445 251092
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 249195 241636 249261 241637
rect 249195 241572 249196 241636
rect 249260 241572 249261 241636
rect 249195 241571 249261 241572
rect 249198 231981 249258 241571
rect 249195 231980 249261 231981
rect 249195 231916 249196 231980
rect 249260 231916 249261 231980
rect 249195 231915 249261 231916
rect 249379 231980 249445 231981
rect 249379 231916 249380 231980
rect 249444 231916 249445 231980
rect 249379 231915 249445 231916
rect 249382 222325 249442 231915
rect 249379 222324 249445 222325
rect 249379 222260 249380 222324
rect 249444 222260 249445 222324
rect 249379 222259 249445 222260
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 249379 214572 249445 214573
rect 249379 214508 249380 214572
rect 249444 214508 249445 214572
rect 249379 214507 249445 214508
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 249382 206410 249442 214507
rect 249382 206350 249626 206410
rect 249566 200021 249626 206350
rect 249563 200020 249629 200021
rect 249563 199956 249564 200020
rect 249628 199956 249629 200020
rect 249563 199955 249629 199956
rect 249563 185604 249629 185605
rect 249563 185540 249564 185604
rect 249628 185540 249629 185604
rect 249563 185539 249629 185540
rect 249566 179349 249626 185539
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 249563 179348 249629 179349
rect 249563 179284 249564 179348
rect 249628 179284 249629 179348
rect 249563 179283 249629 179284
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 248643 170372 248709 170373
rect 248643 170308 248644 170372
rect 248708 170308 248709 170372
rect 248643 170307 248709 170308
rect 248459 170100 248525 170101
rect 248459 170036 248460 170100
rect 248524 170098 248525 170100
rect 248646 170098 248706 170307
rect 248524 170038 248706 170098
rect 248524 170036 248525 170038
rect 248459 170035 248525 170036
rect 249563 169828 249629 169829
rect 249563 169764 249564 169828
rect 249628 169764 249629 169828
rect 249563 169763 249629 169764
rect 249566 167109 249626 169763
rect 249563 167108 249629 167109
rect 249563 167044 249564 167108
rect 249628 167044 249629 167108
rect 249563 167043 249629 167044
rect 249563 166972 249629 166973
rect 249563 166908 249564 166972
rect 249628 166908 249629 166972
rect 249563 166907 249629 166908
rect 249566 160850 249626 166907
rect 249566 160790 249810 160850
rect 249750 154597 249810 160790
rect 249747 154596 249813 154597
rect 249747 154532 249748 154596
rect 249812 154532 249813 154596
rect 249747 154531 249813 154532
rect 249747 154460 249813 154461
rect 249747 154396 249748 154460
rect 249812 154396 249813 154460
rect 249747 154395 249813 154396
rect 249750 144941 249810 154395
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 249379 144940 249445 144941
rect 249379 144876 249380 144940
rect 249444 144876 249445 144940
rect 249379 144875 249445 144876
rect 249747 144940 249813 144941
rect 249747 144876 249748 144940
rect 249812 144876 249813 144940
rect 249747 144875 249813 144876
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 249382 133925 249442 144875
rect 249379 133924 249445 133925
rect 249379 133860 249380 133924
rect 249444 133860 249445 133924
rect 249379 133859 249445 133860
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 243123 77484 243189 77485
rect 243123 77420 243124 77484
rect 243188 77420 243189 77484
rect 243123 77419 243189 77420
rect 243126 75989 243186 77419
rect 243123 75988 243189 75989
rect 243123 75924 243124 75988
rect 243188 75924 243189 75988
rect 243123 75923 243189 75924
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 618054 257004 653498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 257843 639980 257909 639981
rect 257843 639916 257844 639980
rect 257908 639916 257909 639980
rect 257843 639915 257909 639916
rect 257846 639437 257906 639915
rect 257843 639436 257909 639437
rect 257843 639372 257844 639436
rect 257908 639372 257909 639436
rect 257843 639371 257909 639372
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 259499 17236 259565 17237
rect 259499 17172 259500 17236
rect 259564 17172 259565 17236
rect 259499 17171 259565 17172
rect 259502 16965 259562 17171
rect 259499 16964 259565 16965
rect 259499 16900 259500 16964
rect 259564 16900 259565 16964
rect 259499 16899 259565 16900
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 264470 640933 264530 641462
rect 264467 640932 264533 640933
rect 264467 640868 264468 640932
rect 264532 640868 264533 640932
rect 264467 640867 264533 640868
rect 267779 639844 267845 639845
rect 267779 639780 267780 639844
rect 267844 639780 267845 639844
rect 267779 639779 267845 639780
rect 267782 639437 267842 639779
rect 267779 639436 267845 639437
rect 267779 639372 267780 639436
rect 267844 639372 267845 639436
rect 267779 639371 267845 639372
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 287099 639980 287165 639981
rect 287099 639916 287100 639980
rect 287164 639916 287165 639980
rect 287099 639915 287165 639916
rect 282315 639844 282381 639845
rect 282315 639780 282316 639844
rect 282380 639780 282381 639844
rect 282315 639779 282381 639780
rect 282318 639437 282378 639779
rect 287102 639437 287162 639915
rect 282315 639436 282381 639437
rect 282315 639372 282316 639436
rect 282380 639372 282381 639436
rect 282315 639371 282381 639372
rect 287099 639436 287165 639437
rect 287099 639372 287100 639436
rect 287164 639372 287165 639436
rect 287099 639371 287165 639372
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 614454 289404 649898
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299246 640933 299306 641462
rect 299243 640932 299309 640933
rect 299243 640868 299244 640932
rect 299308 640868 299309 640932
rect 299243 640867 299309 640868
rect 297403 639980 297469 639981
rect 297403 639916 297404 639980
rect 297468 639916 297469 639980
rect 297403 639915 297469 639916
rect 297406 639437 297466 639915
rect 297403 639436 297469 639437
rect 297403 639372 297404 639436
rect 297468 639372 297469 639436
rect 297403 639371 297469 639372
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 299604 625254 300204 660698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 302003 640116 302069 640117
rect 302003 640052 302004 640116
rect 302068 640052 302069 640116
rect 302003 640051 302069 640052
rect 302006 638485 302066 640051
rect 306603 639980 306669 639981
rect 306603 639916 306604 639980
rect 306668 639916 306669 639980
rect 306603 639915 306669 639916
rect 306606 639437 306666 639915
rect 306603 639436 306669 639437
rect 306603 639372 306604 639436
rect 306668 639372 306669 639436
rect 306603 639371 306669 639372
rect 302003 638484 302069 638485
rect 302003 638420 302004 638484
rect 302068 638420 302069 638484
rect 302003 638419 302069 638420
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 306804 632454 307404 667898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 304947 134468 305013 134469
rect 304947 134404 304948 134468
rect 305012 134404 305013 134468
rect 304947 134403 305013 134404
rect 304950 133789 305010 134403
rect 304947 133788 305013 133789
rect 304947 133724 304948 133788
rect 305012 133724 305013 133788
rect 304947 133723 305013 133724
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299427 16692 299493 16693
rect 299427 16628 299428 16692
rect 299492 16628 299493 16692
rect 299427 16627 299493 16628
rect 299430 16421 299490 16627
rect 299427 16420 299493 16421
rect 299427 16356 299428 16420
rect 299492 16356 299493 16420
rect 299427 16355 299493 16356
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 316723 639980 316789 639981
rect 316723 639916 316724 639980
rect 316788 639916 316789 639980
rect 316723 639915 316789 639916
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 316726 639437 316786 639915
rect 314004 639334 314604 639418
rect 316723 639436 316789 639437
rect 316723 639372 316724 639436
rect 316788 639372 316789 639436
rect 316723 639371 316789 639372
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 317604 607254 318204 642698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 318379 641612 318445 641613
rect 318379 641548 318380 641612
rect 318444 641548 318445 641612
rect 318379 641547 318445 641548
rect 318382 641018 318442 641547
rect 322062 640933 322122 641462
rect 322059 640932 322125 640933
rect 322059 640868 322060 640932
rect 322124 640868 322125 640932
rect 322059 640867 322125 640868
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 315987 134196 316053 134197
rect 315987 134132 315988 134196
rect 316052 134132 316053 134196
rect 315987 134131 316053 134132
rect 315990 133925 316050 134131
rect 315987 133924 316053 133925
rect 315987 133860 315988 133924
rect 316052 133860 316053 133924
rect 315987 133859 316053 133860
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 614454 325404 649898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 326291 640116 326357 640117
rect 326291 640052 326292 640116
rect 326356 640052 326357 640116
rect 326291 640051 326357 640052
rect 326294 639437 326354 640051
rect 328131 639980 328197 639981
rect 328131 639916 328132 639980
rect 328196 639916 328197 639980
rect 328131 639915 328197 639916
rect 326291 639436 326357 639437
rect 326291 639372 326292 639436
rect 326356 639372 326357 639436
rect 326291 639371 326357 639372
rect 328134 638621 328194 639915
rect 328131 638620 328197 638621
rect 328131 638556 328132 638620
rect 328196 638556 328197 638620
rect 328131 638555 328197 638556
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 325739 17236 325805 17237
rect 325739 17172 325740 17236
rect 325804 17172 325805 17236
rect 325739 17171 325805 17172
rect 325742 16965 325802 17171
rect 325739 16964 325805 16965
rect 325739 16900 325740 16964
rect 325804 16900 325805 16964
rect 325739 16899 325805 16900
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335307 639980 335373 639981
rect 335307 639916 335308 639980
rect 335372 639916 335373 639980
rect 335307 639915 335373 639916
rect 335310 639437 335370 639915
rect 335307 639436 335373 639437
rect 335307 639372 335308 639436
rect 335372 639372 335373 639436
rect 335307 639371 335373 639372
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 335604 625254 336204 660698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 336595 641612 336661 641613
rect 336595 641548 336596 641612
rect 336660 641548 336661 641612
rect 336595 641547 336661 641548
rect 336598 641018 336658 641547
rect 336411 640116 336477 640117
rect 336411 640052 336412 640116
rect 336476 640052 336477 640116
rect 336411 640051 336477 640052
rect 336414 639437 336474 640051
rect 336411 639436 336477 639437
rect 336411 639372 336412 639436
rect 336476 639372 336477 639436
rect 336411 639371 336477 639372
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 332731 328404 332797 328405
rect 332731 328340 332732 328404
rect 332796 328340 332797 328404
rect 332731 328339 332797 328340
rect 332734 319021 332794 328339
rect 332731 319020 332797 319021
rect 332731 318956 332732 319020
rect 332796 318956 332797 319020
rect 332731 318955 332797 318956
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335307 40356 335373 40357
rect 335307 40292 335308 40356
rect 335372 40292 335373 40356
rect 335307 40291 335373 40292
rect 335310 40085 335370 40291
rect 335307 40084 335373 40085
rect 335307 40020 335308 40084
rect 335372 40020 335373 40084
rect 335307 40019 335373 40020
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 632454 343404 667898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 345795 640116 345861 640117
rect 345795 640052 345796 640116
rect 345860 640052 345861 640116
rect 345795 640051 345861 640052
rect 345611 639980 345677 639981
rect 345611 639916 345612 639980
rect 345676 639916 345677 639980
rect 345611 639915 345677 639916
rect 345614 639437 345674 639915
rect 345798 639437 345858 640051
rect 345611 639436 345677 639437
rect 345611 639372 345612 639436
rect 345676 639372 345677 639436
rect 345611 639371 345677 639372
rect 345795 639436 345861 639437
rect 345795 639372 345796 639436
rect 345860 639372 345861 639436
rect 345795 639371 345861 639372
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 346404 636054 347004 671498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 343587 133924 343653 133925
rect 343587 133860 343588 133924
rect 343652 133860 343653 133924
rect 343587 133859 343653 133860
rect 343590 133653 343650 133859
rect 343587 133652 343653 133653
rect 343587 133588 343588 133652
rect 343652 133588 343653 133652
rect 343587 133587 343653 133588
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 639654 350604 675098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 351131 641612 351197 641613
rect 351131 641548 351132 641612
rect 351196 641548 351197 641612
rect 351131 641547 351197 641548
rect 351134 641018 351194 641547
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 607254 354204 642698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 357387 134060 357453 134061
rect 357387 133996 357388 134060
rect 357452 133996 357453 134060
rect 357387 133995 357453 133996
rect 357203 133652 357269 133653
rect 357203 133588 357204 133652
rect 357268 133650 357269 133652
rect 357390 133650 357450 133995
rect 357268 133590 357450 133650
rect 357268 133588 357269 133590
rect 357203 133587 357269 133588
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 354627 40492 354693 40493
rect 354627 40428 354628 40492
rect 354692 40428 354693 40492
rect 354627 40427 354693 40428
rect 354630 40221 354690 40427
rect 354627 40220 354693 40221
rect 354627 40156 354628 40220
rect 354692 40156 354693 40220
rect 354627 40155 354693 40156
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 357387 16964 357453 16965
rect 357387 16900 357388 16964
rect 357452 16900 357453 16964
rect 357387 16899 357453 16900
rect 357390 16690 357450 16899
rect 357571 16692 357637 16693
rect 357571 16690 357572 16692
rect 357390 16630 357572 16690
rect 357571 16628 357572 16630
rect 357636 16628 357637 16692
rect 357571 16627 357637 16628
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 366958 641550 367202 641610
rect 366958 640933 367018 641550
rect 367142 640933 367202 641550
rect 366955 640932 367021 640933
rect 366955 640868 366956 640932
rect 367020 640868 367021 640932
rect 366955 640867 367021 640868
rect 367139 640932 367205 640933
rect 367139 640868 367140 640932
rect 367204 640868 367205 640932
rect 367139 640867 367205 640868
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 372291 639980 372357 639981
rect 372291 639916 372292 639980
rect 372356 639916 372357 639980
rect 372291 639915 372357 639916
rect 372294 639437 372354 639915
rect 372291 639436 372357 639437
rect 372291 639372 372292 639436
rect 372356 639372 372357 639436
rect 372291 639371 372357 639372
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 370083 157588 370149 157589
rect 370083 157524 370084 157588
rect 370148 157524 370149 157588
rect 370083 157523 370149 157524
rect 370086 154597 370146 157523
rect 371604 157254 372204 192698
rect 378804 632454 379404 667898
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 379651 641612 379717 641613
rect 379651 641548 379652 641612
rect 379716 641548 379717 641612
rect 379651 641547 379717 641548
rect 379654 641018 379714 641547
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 376707 170372 376773 170373
rect 376707 170308 376708 170372
rect 376772 170308 376773 170372
rect 376707 170307 376773 170308
rect 376710 170101 376770 170307
rect 376707 170100 376773 170101
rect 376707 170036 376708 170100
rect 376772 170036 376773 170100
rect 376707 170035 376773 170036
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 370083 154596 370149 154597
rect 370083 154532 370084 154596
rect 370148 154532 370149 154596
rect 370083 154531 370149 154532
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 367139 134332 367205 134333
rect 367139 134268 367140 134332
rect 367204 134268 367205 134332
rect 367139 134267 367205 134268
rect 367142 134061 367202 134267
rect 367139 134060 367205 134061
rect 367139 133996 367140 134060
rect 367204 133996 367205 134060
rect 367139 133995 367205 133996
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 368004 117654 368604 153098
rect 370083 138276 370149 138277
rect 370083 138212 370084 138276
rect 370148 138212 370149 138276
rect 370083 138211 370149 138212
rect 370086 135285 370146 138211
rect 370083 135284 370149 135285
rect 370083 135220 370084 135284
rect 370148 135220 370149 135284
rect 370083 135219 370149 135220
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 365667 16692 365733 16693
rect 365667 16628 365668 16692
rect 365732 16628 365733 16692
rect 365667 16627 365733 16628
rect 365670 16421 365730 16627
rect 365667 16420 365733 16421
rect 365667 16356 365668 16420
rect 365732 16356 365733 16420
rect 365667 16355 365733 16356
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 121254 372204 156698
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 376707 134604 376773 134605
rect 376707 134540 376708 134604
rect 376772 134540 376773 134604
rect 376707 134539 376773 134540
rect 376710 134333 376770 134539
rect 376707 134332 376773 134333
rect 376707 134268 376708 134332
rect 376772 134268 376773 134332
rect 376707 134267 376773 134268
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 373947 40628 374013 40629
rect 373947 40564 373948 40628
rect 374012 40564 374013 40628
rect 373947 40563 374013 40564
rect 373950 40357 374010 40563
rect 373947 40356 374013 40357
rect 373947 40292 373948 40356
rect 374012 40292 374013 40356
rect 373947 40291 374013 40292
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 636054 383004 671498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 384251 639980 384317 639981
rect 384251 639916 384252 639980
rect 384316 639916 384317 639980
rect 384251 639915 384317 639916
rect 384254 639437 384314 639915
rect 386004 639654 386604 675098
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 384251 639436 384317 639437
rect 384251 639372 384252 639436
rect 384316 639372 384317 639436
rect 384251 639371 384317 639372
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 607254 390204 642698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 393083 639980 393149 639981
rect 393083 639916 393084 639980
rect 393148 639916 393149 639980
rect 393083 639915 393149 639916
rect 393086 639437 393146 639915
rect 393083 639436 393149 639437
rect 393083 639372 393084 639436
rect 393148 639372 393149 639436
rect 393083 639371 393149 639372
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 614454 397404 649898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 395846 16630 396090 16690
rect 395846 16557 395906 16630
rect 396030 16557 396090 16630
rect 395843 16556 395909 16557
rect 395843 16492 395844 16556
rect 395908 16492 395909 16556
rect 395843 16491 395909 16492
rect 396027 16556 396093 16557
rect 396027 16492 396028 16556
rect 396092 16492 396093 16556
rect 396027 16491 396093 16492
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 618054 401004 653498
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 403571 640116 403637 640117
rect 403571 640052 403572 640116
rect 403636 640052 403637 640116
rect 403571 640051 403637 640052
rect 403574 639437 403634 640051
rect 403571 639436 403637 639437
rect 403571 639372 403572 639436
rect 403636 639372 403637 639436
rect 403571 639371 403637 639372
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 413323 640116 413389 640117
rect 413323 640052 413324 640116
rect 413388 640052 413389 640116
rect 413323 640051 413389 640052
rect 413326 639437 413386 640051
rect 413323 639436 413389 639437
rect 413323 639372 413324 639436
rect 413388 639372 413389 639436
rect 413323 639371 413389 639372
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 607254 426204 642698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432459 641612 432525 641613
rect 432459 641548 432460 641612
rect 432524 641548 432525 641612
rect 432459 641547 432525 641548
rect 432462 641018 432522 641547
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 614454 433404 649898
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 434483 642156 434549 642157
rect 434483 642092 434484 642156
rect 434548 642092 434549 642156
rect 434483 642091 434549 642092
rect 434486 638213 434546 642091
rect 434483 638212 434549 638213
rect 434483 638148 434484 638212
rect 434548 638148 434549 638212
rect 434483 638147 434549 638148
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 618054 437004 653498
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 438534 640933 438594 641462
rect 438531 640932 438597 640933
rect 438531 640868 438532 640932
rect 438596 640868 438597 640932
rect 438531 640867 438597 640868
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 621654 440604 657098
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 441659 639980 441725 639981
rect 441659 639916 441660 639980
rect 441724 639916 441725 639980
rect 441659 639915 441725 639916
rect 441662 639437 441722 639915
rect 441659 639436 441725 639437
rect 441659 639372 441660 639436
rect 441724 639372 441725 639436
rect 441659 639371 441725 639372
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 451963 639980 452029 639981
rect 451963 639916 451964 639980
rect 452028 639916 452029 639980
rect 451963 639915 452029 639916
rect 451966 639437 452026 639915
rect 451963 639436 452029 639437
rect 451963 639372 451964 639436
rect 452028 639372 452029 639436
rect 451963 639371 452029 639372
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 454404 636054 455004 671498
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 456747 640116 456813 640117
rect 456747 640052 456748 640116
rect 456812 640052 456813 640116
rect 456747 640051 456813 640052
rect 456750 639437 456810 640051
rect 458004 639654 458604 675098
rect 456747 639436 456813 639437
rect 456747 639372 456748 639436
rect 456812 639372 456813 639436
rect 456747 639371 456813 639372
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 453987 134060 454053 134061
rect 453987 133996 453988 134060
rect 454052 133996 454053 134060
rect 453987 133995 454053 133996
rect 453990 133789 454050 133995
rect 453987 133788 454053 133789
rect 453987 133724 453988 133788
rect 454052 133724 454053 133788
rect 453987 133723 454053 133724
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 463555 641612 463621 641613
rect 463555 641548 463556 641612
rect 463620 641548 463621 641612
rect 463555 641547 463621 641548
rect 463558 641018 463618 641547
rect 463926 640253 463986 640782
rect 463923 640252 463989 640253
rect 463923 640188 463924 640252
rect 463988 640188 463989 640252
rect 463923 640187 463989 640188
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 473307 134060 473373 134061
rect 473307 133996 473308 134060
rect 473372 133996 473373 134060
rect 473307 133995 473373 133996
rect 473310 133653 473370 133995
rect 473307 133652 473373 133653
rect 473307 133588 473308 133652
rect 473372 133588 473373 133652
rect 473307 133587 473373 133588
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 480854 640253 480914 641462
rect 480851 640252 480917 640253
rect 480851 640188 480852 640252
rect 480916 640188 480917 640252
rect 480851 640187 480917 640188
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 493363 639708 493429 639709
rect 493363 639644 493364 639708
rect 493428 639644 493429 639708
rect 493363 639643 493429 639644
rect 494004 639654 494604 675098
rect 493366 639165 493426 639643
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 493363 639164 493429 639165
rect 493363 639100 493364 639164
rect 493428 639100 493429 639164
rect 493363 639099 493429 639100
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 502195 134196 502261 134197
rect 502195 134132 502196 134196
rect 502260 134132 502261 134196
rect 502195 134131 502261 134132
rect 502198 133925 502258 134131
rect 502195 133924 502261 133925
rect 502195 133860 502196 133924
rect 502260 133860 502261 133924
rect 502195 133859 502261 133860
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 502195 40356 502261 40357
rect 502195 40292 502196 40356
rect 502260 40292 502261 40356
rect 502195 40291 502261 40292
rect 502198 40085 502258 40291
rect 502195 40084 502261 40085
rect 502195 40020 502196 40084
rect 502260 40020 502261 40084
rect 502195 40019 502261 40020
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 502011 17100 502077 17101
rect 502011 17036 502012 17100
rect 502076 17036 502077 17100
rect 502011 17035 502077 17036
rect 502014 16690 502074 17035
rect 502195 16692 502261 16693
rect 502195 16690 502196 16692
rect 502014 16630 502196 16690
rect 502195 16628 502196 16630
rect 502260 16628 502261 16692
rect 502195 16627 502261 16628
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 509187 639708 509253 639709
rect 509187 639644 509188 639708
rect 509252 639644 509253 639708
rect 509187 639643 509253 639644
rect 509190 639029 509250 639643
rect 509187 639028 509253 639029
rect 509187 638964 509188 639028
rect 509252 638964 509253 639028
rect 509187 638963 509253 638964
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526115 642972 526181 642973
rect 526115 642908 526116 642972
rect 526180 642908 526181 642972
rect 526115 642907 526181 642908
rect 526118 637805 526178 642907
rect 526115 637804 526181 637805
rect 526115 637740 526116 637804
rect 526180 637740 526181 637804
rect 526115 637739 526181 637740
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 636054 527004 671498
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 527403 639708 527469 639709
rect 527403 639644 527404 639708
rect 527468 639644 527469 639708
rect 527403 639643 527469 639644
rect 530004 639654 530604 675098
rect 527219 637804 527285 637805
rect 527219 637740 527220 637804
rect 527284 637740 527285 637804
rect 527219 637739 527285 637740
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 527222 634405 527282 637739
rect 527219 634404 527285 634405
rect 527219 634340 527220 634404
rect 527284 634340 527285 634404
rect 527219 634339 527285 634340
rect 527406 634269 527466 639643
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 527587 634404 527653 634405
rect 527587 634340 527588 634404
rect 527652 634340 527653 634404
rect 527587 634339 527653 634340
rect 527403 634268 527469 634269
rect 527403 634204 527404 634268
rect 527468 634204 527469 634268
rect 527403 634203 527469 634204
rect 527219 633996 527285 633997
rect 527219 633932 527220 633996
rect 527284 633932 527285 633996
rect 527219 633931 527285 633932
rect 527222 623117 527282 633931
rect 527590 630733 527650 634339
rect 527587 630732 527653 630733
rect 527587 630668 527588 630732
rect 527652 630668 527653 630732
rect 527587 630667 527653 630668
rect 527403 630596 527469 630597
rect 527403 630532 527404 630596
rect 527468 630532 527469 630596
rect 527403 630531 527469 630532
rect 527406 628010 527466 630531
rect 527406 627950 527834 628010
rect 527774 627877 527834 627950
rect 527771 627876 527837 627877
rect 527771 627812 527772 627876
rect 527836 627812 527837 627876
rect 527771 627811 527837 627812
rect 528507 627876 528573 627877
rect 528507 627812 528508 627876
rect 528572 627812 528573 627876
rect 528507 627811 528573 627812
rect 527219 623116 527285 623117
rect 527219 623052 527220 623116
rect 527284 623052 527285 623116
rect 527219 623051 527285 623052
rect 528139 623116 528205 623117
rect 528139 623052 528140 623116
rect 528204 623052 528205 623116
rect 528139 623051 528205 623052
rect 527587 618356 527653 618357
rect 527587 618292 527588 618356
rect 527652 618292 527653 618356
rect 527587 618291 527653 618292
rect 527590 618085 527650 618291
rect 528142 618221 528202 623051
rect 528510 618357 528570 627811
rect 528507 618356 528573 618357
rect 528507 618292 528508 618356
rect 528572 618292 528573 618356
rect 528507 618291 528573 618292
rect 528139 618220 528205 618221
rect 528139 618156 528140 618220
rect 528204 618156 528205 618220
rect 528139 618155 528205 618156
rect 528691 618220 528757 618221
rect 528691 618156 528692 618220
rect 528756 618156 528757 618220
rect 528691 618155 528757 618156
rect 527219 618084 527285 618085
rect 527219 618020 527220 618084
rect 527284 618020 527285 618084
rect 527219 618019 527285 618020
rect 527587 618084 527653 618085
rect 527587 618020 527588 618084
rect 527652 618020 527653 618084
rect 527587 618019 527653 618020
rect 527222 608701 527282 618019
rect 528694 608701 528754 618155
rect 527219 608700 527285 608701
rect 527219 608636 527220 608700
rect 527284 608636 527285 608700
rect 527219 608635 527285 608636
rect 527955 608700 528021 608701
rect 527955 608636 527956 608700
rect 528020 608636 528021 608700
rect 527955 608635 528021 608636
rect 528323 608700 528389 608701
rect 528323 608636 528324 608700
rect 528388 608636 528389 608700
rect 528323 608635 528389 608636
rect 528691 608700 528757 608701
rect 528691 608636 528692 608700
rect 528756 608636 528757 608700
rect 528691 608635 528757 608636
rect 527587 603804 527653 603805
rect 527587 603740 527588 603804
rect 527652 603740 527653 603804
rect 527587 603739 527653 603740
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 527590 596050 527650 603739
rect 527222 595990 527650 596050
rect 527222 587213 527282 595990
rect 527958 589250 528018 608635
rect 528326 603805 528386 608635
rect 528323 603804 528389 603805
rect 528323 603740 528324 603804
rect 528388 603740 528389 603804
rect 528323 603739 528389 603740
rect 527590 589190 528018 589250
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 527219 587212 527285 587213
rect 527219 587148 527220 587212
rect 527284 587148 527285 587212
rect 527219 587147 527285 587148
rect 527590 582450 527650 589190
rect 527955 587212 528021 587213
rect 527955 587148 527956 587212
rect 528020 587148 528021 587212
rect 527955 587147 528021 587148
rect 527406 582390 527650 582450
rect 527406 579869 527466 582390
rect 527403 579868 527469 579869
rect 527403 579804 527404 579868
rect 527468 579804 527469 579868
rect 527403 579803 527469 579804
rect 527958 579597 528018 587147
rect 527955 579596 528021 579597
rect 527955 579532 527956 579596
rect 528020 579532 528021 579596
rect 527955 579531 528021 579532
rect 528323 579596 528389 579597
rect 528323 579532 528324 579596
rect 528388 579532 528389 579596
rect 528323 579531 528389 579532
rect 528326 570213 528386 579531
rect 528323 570212 528389 570213
rect 528323 570148 528324 570212
rect 528388 570148 528389 570212
rect 528323 570147 528389 570148
rect 527771 570076 527837 570077
rect 527771 570012 527772 570076
rect 527836 570012 527837 570076
rect 527771 570011 527837 570012
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 527774 563141 527834 570011
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 527771 563140 527837 563141
rect 527771 563076 527772 563140
rect 527836 563076 527837 563140
rect 527771 563075 527837 563076
rect 527955 562868 528021 562869
rect 527955 562804 527956 562868
rect 528020 562804 528021 562868
rect 527955 562803 528021 562804
rect 527958 560285 528018 562803
rect 527403 560284 527469 560285
rect 527403 560220 527404 560284
rect 527468 560220 527469 560284
rect 527403 560219 527469 560220
rect 527955 560284 528021 560285
rect 527955 560220 527956 560284
rect 528020 560220 528021 560284
rect 527955 560219 528021 560220
rect 527406 550901 527466 560219
rect 527403 550900 527469 550901
rect 527403 550836 527404 550900
rect 527468 550836 527469 550900
rect 527403 550835 527469 550836
rect 527771 550764 527837 550765
rect 527771 550700 527772 550764
rect 527836 550700 527837 550764
rect 527771 550699 527837 550700
rect 527774 543965 527834 550699
rect 527771 543964 527837 543965
rect 527771 543900 527772 543964
rect 527836 543900 527837 543964
rect 527771 543899 527837 543900
rect 527219 543556 527285 543557
rect 527219 543492 527220 543556
rect 527284 543492 527285 543556
rect 527219 543491 527285 543492
rect 527222 534037 527282 543491
rect 527219 534036 527285 534037
rect 527219 533972 527220 534036
rect 527284 533972 527285 534036
rect 527219 533971 527285 533972
rect 528139 534036 528205 534037
rect 528139 533972 528140 534036
rect 528204 533972 528205 534036
rect 528139 533971 528205 533972
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 528142 524653 528202 533971
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 528139 524652 528205 524653
rect 528139 524588 528140 524652
rect 528204 524588 528205 524652
rect 528139 524587 528205 524588
rect 527955 524244 528021 524245
rect 527955 524180 527956 524244
rect 528020 524180 528021 524244
rect 527955 524179 528021 524180
rect 527958 521661 528018 524179
rect 527219 521660 527285 521661
rect 527219 521596 527220 521660
rect 527284 521596 527285 521660
rect 527219 521595 527285 521596
rect 527955 521660 528021 521661
rect 527955 521596 527956 521660
rect 528020 521596 528021 521660
rect 527955 521595 528021 521596
rect 527222 512277 527282 521595
rect 527219 512276 527285 512277
rect 527219 512212 527220 512276
rect 527284 512212 527285 512276
rect 527219 512211 527285 512212
rect 527587 512140 527653 512141
rect 527587 512076 527588 512140
rect 527652 512076 527653 512140
rect 527587 512075 527653 512076
rect 527590 505205 527650 512075
rect 527587 505204 527653 505205
rect 527587 505140 527588 505204
rect 527652 505140 527653 505204
rect 527587 505139 527653 505140
rect 527771 504932 527837 504933
rect 527771 504868 527772 504932
rect 527836 504868 527837 504932
rect 527771 504867 527837 504868
rect 527774 502349 527834 504867
rect 527403 502348 527469 502349
rect 527403 502284 527404 502348
rect 527468 502284 527469 502348
rect 527403 502283 527469 502284
rect 527771 502348 527837 502349
rect 527771 502284 527772 502348
rect 527836 502284 527837 502348
rect 527771 502283 527837 502284
rect 527406 492693 527466 502283
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 527403 492692 527469 492693
rect 527403 492628 527404 492692
rect 527468 492628 527469 492692
rect 527403 492627 527469 492628
rect 527955 492692 528021 492693
rect 527955 492628 527956 492692
rect 528020 492628 528021 492692
rect 527955 492627 528021 492628
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 527958 485893 528018 492627
rect 527955 485892 528021 485893
rect 527955 485828 527956 485892
rect 528020 485828 528021 485892
rect 527955 485827 528021 485828
rect 527771 485620 527837 485621
rect 527771 485556 527772 485620
rect 527836 485556 527837 485620
rect 527771 485555 527837 485556
rect 527774 482901 527834 485555
rect 527771 482900 527837 482901
rect 527771 482836 527772 482900
rect 527836 482836 527837 482900
rect 527771 482835 527837 482836
rect 528139 482900 528205 482901
rect 528139 482836 528140 482900
rect 528204 482836 528205 482900
rect 528139 482835 528205 482836
rect 528142 473381 528202 482835
rect 527587 473380 527653 473381
rect 527587 473316 527588 473380
rect 527652 473316 527653 473380
rect 527587 473315 527653 473316
rect 528139 473380 528205 473381
rect 528139 473316 528140 473380
rect 528204 473316 528205 473380
rect 528139 473315 528205 473316
rect 527590 466309 527650 473315
rect 527219 466308 527285 466309
rect 527219 466244 527220 466308
rect 527284 466244 527285 466308
rect 527219 466243 527285 466244
rect 527587 466308 527653 466309
rect 527587 466244 527588 466308
rect 527652 466244 527653 466308
rect 527587 466243 527653 466244
rect 527222 456789 527282 466243
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 527219 456788 527285 456789
rect 527219 456724 527220 456788
rect 527284 456724 527285 456788
rect 527219 456723 527285 456724
rect 527771 456788 527837 456789
rect 527771 456724 527772 456788
rect 527836 456724 527837 456788
rect 527771 456723 527837 456724
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 527774 453930 527834 456723
rect 527590 453870 527834 453930
rect 527590 444413 527650 453870
rect 527219 444412 527285 444413
rect 527219 444348 527220 444412
rect 527284 444348 527285 444412
rect 527219 444347 527285 444348
rect 527587 444412 527653 444413
rect 527587 444348 527588 444412
rect 527652 444348 527653 444412
rect 527587 444347 527653 444348
rect 527222 437477 527282 444347
rect 527219 437476 527285 437477
rect 527219 437412 527220 437476
rect 527284 437412 527285 437476
rect 527219 437411 527285 437412
rect 527955 437476 528021 437477
rect 527955 437412 527956 437476
rect 528020 437412 528021 437476
rect 527955 437411 528021 437412
rect 527958 427957 528018 437411
rect 527955 427956 528021 427957
rect 527955 427892 527956 427956
rect 528020 427892 528021 427956
rect 527955 427891 528021 427892
rect 527771 427684 527837 427685
rect 527771 427620 527772 427684
rect 527836 427620 527837 427684
rect 527771 427619 527837 427620
rect 527774 424965 527834 427619
rect 527771 424964 527837 424965
rect 527771 424900 527772 424964
rect 527836 424900 527837 424964
rect 527771 424899 527837 424900
rect 527403 424828 527469 424829
rect 527403 424764 527404 424828
rect 527468 424764 527469 424828
rect 527403 424763 527469 424764
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 527406 415445 527466 424763
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 527403 415444 527469 415445
rect 527403 415380 527404 415444
rect 527468 415380 527469 415444
rect 527403 415379 527469 415380
rect 527955 415444 528021 415445
rect 527955 415380 527956 415444
rect 528020 415380 528021 415444
rect 527955 415379 528021 415380
rect 527958 408645 528018 415379
rect 527955 408644 528021 408645
rect 527955 408580 527956 408644
rect 528020 408580 528021 408644
rect 527955 408579 528021 408580
rect 527771 408372 527837 408373
rect 527771 408308 527772 408372
rect 527836 408308 527837 408372
rect 527771 408307 527837 408308
rect 527774 405653 527834 408307
rect 527219 405652 527285 405653
rect 527219 405588 527220 405652
rect 527284 405588 527285 405652
rect 527219 405587 527285 405588
rect 527771 405652 527837 405653
rect 527771 405588 527772 405652
rect 527836 405588 527837 405652
rect 527771 405587 527837 405588
rect 527222 396133 527282 405587
rect 527219 396132 527285 396133
rect 527219 396068 527220 396132
rect 527284 396068 527285 396132
rect 527219 396067 527285 396068
rect 527587 396132 527653 396133
rect 527587 396068 527588 396132
rect 527652 396068 527653 396132
rect 527587 396067 527653 396068
rect 527590 389333 527650 396067
rect 527587 389332 527653 389333
rect 527587 389268 527588 389332
rect 527652 389268 527653 389332
rect 527587 389267 527653 389268
rect 527403 389060 527469 389061
rect 527403 388996 527404 389060
rect 527468 388996 527469 389060
rect 527403 388995 527469 388996
rect 527406 386341 527466 388995
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 527403 386340 527469 386341
rect 527403 386276 527404 386340
rect 527468 386276 527469 386340
rect 527403 386275 527469 386276
rect 527955 386204 528021 386205
rect 527955 386140 527956 386204
rect 528020 386140 528021 386204
rect 527955 386139 528021 386140
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 527958 376821 528018 386139
rect 527587 376820 527653 376821
rect 527587 376756 527588 376820
rect 527652 376756 527653 376820
rect 527587 376755 527653 376756
rect 527955 376820 528021 376821
rect 527955 376756 527956 376820
rect 528020 376756 528021 376820
rect 527955 376755 528021 376756
rect 527590 370021 527650 376755
rect 527587 370020 527653 370021
rect 527587 369956 527588 370020
rect 527652 369956 527653 370020
rect 527587 369955 527653 369956
rect 527771 369748 527837 369749
rect 527771 369684 527772 369748
rect 527836 369684 527837 369748
rect 527771 369683 527837 369684
rect 527774 367029 527834 369683
rect 527771 367028 527837 367029
rect 527771 366964 527772 367028
rect 527836 366964 527837 367028
rect 527771 366963 527837 366964
rect 528323 366892 528389 366893
rect 528323 366828 528324 366892
rect 528388 366828 528389 366892
rect 528323 366827 528389 366828
rect 528326 357509 528386 366827
rect 527955 357508 528021 357509
rect 527955 357444 527956 357508
rect 528020 357444 528021 357508
rect 527955 357443 528021 357444
rect 528323 357508 528389 357509
rect 528323 357444 528324 357508
rect 528388 357444 528389 357508
rect 528323 357443 528389 357444
rect 527958 350709 528018 357443
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 527955 350708 528021 350709
rect 527955 350644 527956 350708
rect 528020 350644 528021 350708
rect 527955 350643 528021 350644
rect 527771 350436 527837 350437
rect 527771 350372 527772 350436
rect 527836 350372 527837 350436
rect 527771 350371 527837 350372
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 527774 347717 527834 350371
rect 527771 347716 527837 347717
rect 527771 347652 527772 347716
rect 527836 347652 527837 347716
rect 527771 347651 527837 347652
rect 528323 347716 528389 347717
rect 528323 347652 528324 347716
rect 528388 347652 528389 347716
rect 528323 347651 528389 347652
rect 526404 312054 527004 347498
rect 528326 340373 528386 347651
rect 527587 340372 527653 340373
rect 527587 340308 527588 340372
rect 527652 340308 527653 340372
rect 527587 340307 527653 340308
rect 528323 340372 528389 340373
rect 528323 340308 528324 340372
rect 528388 340308 528389 340372
rect 528323 340307 528389 340308
rect 527590 336701 527650 340307
rect 527587 336700 527653 336701
rect 527587 336636 527588 336700
rect 527652 336636 527653 336700
rect 527587 336635 527653 336636
rect 527403 318884 527469 318885
rect 527403 318820 527404 318884
rect 527468 318820 527469 318884
rect 527403 318819 527469 318820
rect 527406 312085 527466 318819
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 527403 312084 527469 312085
rect 527403 312020 527404 312084
rect 527468 312020 527469 312084
rect 527403 312019 527469 312020
rect 526404 311734 527004 311818
rect 527587 311812 527653 311813
rect 527587 311748 527588 311812
rect 527652 311748 527653 311812
rect 527587 311747 527653 311748
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 527590 309093 527650 311747
rect 527587 309092 527653 309093
rect 527587 309028 527588 309092
rect 527652 309028 527653 309092
rect 527587 309027 527653 309028
rect 527403 302156 527469 302157
rect 527403 302092 527404 302156
rect 527468 302092 527469 302156
rect 527403 302091 527469 302092
rect 527406 292770 527466 302091
rect 527406 292710 527650 292770
rect 527590 289781 527650 292710
rect 527587 289780 527653 289781
rect 527587 289716 527588 289780
rect 527652 289716 527653 289780
rect 527587 289715 527653 289716
rect 527403 280260 527469 280261
rect 527403 280196 527404 280260
rect 527468 280196 527469 280260
rect 527403 280195 527469 280196
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 527406 273461 527466 280195
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 527403 273460 527469 273461
rect 527403 273396 527404 273460
rect 527468 273396 527469 273460
rect 527403 273395 527469 273396
rect 527587 273052 527653 273053
rect 527587 272988 527588 273052
rect 527652 272988 527653 273052
rect 527587 272987 527653 272988
rect 527590 270469 527650 272987
rect 527587 270468 527653 270469
rect 527587 270404 527588 270468
rect 527652 270404 527653 270468
rect 527587 270403 527653 270404
rect 527403 260948 527469 260949
rect 527403 260884 527404 260948
rect 527468 260884 527469 260948
rect 527403 260883 527469 260884
rect 527406 254013 527466 260883
rect 527403 254012 527469 254013
rect 527403 253948 527404 254012
rect 527468 253948 527469 254012
rect 527403 253947 527469 253948
rect 527587 253740 527653 253741
rect 527587 253676 527588 253740
rect 527652 253676 527653 253740
rect 527587 253675 527653 253676
rect 527590 251157 527650 253675
rect 527587 251156 527653 251157
rect 527587 251092 527588 251156
rect 527652 251092 527653 251156
rect 527587 251091 527653 251092
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 527403 241636 527469 241637
rect 527403 241572 527404 241636
rect 527468 241572 527469 241636
rect 527403 241571 527469 241572
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 527406 234701 527466 241571
rect 527403 234700 527469 234701
rect 527403 234636 527404 234700
rect 527468 234636 527469 234700
rect 527403 234635 527469 234636
rect 527587 234428 527653 234429
rect 527587 234364 527588 234428
rect 527652 234364 527653 234428
rect 527587 234363 527653 234364
rect 527590 231845 527650 234363
rect 527587 231844 527653 231845
rect 527587 231780 527588 231844
rect 527652 231780 527653 231844
rect 527587 231779 527653 231780
rect 527771 222324 527837 222325
rect 527771 222260 527772 222324
rect 527836 222260 527837 222324
rect 527771 222259 527837 222260
rect 527774 215525 527834 222259
rect 527771 215524 527837 215525
rect 527771 215460 527772 215524
rect 527836 215460 527837 215524
rect 527771 215459 527837 215460
rect 527587 215252 527653 215253
rect 527587 215188 527588 215252
rect 527652 215188 527653 215252
rect 527587 215187 527653 215188
rect 527590 212533 527650 215187
rect 527587 212532 527653 212533
rect 527587 212468 527588 212532
rect 527652 212468 527653 212532
rect 527587 212467 527653 212468
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 527403 203012 527469 203013
rect 527403 202948 527404 203012
rect 527468 202948 527469 203012
rect 527403 202947 527469 202948
rect 527406 196077 527466 202947
rect 527403 196076 527469 196077
rect 527403 196012 527404 196076
rect 527468 196012 527469 196076
rect 527403 196011 527469 196012
rect 527587 195804 527653 195805
rect 527587 195740 527588 195804
rect 527652 195740 527653 195804
rect 527587 195739 527653 195740
rect 527590 193221 527650 195739
rect 527587 193220 527653 193221
rect 527587 193156 527588 193220
rect 527652 193156 527653 193220
rect 527587 193155 527653 193156
rect 527403 183700 527469 183701
rect 527403 183636 527404 183700
rect 527468 183636 527469 183700
rect 527403 183635 527469 183636
rect 527406 176765 527466 183635
rect 527403 176764 527469 176765
rect 527403 176700 527404 176764
rect 527468 176700 527469 176764
rect 527403 176699 527469 176700
rect 527219 176492 527285 176493
rect 527219 176428 527220 176492
rect 527284 176428 527285 176492
rect 527219 176427 527285 176428
rect 527222 173909 527282 176427
rect 527219 173908 527285 173909
rect 527219 173844 527220 173908
rect 527284 173844 527285 173908
rect 527219 173843 527285 173844
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 527403 164252 527469 164253
rect 527403 164188 527404 164252
rect 527468 164188 527469 164252
rect 527403 164187 527469 164188
rect 527406 157453 527466 164187
rect 527403 157452 527469 157453
rect 527403 157388 527404 157452
rect 527468 157388 527469 157452
rect 527403 157387 527469 157388
rect 527219 157180 527285 157181
rect 527219 157116 527220 157180
rect 527284 157116 527285 157180
rect 527219 157115 527285 157116
rect 527222 154461 527282 157115
rect 527219 154460 527285 154461
rect 527219 154396 527220 154460
rect 527284 154396 527285 154460
rect 527219 154395 527285 154396
rect 527403 144940 527469 144941
rect 527403 144876 527404 144940
rect 527468 144876 527469 144940
rect 527403 144875 527469 144876
rect 527406 140045 527466 144875
rect 527403 140044 527469 140045
rect 527403 139980 527404 140044
rect 527468 139980 527469 140044
rect 527403 139979 527469 139980
rect 527771 140044 527837 140045
rect 527771 139980 527772 140044
rect 527836 139980 527837 140044
rect 527771 139979 527837 139980
rect 527774 135149 527834 139979
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 527771 135148 527837 135149
rect 527771 135084 527772 135148
rect 527836 135084 527837 135148
rect 527771 135083 527837 135084
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 527403 125628 527469 125629
rect 527403 125564 527404 125628
rect 527468 125564 527469 125628
rect 527403 125563 527469 125564
rect 527406 118829 527466 125563
rect 527403 118828 527469 118829
rect 527403 118764 527404 118828
rect 527468 118764 527469 118828
rect 527403 118763 527469 118764
rect 527587 118556 527653 118557
rect 527587 118492 527588 118556
rect 527652 118492 527653 118556
rect 527587 118491 527653 118492
rect 527590 109170 527650 118491
rect 527222 109110 527650 109170
rect 527222 109037 527282 109110
rect 527219 109036 527285 109037
rect 527219 108972 527220 109036
rect 527284 108972 527285 109036
rect 527219 108971 527285 108972
rect 527771 109036 527837 109037
rect 527771 108972 527772 109036
rect 527836 108972 527837 109036
rect 527771 108971 527837 108972
rect 527774 99517 527834 108971
rect 530004 99654 530604 135098
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 531267 134060 531333 134061
rect 531267 133996 531268 134060
rect 531332 133996 531333 134060
rect 531267 133995 531333 133996
rect 531270 133653 531330 133995
rect 531267 133652 531333 133653
rect 531267 133588 531268 133652
rect 531332 133588 531333 133652
rect 531267 133587 531333 133588
rect 527771 99516 527837 99517
rect 527771 99452 527772 99516
rect 527836 99452 527837 99516
rect 527771 99451 527837 99452
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 527587 99244 527653 99245
rect 527587 99180 527588 99244
rect 527652 99180 527653 99244
rect 527587 99179 527653 99180
rect 527590 96525 527650 99179
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 527587 96524 527653 96525
rect 527587 96460 527588 96524
rect 527652 96460 527653 96524
rect 527587 96459 527653 96460
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 527403 87004 527469 87005
rect 527403 86940 527404 87004
rect 527468 86940 527469 87004
rect 527403 86939 527469 86940
rect 527406 80205 527466 86939
rect 527403 80204 527469 80205
rect 527403 80140 527404 80204
rect 527468 80140 527469 80204
rect 527403 80139 527469 80140
rect 527219 79932 527285 79933
rect 527219 79868 527220 79932
rect 527284 79868 527285 79932
rect 527219 79867 527285 79868
rect 527222 70549 527282 79867
rect 527219 70548 527285 70549
rect 527219 70484 527220 70548
rect 527284 70484 527285 70548
rect 527219 70483 527285 70484
rect 527587 70276 527653 70277
rect 527587 70212 527588 70276
rect 527652 70212 527653 70276
rect 527587 70211 527653 70212
rect 527590 67690 527650 70211
rect 527590 67630 527834 67690
rect 527774 62797 527834 67630
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 527219 62796 527285 62797
rect 527219 62732 527220 62796
rect 527284 62732 527285 62796
rect 527219 62731 527285 62732
rect 527771 62796 527837 62797
rect 527771 62732 527772 62796
rect 527836 62732 527837 62796
rect 527771 62731 527837 62732
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 527222 57901 527282 62731
rect 527219 57900 527285 57901
rect 527219 57836 527220 57900
rect 527284 57836 527285 57900
rect 527219 57835 527285 57836
rect 527403 48380 527469 48381
rect 527403 48316 527404 48380
rect 527468 48316 527469 48380
rect 527403 48315 527469 48316
rect 527406 41581 527466 48315
rect 527403 41580 527469 41581
rect 527403 41516 527404 41580
rect 527468 41516 527469 41580
rect 527403 41515 527469 41516
rect 527587 41308 527653 41309
rect 527587 41244 527588 41308
rect 527652 41244 527653 41308
rect 527587 41243 527653 41244
rect 527590 38589 527650 41243
rect 527587 38588 527653 38589
rect 527587 38524 527588 38588
rect 527652 38524 527653 38588
rect 527587 38523 527653 38524
rect 527403 29068 527469 29069
rect 527403 29004 527404 29068
rect 527468 29004 527469 29068
rect 527403 29003 527469 29004
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 527406 22269 527466 29003
rect 530004 27654 530604 63098
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 531267 40220 531333 40221
rect 531267 40156 531268 40220
rect 531332 40156 531333 40220
rect 531267 40155 531333 40156
rect 531270 39813 531330 40155
rect 531267 39812 531333 39813
rect 531267 39748 531268 39812
rect 531332 39748 531333 39812
rect 531267 39747 531333 39748
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 527403 22268 527469 22269
rect 527403 22204 527404 22268
rect 527468 22204 527469 22268
rect 527403 22203 527469 22204
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 -4946 530604 27098
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 531267 17236 531333 17237
rect 531267 17172 531268 17236
rect 531332 17172 531333 17236
rect 531267 17171 531333 17172
rect 531270 16965 531330 17171
rect 531267 16964 531333 16965
rect 531267 16900 531268 16964
rect 531332 16900 531333 16964
rect 531267 16899 531333 16900
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 550587 170508 550653 170509
rect 550587 170444 550588 170508
rect 550652 170444 550653 170508
rect 550587 170443 550653 170444
rect 550590 170237 550650 170443
rect 550587 170236 550653 170237
rect 550587 170172 550588 170236
rect 550652 170172 550653 170236
rect 550587 170171 550653 170172
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 550587 134060 550653 134061
rect 550587 133996 550588 134060
rect 550652 133996 550653 134060
rect 550587 133995 550653 133996
rect 550590 133789 550650 133995
rect 550587 133788 550653 133789
rect 550587 133724 550588 133788
rect 550652 133724 550653 133788
rect 550587 133723 550653 133724
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 550587 40220 550653 40221
rect 550587 40156 550588 40220
rect 550652 40156 550653 40220
rect 550587 40155 550653 40156
rect 550590 39949 550650 40155
rect 550587 39948 550653 39949
rect 550587 39884 550588 39948
rect 550652 39884 550653 39948
rect 550587 39883 550653 39884
rect 550587 17372 550653 17373
rect 550587 17308 550588 17372
rect 550652 17308 550653 17372
rect 550587 17307 550653 17308
rect 550590 17101 550650 17307
rect 550587 17100 550653 17101
rect 550587 17036 550588 17100
rect 550652 17036 550653 17100
rect 550587 17035 550653 17036
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 5310 641462 5546 641698
rect 7334 641612 7570 641698
rect 7334 641548 7420 641612
rect 7420 641548 7484 641612
rect 7484 641548 7570 641612
rect 7334 641462 7570 641548
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 12854 640782 13090 641018
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 27574 641612 27810 641698
rect 27574 641548 27660 641612
rect 27660 641548 27724 641612
rect 27724 641548 27810 641612
rect 27574 641462 27810 641548
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 79646 641612 79882 641698
rect 79646 641548 79732 641612
rect 79732 641548 79796 641612
rect 79796 641548 79882 641612
rect 79646 641462 79882 641548
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 80750 641462 80986 641698
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108350 640932 108586 641018
rect 108350 640868 108436 640932
rect 108436 640868 108500 640932
rect 108500 640868 108586 640932
rect 108350 640782 108586 640868
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 109638 640782 109874 641018
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137238 641612 137474 641698
rect 137238 641548 137324 641612
rect 137324 641548 137388 641612
rect 137388 641548 137474 641612
rect 137238 641462 137474 641548
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 138342 641462 138578 641698
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 165942 640932 166178 641018
rect 165942 640868 166028 640932
rect 166028 640868 166092 640932
rect 166092 640868 166178 640932
rect 165942 640782 166178 640868
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 167230 640782 167466 641018
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 215070 641612 215306 641698
rect 215070 641548 215156 641612
rect 215156 641548 215220 641612
rect 215220 641548 215306 641612
rect 215070 641462 215306 641548
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 222062 641612 222298 641698
rect 222062 641548 222148 641612
rect 222148 641548 222212 641612
rect 222212 641548 222298 641612
rect 222062 641462 222298 641548
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 225926 640782 226162 641018
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 231814 640782 232050 641018
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 251686 640932 251922 641018
rect 251686 640868 251772 640932
rect 251772 640868 251836 640932
rect 251836 640868 251922 640932
rect 251686 640782 251922 640868
rect 249478 629902 249714 630138
rect 249294 627182 249530 627418
rect 249294 615622 249530 615858
rect 249478 614942 249714 615178
rect 249294 612902 249530 613138
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 249110 608822 249346 609058
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 249478 342262 249714 342498
rect 249110 341582 249346 341818
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 264382 641462 264618 641698
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 282598 641612 282834 641698
rect 282598 641548 282684 641612
rect 282684 641548 282748 641612
rect 282748 641548 282834 641612
rect 282598 641462 282834 641548
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 289774 640932 290010 641018
rect 289774 640868 289860 640932
rect 289860 640868 289924 640932
rect 289924 640868 290010 640932
rect 289774 640782 290010 640868
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299158 641462 299394 641698
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 301550 641612 301786 641698
rect 301550 641548 301636 641612
rect 301636 641548 301700 641612
rect 301700 641548 301786 641612
rect 301550 641462 301786 641548
rect 302838 641612 303074 641698
rect 302838 641548 302924 641612
rect 302924 641548 302988 641612
rect 302988 641548 303074 641612
rect 302838 641462 303074 641548
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 309278 641612 309514 641698
rect 309278 641548 309364 641612
rect 309364 641548 309428 641612
rect 309428 641548 309514 641612
rect 309278 641462 309514 641548
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 321974 641462 322210 641698
rect 318294 640782 318530 641018
rect 318662 640932 318898 641018
rect 318662 640868 318748 640932
rect 318748 640868 318812 640932
rect 318812 640868 318898 640932
rect 318662 640782 318898 640868
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 326942 641612 327178 641698
rect 326942 641548 327028 641612
rect 327028 641548 327092 641612
rect 327092 641548 327178 641612
rect 326942 641462 327178 641548
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 336510 640782 336746 641018
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 348286 641612 348522 641698
rect 348286 641548 348372 641612
rect 348372 641548 348436 641612
rect 348436 641548 348522 641612
rect 348286 641462 348522 641548
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 351046 640782 351282 641018
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 357302 640932 357538 641018
rect 357302 640868 357388 640932
rect 357388 640868 357452 640932
rect 357452 640868 357538 640932
rect 357302 640782 357538 640868
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 376622 641612 376858 641698
rect 376622 641548 376708 641612
rect 376708 641548 376772 641612
rect 376772 641548 376858 641612
rect 376622 641462 376858 641548
rect 376438 640932 376674 641018
rect 376438 640868 376524 640932
rect 376524 640868 376588 640932
rect 376588 640868 376674 640932
rect 376438 640782 376674 640868
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 379566 640782 379802 641018
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 388950 640932 389186 641018
rect 388950 640868 389036 640932
rect 389036 640868 389100 640932
rect 389100 640868 389186 640932
rect 388950 640782 389186 640868
rect 386186 639418 386422 639654
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 395574 640932 395810 641018
rect 395574 640868 395660 640932
rect 395660 640868 395724 640932
rect 395724 640868 395810 640932
rect 395574 640782 395810 640868
rect 395942 640932 396178 641018
rect 395942 640868 396028 640932
rect 396028 640868 396092 640932
rect 396092 640868 396178 640932
rect 395942 640782 396178 640868
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 399254 640932 399490 641018
rect 399254 640868 399340 640932
rect 399340 640868 399404 640932
rect 399404 640868 399490 640932
rect 399254 640782 399490 640868
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 423542 641612 423778 641698
rect 423542 641548 423628 641612
rect 423628 641548 423692 641612
rect 423692 641548 423778 641612
rect 423542 641462 423778 641548
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432374 640782 432610 641018
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436054 640932 436290 641018
rect 436054 640868 436140 640932
rect 436140 640868 436204 640932
rect 436204 640868 436290 640932
rect 436054 640782 436290 640868
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 438446 641462 438682 641698
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 453902 641612 454138 641698
rect 453902 641548 453988 641612
rect 453988 641548 454052 641612
rect 454052 641548 454138 641612
rect 453902 641462 454138 641548
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 463470 640782 463706 641018
rect 463838 640782 464074 641018
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 480766 641462 481002 641698
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 509102 640252 509338 640338
rect 509102 640188 509188 640252
rect 509188 640188 509252 640252
rect 509252 640188 509338 640252
rect 509102 640102 509338 640188
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect 5268 641698 7612 641740
rect 5268 641462 5310 641698
rect 5546 641462 7334 641698
rect 7570 641462 7612 641698
rect 5268 641420 7612 641462
rect 19804 641698 27852 641740
rect 19804 641462 27574 641698
rect 27810 641462 27852 641698
rect 19804 641420 27852 641462
rect 79604 641698 81028 641740
rect 79604 641462 79646 641698
rect 79882 641462 80750 641698
rect 80986 641462 81028 641698
rect 79604 641420 81028 641462
rect 137196 641698 138620 641740
rect 137196 641462 137238 641698
rect 137474 641462 138342 641698
rect 138578 641462 138620 641698
rect 137196 641420 138620 641462
rect 215028 641698 222340 641740
rect 215028 641462 215070 641698
rect 215306 641462 222062 641698
rect 222298 641462 222340 641698
rect 215028 641420 222340 641462
rect 263052 641698 264660 641740
rect 263052 641462 264382 641698
rect 264618 641462 264660 641698
rect 263052 641420 264660 641462
rect 282400 641698 283060 641740
rect 282400 641462 282598 641698
rect 282834 641462 283060 641698
rect 282400 641420 283060 641462
rect 299116 641698 301828 641740
rect 299116 641462 299158 641698
rect 299394 641462 301550 641698
rect 301786 641462 301828 641698
rect 299116 641420 301828 641462
rect 302796 641698 309556 641740
rect 302796 641462 302838 641698
rect 303074 641462 309278 641698
rect 309514 641462 309556 641698
rect 302796 641420 309556 641462
rect 321932 641698 327220 641740
rect 321932 641462 321974 641698
rect 322210 641462 326942 641698
rect 327178 641462 327220 641698
rect 321932 641420 327220 641462
rect 340884 641698 348564 641740
rect 340884 641462 348286 641698
rect 348522 641462 348564 641698
rect 340884 641420 348564 641462
rect 376580 641698 376900 641740
rect 376580 641462 376622 641698
rect 376858 641462 376900 641698
rect 19804 641060 20124 641420
rect 263052 641060 263372 641420
rect 12812 641018 20124 641060
rect 12812 640782 12854 641018
rect 13090 640782 20124 641018
rect 12812 640740 20124 640782
rect 108308 641018 109916 641060
rect 108308 640782 108350 641018
rect 108586 640782 109638 641018
rect 109874 640782 109916 641018
rect 108308 640740 109916 640782
rect 165900 641018 167508 641060
rect 165900 640782 165942 641018
rect 166178 640782 167230 641018
rect 167466 640782 167508 641018
rect 165900 640740 167508 640782
rect 225884 641018 232092 641060
rect 225884 640782 225926 641018
rect 226162 640782 231814 641018
rect 232050 640782 232092 641018
rect 225884 640740 232092 640782
rect 251644 641018 263372 641060
rect 251644 640782 251686 641018
rect 251922 640782 263372 641018
rect 251644 640740 263372 640782
rect 282740 641060 283060 641420
rect 282740 641018 290052 641060
rect 282740 640782 289774 641018
rect 290010 640782 290052 641018
rect 282740 640740 290052 640782
rect 318252 641018 318940 641060
rect 318252 640782 318294 641018
rect 318530 640782 318662 641018
rect 318898 640782 318940 641018
rect 318252 640740 318940 640782
rect 336468 641018 340284 641060
rect 336468 640782 336510 641018
rect 336746 640782 340284 641018
rect 336468 640740 340284 640782
rect 339964 640380 340284 640740
rect 340884 640380 341204 641420
rect 376580 641060 376900 641462
rect 386148 641060 386652 641740
rect 417796 641698 423820 641740
rect 417796 641462 423542 641698
rect 423778 641462 423820 641698
rect 417796 641420 423820 641462
rect 438404 641698 444980 641740
rect 438404 641462 438446 641698
rect 438682 641462 444980 641698
rect 438404 641420 444980 641462
rect 417796 641060 418116 641420
rect 351004 641018 357580 641060
rect 351004 640782 351046 641018
rect 351282 640782 357302 641018
rect 357538 640782 357580 641018
rect 351004 640740 357580 640782
rect 376396 641018 376900 641060
rect 376396 640782 376438 641018
rect 376674 640782 376900 641018
rect 376396 640740 376900 640782
rect 379524 641018 389228 641060
rect 379524 640782 379566 641018
rect 379802 640782 388950 641018
rect 389186 640782 389228 641018
rect 379524 640740 389228 640782
rect 395532 641018 396220 641060
rect 395532 640782 395574 641018
rect 395810 640782 395942 641018
rect 396178 640782 396220 641018
rect 395532 640740 396220 640782
rect 399212 641018 418116 641060
rect 399212 640782 399254 641018
rect 399490 640782 418116 641018
rect 399212 640740 418116 640782
rect 432332 641018 436332 641060
rect 432332 640782 432374 641018
rect 432610 640782 436054 641018
rect 436290 640782 436332 641018
rect 432332 640740 436332 640782
rect 339964 640060 341204 640380
rect 444660 640380 444980 641420
rect 453492 641698 454180 641740
rect 453492 641462 453902 641698
rect 454138 641462 454180 641698
rect 453492 641420 454180 641462
rect 480724 641698 495764 641740
rect 480724 641462 480766 641698
rect 481002 641462 495764 641698
rect 480724 641420 495764 641462
rect 453492 640380 453812 641420
rect 495444 641060 495764 641420
rect 463428 641018 464116 641060
rect 463428 640782 463470 641018
rect 463706 640782 463838 641018
rect 464074 640782 464116 641018
rect 463428 640740 464116 640782
rect 495444 640740 509380 641060
rect 444660 640060 453812 640380
rect 509060 640338 509380 640740
rect 509060 640102 509102 640338
rect 509338 640102 509380 640338
rect 509060 640060 509380 640102
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect 249436 630138 249940 630180
rect 249436 629902 249478 630138
rect 249714 629902 249940 630138
rect 249436 629860 249940 629902
rect 249620 627460 249940 629860
rect 249252 627418 249940 627460
rect 249252 627182 249294 627418
rect 249530 627182 249940 627418
rect 249252 627140 249940 627182
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect 249252 615858 249940 615900
rect 249252 615622 249294 615858
rect 249530 615622 249940 615858
rect 249252 615580 249940 615622
rect 249620 615220 249940 615580
rect 249436 615178 249940 615220
rect 249436 614942 249478 615178
rect 249714 614942 249940 615178
rect 249436 614900 249940 614942
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect 248700 613138 249572 613180
rect 248700 612902 249294 613138
rect 249530 612902 249572 613138
rect 248700 612860 249572 612902
rect 248700 609100 249020 612860
rect 248700 609058 249388 609100
rect 248700 608822 249110 609058
rect 249346 608822 249388 609058
rect 248700 608780 249388 608822
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect 249252 342498 249756 342540
rect 249252 342262 249478 342498
rect 249714 342262 249756 342498
rect 249252 342220 249756 342262
rect 249252 341860 249572 342220
rect 249068 341818 249572 341860
rect 249068 341582 249110 341818
rect 249346 341582 249572 341818
rect 249068 341540 249572 341582
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1607618424
transform 1 0 230000 0 1 340000
box 0 0 299432 300000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
