magic
tech sky130A
magscale 1 2
timestamp 1608085893
<< locali >>
rect 364533 676243 364567 685797
rect 429577 666587 429611 684437
rect 494069 666587 494103 676141
rect 559297 666587 559331 684437
rect 364533 608651 364567 618205
rect 429393 601715 429427 608549
rect 559113 601715 559147 608549
rect 364625 589339 364659 598893
rect 429577 589339 429611 598893
rect 559297 589339 559331 598893
rect 292129 579071 292163 579309
rect 396733 578595 396767 579309
rect 415685 578527 415719 579309
rect 428381 578459 428415 579309
rect 441077 578391 441111 579309
rect 453589 578323 453623 579309
rect 455797 578255 455831 579309
rect 287069 338011 287103 338113
rect 278789 337807 278823 337977
rect 296637 337875 296671 338113
rect 306389 337875 306423 338113
rect 315957 337875 315991 338113
rect 327215 337909 327273 337943
rect 99389 336855 99423 337093
rect 108957 336855 108991 337229
rect 113189 336787 113223 337229
rect 122757 336787 122791 337229
rect 275293 337195 275327 337773
rect 307033 337467 307067 337773
rect 327089 337467 327123 337841
rect 327181 336855 327215 337501
rect 336749 337467 336783 338793
rect 342821 337535 342855 338113
rect 344661 337875 344695 338113
rect 346409 337739 346443 338657
rect 341717 337127 341751 337501
rect 345581 336991 345615 337569
rect 353953 337263 353987 337501
rect 363981 337263 364015 337637
rect 350549 336855 350583 337229
rect 250177 327131 250211 335529
rect 259837 318835 259871 328389
rect 323317 327131 323351 336685
rect 230857 309179 230891 318733
rect 235089 311831 235123 318733
rect 236285 309179 236319 318733
rect 265265 317475 265299 327029
rect 266645 318835 266679 321589
rect 267749 318835 267783 321589
rect 273545 317543 273579 321725
rect 250177 312579 250211 317373
rect 251557 307819 251591 317373
rect 267749 311151 267783 315945
rect 235089 289867 235123 299421
rect 236285 289867 236319 299421
rect 251373 288439 251407 298061
rect 259653 296735 259687 302277
rect 265265 300135 265299 309077
rect 266645 305031 266679 309213
rect 270785 307819 270819 317373
rect 272257 307819 272291 317373
rect 281733 316047 281767 321589
rect 301053 317475 301087 327029
rect 327273 317475 327307 327029
rect 331413 318903 331447 331857
rect 366925 328491 366959 337841
rect 372261 337807 372295 338045
rect 412557 337671 412591 337977
rect 368213 337195 368247 337569
rect 413477 337059 413511 337637
rect 422309 337603 422343 337977
rect 415501 337195 415535 337569
rect 426081 337127 426115 337501
rect 431601 337195 431635 337365
rect 427829 336855 427863 337093
rect 432613 337059 432647 337501
rect 432705 337127 432739 337501
rect 435189 337127 435223 337569
rect 437121 336651 437155 337501
rect 440157 336855 440191 337977
rect 440249 337739 440283 337909
rect 440341 337399 440375 337909
rect 441905 337467 441939 337909
rect 441997 337671 442031 337909
rect 448529 337501 448713 337535
rect 448529 337467 448563 337501
rect 451105 337467 451139 337977
rect 453221 337467 453255 337773
rect 444423 337161 444573 337195
rect 444515 337093 444665 337127
rect 444515 336957 444573 336991
rect 444297 336651 444331 336889
rect 446965 336855 446999 337365
rect 454693 336855 454727 337977
rect 461501 337977 461719 338011
rect 459017 337331 459051 337773
rect 461501 337671 461535 337977
rect 461685 337943 461719 337977
rect 461593 337671 461627 337909
rect 463433 337875 463467 337909
rect 463433 337841 463617 337875
rect 469137 337807 469171 337977
rect 459109 336923 459143 337297
rect 469229 337263 469263 337977
rect 461593 336855 461627 337229
rect 465031 336889 465215 336923
rect 465181 336719 465215 336889
rect 341349 318835 341383 328389
rect 367017 318835 367051 328321
rect 389465 318835 389499 328389
rect 288725 306391 288759 307717
rect 262597 296735 262631 299625
rect 266737 288439 266771 298061
rect 267841 287079 267875 296565
rect 270785 289867 270819 299421
rect 272257 289323 272291 299421
rect 291577 296531 291611 303569
rect 306849 299523 306883 317373
rect 310897 307887 310931 311933
rect 330217 307819 330251 317373
rect 310713 298163 310747 307717
rect 323225 299523 323259 304249
rect 331413 299591 331447 317373
rect 337117 309111 337151 311933
rect 372721 309179 372755 318733
rect 301053 292519 301087 298061
rect 235089 270555 235123 280109
rect 236285 270555 236319 280109
rect 270693 275315 270727 280109
rect 273545 270555 273579 280109
rect 288909 274703 288943 284257
rect 291393 274703 291427 292485
rect 310897 282795 310931 293029
rect 324697 289867 324731 299421
rect 337117 298163 337151 307717
rect 341165 299523 341199 309077
rect 367017 299523 367051 309077
rect 393605 307819 393639 317373
rect 460213 307819 460247 317373
rect 372721 289867 372755 299421
rect 327181 278783 327215 280177
rect 337117 278783 337151 288337
rect 341165 280211 341199 289765
rect 367017 280211 367051 289765
rect 389373 280211 389407 289765
rect 393605 280211 393639 298061
rect 460029 288439 460063 298061
rect 297005 266407 297039 275961
rect 235089 251243 235123 260797
rect 236285 251243 236319 260797
rect 247233 259607 247267 260865
rect 250177 259471 250211 264265
rect 266737 259471 266771 263585
rect 310897 263483 310931 278681
rect 323317 267767 323351 273309
rect 331413 267767 331447 277321
rect 372721 270555 372755 280109
rect 375849 270555 375883 280109
rect 377137 270555 377171 280109
rect 341165 260899 341199 270453
rect 247233 249747 247267 258009
rect 270693 256003 270727 260797
rect 250177 241519 250211 251141
rect 259653 241587 259687 254609
rect 273545 251243 273579 260797
rect 281825 259471 281859 260865
rect 367017 260899 367051 270453
rect 389373 260899 389407 270453
rect 393605 260899 393639 278681
rect 460121 273139 460155 280109
rect 463801 270555 463835 275281
rect 460029 260967 460063 270453
rect 281825 241519 281859 251141
rect 284677 238799 284711 248353
rect 286057 247095 286091 255901
rect 288817 241519 288851 259097
rect 324605 258111 324639 260865
rect 294245 238799 294279 251821
rect 296821 249475 296855 257941
rect 310897 251311 310931 256037
rect 301053 248455 301087 249849
rect 250177 230503 250211 234617
rect 299489 231863 299523 241417
rect 306757 240091 306791 248353
rect 310713 241519 310747 251141
rect 323409 249815 323443 253929
rect 331413 236691 331447 259369
rect 372721 251243 372755 260797
rect 375849 251243 375883 260797
rect 377137 251243 377171 260797
rect 463709 251243 463743 260797
rect 367017 241519 367051 251073
rect 460029 241519 460063 251141
rect 375849 231863 375883 241417
rect 463801 234651 463835 241417
rect 310805 222207 310839 231761
rect 337301 222207 337335 225301
rect 367017 222207 367051 231761
rect 244381 212483 244415 220745
rect 270693 212551 270727 222105
rect 331413 220847 331447 222173
rect 286057 202895 286091 212449
rect 290197 211123 290231 219385
rect 291669 204323 291703 219385
rect 341165 215271 341199 220745
rect 375849 212551 375883 222105
rect 310805 202895 310839 212449
rect 330125 202827 330159 211089
rect 367017 202895 367051 212449
rect 245853 189091 245887 191845
rect 290013 190519 290047 200073
rect 324605 193171 324639 201433
rect 327181 193171 327215 201433
rect 331413 191811 331447 200073
rect 375849 193239 375883 202793
rect 337117 186303 337151 191777
rect 367017 183583 367051 193137
rect 393513 193103 393547 204901
rect 393513 183515 393547 191777
rect 245761 179435 245795 180897
rect 235089 154615 235123 164169
rect 247141 161483 247175 171037
rect 266645 161483 266679 171037
rect 267841 169779 267875 179333
rect 273545 172567 273579 182121
rect 290013 172567 290047 182121
rect 291669 173723 291703 182121
rect 299857 171139 299891 176749
rect 301053 171139 301087 180761
rect 306849 171139 306883 180761
rect 460121 176511 460155 183481
rect 232329 145027 232363 154513
rect 259745 147611 259779 154513
rect 265357 150467 265391 160021
rect 272349 148291 272383 160021
rect 273545 144891 273579 153153
rect 285965 151827 285999 161381
rect 281733 143599 281767 148325
rect 310805 147611 310839 153153
rect 330217 144959 330251 162741
rect 331597 161483 331631 171037
rect 337117 161483 337151 171037
rect 367017 154683 367051 164169
rect 375849 154615 375883 164169
rect 393605 153255 393639 162809
rect 230857 133943 230891 143497
rect 232329 133943 232363 143497
rect 245853 137955 245887 143497
rect 250177 137955 250211 143497
rect 251373 132515 251407 142069
rect 232329 114563 232363 124117
rect 235089 115991 235123 125545
rect 245945 114563 245979 115957
rect 247325 114563 247359 124117
rect 259653 122859 259687 132413
rect 262597 122859 262631 132413
rect 291393 129659 291427 129897
rect 251373 113203 251407 122757
rect 270785 113203 270819 122757
rect 232329 95251 232363 104805
rect 235089 96679 235123 106233
rect 244381 103547 244415 113101
rect 245945 96679 245979 106233
rect 262505 104907 262539 109701
rect 285965 103547 285999 113101
rect 290013 104227 290047 111741
rect 291485 110483 291519 120037
rect 294429 113203 294463 122757
rect 295717 116603 295751 122757
rect 296913 122723 296947 139349
rect 324789 133943 324823 139893
rect 326077 133943 326111 137717
rect 331413 133943 331447 146013
rect 299765 124219 299799 133841
rect 301053 124219 301087 133841
rect 303905 113203 303939 122757
rect 310805 121499 310839 125749
rect 339785 124287 339819 135201
rect 341349 128299 341383 138669
rect 357633 137955 357667 144857
rect 367017 135371 367051 144857
rect 393605 142171 393639 148461
rect 463709 144959 463743 147713
rect 357541 124219 357575 133841
rect 367017 125647 367051 135201
rect 324605 113203 324639 122757
rect 325893 114427 325927 122757
rect 339785 118031 339819 122757
rect 247141 93891 247175 103445
rect 295717 102187 295751 111741
rect 232329 75939 232363 85493
rect 235089 77299 235123 86921
rect 236285 77299 236319 86921
rect 247141 73219 247175 80053
rect 259745 77299 259779 95149
rect 262597 84303 262631 93789
rect 265265 92531 265299 95285
rect 290013 93823 290047 97937
rect 230765 48331 230799 60605
rect 232329 56627 232363 66045
rect 235089 62747 235123 67541
rect 236285 57987 236319 67541
rect 244381 56627 244415 66181
rect 251373 64923 251407 77197
rect 267841 73219 267875 82773
rect 270693 77299 270727 90389
rect 272165 77299 272199 90389
rect 310805 89675 310839 98685
rect 317705 95251 317739 103377
rect 323409 95251 323443 108001
rect 337025 104907 337059 114461
rect 341165 106335 341199 115889
rect 372813 113203 372847 122757
rect 375757 115991 375791 125545
rect 377045 114563 377079 124117
rect 324605 95251 324639 104805
rect 327181 96611 327215 103445
rect 330125 98719 330159 103377
rect 331413 93891 331447 103445
rect 337209 95251 337243 104737
rect 357633 99331 357667 109701
rect 367017 96747 367051 106233
rect 389373 103547 389407 121397
rect 393605 110483 393639 120037
rect 463893 104907 463927 114461
rect 273545 75939 273579 79985
rect 281825 75939 281859 88961
rect 286057 75939 286091 84949
rect 310805 75939 310839 85493
rect 329941 84235 329975 93789
rect 366925 87091 366959 87193
rect 341073 77299 341107 86921
rect 357633 77299 357667 86921
rect 272165 67643 272199 70533
rect 230765 37315 230799 38709
rect 236285 38675 236319 48229
rect 247233 45611 247267 55165
rect 250177 53839 250211 56593
rect 259929 45679 259963 56525
rect 265265 50915 265299 66181
rect 273545 56627 273579 66181
rect 294245 64923 294279 74477
rect 341073 70295 341107 77129
rect 367017 75939 367051 85493
rect 372721 77299 372755 103377
rect 389281 89675 389315 98685
rect 375849 77299 375883 86921
rect 377137 77299 377171 86921
rect 393605 86887 393639 100657
rect 431325 77299 431359 86921
rect 463709 85595 463743 94129
rect 377137 67643 377171 70465
rect 389373 66283 389407 75837
rect 278881 48331 278915 51153
rect 281733 48331 281767 61421
rect 288725 48331 288759 57001
rect 295533 48331 295567 61421
rect 303905 53839 303939 63461
rect 310805 60707 310839 66181
rect 323409 56627 323443 66181
rect 327181 56627 327215 66181
rect 330125 57851 330159 61421
rect 339785 56627 339819 60809
rect 337117 48331 337151 51085
rect 341349 50643 341383 56525
rect 357633 48331 357667 57885
rect 367017 48399 367051 66181
rect 393697 64923 393731 74477
rect 431325 67643 431359 77129
rect 389189 48331 389223 57545
rect 460029 48331 460063 57885
rect 327365 46971 327399 48297
rect 232237 27659 232271 37145
rect 245761 34527 245795 44081
rect 251373 35955 251407 45509
rect 265173 37315 265207 46869
rect 266737 37315 266771 46869
rect 230765 18003 230799 27557
rect 247233 26367 247267 35853
rect 250085 26299 250119 35785
rect 259561 26367 259595 35853
rect 232145 14127 232179 22729
rect 244197 16643 244231 22117
rect 245853 16643 245887 26197
rect 230673 11203 230707 12461
rect 247141 9163 247175 26197
rect 249993 16643 250027 22117
rect 259561 17935 259595 26197
rect 265265 18071 265299 27557
rect 270785 26299 270819 35853
rect 281733 29019 281767 38573
rect 284769 37315 284803 46869
rect 291485 35955 291519 46869
rect 299765 35955 299799 45509
rect 306941 35955 306975 40749
rect 323317 37315 323351 46869
rect 339785 42075 339819 46869
rect 366833 37315 366867 46869
rect 460029 41395 460063 48161
rect 306665 26367 306699 31093
rect 339693 29019 339727 31773
rect 393605 27659 393639 37213
rect 460121 31739 460155 38573
rect 267749 10659 267783 22593
rect 272073 10863 272107 26197
rect 273453 10931 273487 17901
rect 291577 16643 291611 26197
rect 303997 24871 304031 26265
rect 295533 12223 295567 19261
rect 310897 16643 310931 26197
rect 330217 9707 330251 25857
rect 331413 9707 331447 26197
rect 339693 9707 339727 19193
rect 366833 9707 366867 27557
rect 375849 20859 375883 27557
rect 389373 16643 389407 26197
rect 227545 6987 227579 7633
rect 321569 4947 321603 5049
rect 327181 4947 327215 5049
rect 321569 4913 321753 4947
rect 327031 4913 327215 4947
rect 224233 4811 224267 4913
rect 224141 4267 224175 4777
rect 269129 4063 269163 4233
rect 82829 3043 82863 3213
rect 94973 3009 95249 3043
rect 94973 2975 95007 3009
rect 264621 1139 264655 4029
rect 273453 3859 273487 4097
rect 278697 4063 278731 4233
rect 282929 3723 282963 4029
rect 287621 3995 287655 4165
rect 287713 3723 287747 3961
rect 332333 3927 332367 4097
rect 273269 3043 273303 3213
rect 282837 3043 282871 3349
rect 288633 3315 288667 3825
rect 292497 3315 292531 3689
rect 320649 3451 320683 3621
rect 320833 3587 320867 3893
rect 326353 3723 326387 3893
rect 332241 3791 332275 3893
rect 332149 3587 332183 3757
rect 335369 3587 335403 4097
rect 340797 4097 340889 4131
rect 335921 3723 335955 3893
rect 322765 3111 322799 3553
rect 335737 3043 335771 3553
rect 340647 3145 340739 3179
rect 335829 2975 335863 3145
rect 335645 2839 335679 2941
rect 340705 2907 340739 3145
rect 340797 2839 340831 4097
rect 345489 3315 345523 3349
rect 345489 3281 345707 3315
rect 345673 3247 345707 3281
rect 345581 2839 345615 3213
rect 345949 3179 345983 3349
rect 349169 2975 349203 4097
rect 350181 3247 350215 4437
rect 350549 4403 350583 4505
rect 350583 4029 350675 4063
rect 350641 3655 350675 4029
rect 352389 3995 352423 4097
rect 350549 2907 350583 3621
rect 352481 3247 352515 3961
rect 352941 3383 352975 3961
rect 355057 3961 355425 3995
rect 355057 3655 355091 3961
rect 376769 3927 376803 4913
rect 355425 3451 355459 3621
rect 355517 3383 355551 3621
rect 376861 3519 376895 4981
rect 376803 3485 376895 3519
rect 354873 3349 355551 3383
rect 354873 2975 354907 3349
rect 370329 3315 370363 3417
rect 369903 3281 370363 3315
rect 350549 2873 350825 2907
rect 355517 2771 355551 3077
rect 355609 2907 355643 3077
rect 356069 2975 356103 3213
rect 364993 3111 365027 3281
rect 360301 2975 360335 3009
rect 360301 2941 360485 2975
rect 355735 2805 355977 2839
rect 389465 595 389499 3485
rect 422309 2907 422343 3689
rect 425253 3451 425287 3961
rect 427001 3655 427035 3961
rect 427035 3213 427185 3247
rect 428105 3043 428139 3689
rect 428197 2839 428231 3009
rect 431877 2771 431911 3689
rect 432521 2907 432555 3281
rect 433935 3213 434821 3247
rect 435925 2907 435959 3009
rect 436017 2907 436051 3213
rect 449081 2907 449115 3961
rect 454693 2771 454727 4913
rect 461225 4879 461259 5117
rect 466101 4947 466135 5253
rect 468861 5049 469505 5083
rect 468861 4811 468895 5049
rect 466193 3825 466377 3859
rect 460213 3519 460247 3689
rect 461593 2975 461627 3621
rect 466193 3519 466227 3825
rect 518173 3043 518207 3213
rect 394249 595 394283 1037
<< viali >>
rect 364533 685797 364567 685831
rect 364533 676209 364567 676243
rect 429577 684437 429611 684471
rect 559297 684437 559331 684471
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559297 666553 559331 666587
rect 364533 618205 364567 618239
rect 364533 608617 364567 608651
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 364625 598893 364659 598927
rect 364625 589305 364659 589339
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 292129 579309 292163 579343
rect 292129 579037 292163 579071
rect 396733 579309 396767 579343
rect 396733 578561 396767 578595
rect 415685 579309 415719 579343
rect 415685 578493 415719 578527
rect 428381 579309 428415 579343
rect 428381 578425 428415 578459
rect 441077 579309 441111 579343
rect 441077 578357 441111 578391
rect 453589 579309 453623 579343
rect 453589 578289 453623 578323
rect 455797 579309 455831 579343
rect 455797 578221 455831 578255
rect 336749 338793 336783 338827
rect 287069 338113 287103 338147
rect 278789 337977 278823 338011
rect 287069 337977 287103 338011
rect 296637 338113 296671 338147
rect 296637 337841 296671 337875
rect 306389 338113 306423 338147
rect 306389 337841 306423 337875
rect 315957 338113 315991 338147
rect 327181 337909 327215 337943
rect 327273 337909 327307 337943
rect 315957 337841 315991 337875
rect 327089 337841 327123 337875
rect 275293 337773 275327 337807
rect 278789 337773 278823 337807
rect 307033 337773 307067 337807
rect 108957 337229 108991 337263
rect 99389 337093 99423 337127
rect 99389 336821 99423 336855
rect 108957 336821 108991 336855
rect 113189 337229 113223 337263
rect 113189 336753 113223 336787
rect 122757 337229 122791 337263
rect 307033 337433 307067 337467
rect 327089 337433 327123 337467
rect 327181 337501 327215 337535
rect 275293 337161 275327 337195
rect 346409 338657 346443 338691
rect 342821 338113 342855 338147
rect 344661 338113 344695 338147
rect 344661 337841 344695 337875
rect 372261 338045 372295 338079
rect 346409 337705 346443 337739
rect 366925 337841 366959 337875
rect 363981 337637 364015 337671
rect 336749 337433 336783 337467
rect 341717 337501 341751 337535
rect 342821 337501 342855 337535
rect 345581 337569 345615 337603
rect 341717 337093 341751 337127
rect 353953 337501 353987 337535
rect 345581 336957 345615 336991
rect 350549 337229 350583 337263
rect 353953 337229 353987 337263
rect 363981 337229 364015 337263
rect 327181 336821 327215 336855
rect 350549 336821 350583 336855
rect 122757 336753 122791 336787
rect 323317 336685 323351 336719
rect 250177 335529 250211 335563
rect 250177 327097 250211 327131
rect 259837 328389 259871 328423
rect 323317 327097 323351 327131
rect 331413 331857 331447 331891
rect 259837 318801 259871 318835
rect 265265 327029 265299 327063
rect 230857 318733 230891 318767
rect 235089 318733 235123 318767
rect 235089 311797 235123 311831
rect 236285 318733 236319 318767
rect 230857 309145 230891 309179
rect 301053 327029 301087 327063
rect 273545 321725 273579 321759
rect 266645 321589 266679 321623
rect 266645 318801 266679 318835
rect 267749 321589 267783 321623
rect 267749 318801 267783 318835
rect 273545 317509 273579 317543
rect 281733 321589 281767 321623
rect 265265 317441 265299 317475
rect 250177 317373 250211 317407
rect 250177 312545 250211 312579
rect 251557 317373 251591 317407
rect 236285 309145 236319 309179
rect 270785 317373 270819 317407
rect 267749 315945 267783 315979
rect 267749 311117 267783 311151
rect 266645 309213 266679 309247
rect 251557 307785 251591 307819
rect 265265 309077 265299 309111
rect 259653 302277 259687 302311
rect 235089 299421 235123 299455
rect 235089 289833 235123 289867
rect 236285 299421 236319 299455
rect 236285 289833 236319 289867
rect 251373 298061 251407 298095
rect 270785 307785 270819 307819
rect 272257 317373 272291 317407
rect 301053 317441 301087 317475
rect 327273 327029 327307 327063
rect 372261 337773 372295 337807
rect 412557 337977 412591 338011
rect 422309 337977 422343 338011
rect 412557 337637 412591 337671
rect 413477 337637 413511 337671
rect 368213 337569 368247 337603
rect 368213 337161 368247 337195
rect 440157 337977 440191 338011
rect 415501 337569 415535 337603
rect 422309 337569 422343 337603
rect 435189 337569 435223 337603
rect 415501 337161 415535 337195
rect 426081 337501 426115 337535
rect 432613 337501 432647 337535
rect 431601 337365 431635 337399
rect 431601 337161 431635 337195
rect 426081 337093 426115 337127
rect 427829 337093 427863 337127
rect 413477 337025 413511 337059
rect 432705 337501 432739 337535
rect 432705 337093 432739 337127
rect 435189 337093 435223 337127
rect 437121 337501 437155 337535
rect 432613 337025 432647 337059
rect 427829 336821 427863 336855
rect 451105 337977 451139 338011
rect 440249 337909 440283 337943
rect 440249 337705 440283 337739
rect 440341 337909 440375 337943
rect 441905 337909 441939 337943
rect 441997 337909 442031 337943
rect 441997 337637 442031 337671
rect 441905 337433 441939 337467
rect 448713 337501 448747 337535
rect 448529 337433 448563 337467
rect 454693 337977 454727 338011
rect 451105 337433 451139 337467
rect 453221 337773 453255 337807
rect 453221 337433 453255 337467
rect 440341 337365 440375 337399
rect 446965 337365 446999 337399
rect 444389 337161 444423 337195
rect 444573 337161 444607 337195
rect 444481 337093 444515 337127
rect 444665 337093 444699 337127
rect 444481 336957 444515 336991
rect 444573 336957 444607 336991
rect 440157 336821 440191 336855
rect 444297 336889 444331 336923
rect 437121 336617 437155 336651
rect 446965 336821 446999 336855
rect 459017 337773 459051 337807
rect 469137 337977 469171 338011
rect 461501 337637 461535 337671
rect 461593 337909 461627 337943
rect 461685 337909 461719 337943
rect 463433 337909 463467 337943
rect 463617 337841 463651 337875
rect 469137 337773 469171 337807
rect 469229 337977 469263 338011
rect 461593 337637 461627 337671
rect 459017 337297 459051 337331
rect 459109 337297 459143 337331
rect 459109 336889 459143 336923
rect 461593 337229 461627 337263
rect 469229 337229 469263 337263
rect 454693 336821 454727 336855
rect 464997 336889 465031 336923
rect 461593 336821 461627 336855
rect 465181 336685 465215 336719
rect 444297 336617 444331 336651
rect 366925 328457 366959 328491
rect 331413 318869 331447 318903
rect 341349 328389 341383 328423
rect 389465 328389 389499 328423
rect 341349 318801 341383 318835
rect 367017 328321 367051 328355
rect 367017 318801 367051 318835
rect 389465 318801 389499 318835
rect 327273 317441 327307 317475
rect 372721 318733 372755 318767
rect 281733 316013 281767 316047
rect 306849 317373 306883 317407
rect 272257 307785 272291 307819
rect 288725 307717 288759 307751
rect 288725 306357 288759 306391
rect 266645 304997 266679 305031
rect 265265 300101 265299 300135
rect 291577 303569 291611 303603
rect 259653 296701 259687 296735
rect 262597 299625 262631 299659
rect 270785 299421 270819 299455
rect 262597 296701 262631 296735
rect 266737 298061 266771 298095
rect 251373 288405 251407 288439
rect 266737 288405 266771 288439
rect 267841 296565 267875 296599
rect 270785 289833 270819 289867
rect 272257 299421 272291 299455
rect 330217 317373 330251 317407
rect 310897 311933 310931 311967
rect 310897 307853 310931 307887
rect 330217 307785 330251 307819
rect 331413 317373 331447 317407
rect 306849 299489 306883 299523
rect 310713 307717 310747 307751
rect 323225 304249 323259 304283
rect 337117 311933 337151 311967
rect 372721 309145 372755 309179
rect 393605 317373 393639 317407
rect 337117 309077 337151 309111
rect 341165 309077 341199 309111
rect 331413 299557 331447 299591
rect 337117 307717 337151 307751
rect 323225 299489 323259 299523
rect 310713 298129 310747 298163
rect 324697 299421 324731 299455
rect 291577 296497 291611 296531
rect 301053 298061 301087 298095
rect 272257 289289 272291 289323
rect 291393 292485 291427 292519
rect 301053 292485 301087 292519
rect 310897 293029 310931 293063
rect 267841 287045 267875 287079
rect 288909 284257 288943 284291
rect 235089 280109 235123 280143
rect 235089 270521 235123 270555
rect 236285 280109 236319 280143
rect 270693 280109 270727 280143
rect 270693 275281 270727 275315
rect 273545 280109 273579 280143
rect 236285 270521 236319 270555
rect 288909 274669 288943 274703
rect 341165 299489 341199 299523
rect 367017 309077 367051 309111
rect 393605 307785 393639 307819
rect 460213 317373 460247 317407
rect 460213 307785 460247 307819
rect 367017 299489 367051 299523
rect 337117 298129 337151 298163
rect 372721 299421 372755 299455
rect 324697 289833 324731 289867
rect 372721 289833 372755 289867
rect 393605 298061 393639 298095
rect 341165 289765 341199 289799
rect 310897 282761 310931 282795
rect 337117 288337 337151 288371
rect 327181 280177 327215 280211
rect 327181 278749 327215 278783
rect 341165 280177 341199 280211
rect 367017 289765 367051 289799
rect 367017 280177 367051 280211
rect 389373 289765 389407 289799
rect 389373 280177 389407 280211
rect 460029 298061 460063 298095
rect 460029 288405 460063 288439
rect 393605 280177 393639 280211
rect 337117 278749 337151 278783
rect 372721 280109 372755 280143
rect 310897 278681 310931 278715
rect 291393 274669 291427 274703
rect 297005 275961 297039 275995
rect 273545 270521 273579 270555
rect 297005 266373 297039 266407
rect 250177 264265 250211 264299
rect 247233 260865 247267 260899
rect 235089 260797 235123 260831
rect 235089 251209 235123 251243
rect 236285 260797 236319 260831
rect 247233 259573 247267 259607
rect 250177 259437 250211 259471
rect 266737 263585 266771 263619
rect 331413 277321 331447 277355
rect 323317 273309 323351 273343
rect 323317 267733 323351 267767
rect 372721 270521 372755 270555
rect 375849 280109 375883 280143
rect 375849 270521 375883 270555
rect 377137 280109 377171 280143
rect 460121 280109 460155 280143
rect 377137 270521 377171 270555
rect 393605 278681 393639 278715
rect 331413 267733 331447 267767
rect 341165 270453 341199 270487
rect 310897 263449 310931 263483
rect 281825 260865 281859 260899
rect 266737 259437 266771 259471
rect 270693 260797 270727 260831
rect 236285 251209 236319 251243
rect 247233 258009 247267 258043
rect 270693 255969 270727 256003
rect 273545 260797 273579 260831
rect 259653 254609 259687 254643
rect 247233 249713 247267 249747
rect 250177 251141 250211 251175
rect 281825 259437 281859 259471
rect 324605 260865 324639 260899
rect 341165 260865 341199 260899
rect 367017 270453 367051 270487
rect 367017 260865 367051 260899
rect 389373 270453 389407 270487
rect 389373 260865 389407 260899
rect 460121 273105 460155 273139
rect 463801 275281 463835 275315
rect 463801 270521 463835 270555
rect 460029 270453 460063 270487
rect 460029 260933 460063 260967
rect 393605 260865 393639 260899
rect 288817 259097 288851 259131
rect 273545 251209 273579 251243
rect 286057 255901 286091 255935
rect 259653 241553 259687 241587
rect 281825 251141 281859 251175
rect 250177 241485 250211 241519
rect 281825 241485 281859 241519
rect 284677 248353 284711 248387
rect 286057 247061 286091 247095
rect 372721 260797 372755 260831
rect 324605 258077 324639 258111
rect 331413 259369 331447 259403
rect 296821 257941 296855 257975
rect 288817 241485 288851 241519
rect 294245 251821 294279 251855
rect 284677 238765 284711 238799
rect 310897 256037 310931 256071
rect 310897 251277 310931 251311
rect 323409 253929 323443 253963
rect 310713 251141 310747 251175
rect 296821 249441 296855 249475
rect 301053 249849 301087 249883
rect 301053 248421 301087 248455
rect 306757 248353 306791 248387
rect 294245 238765 294279 238799
rect 299489 241417 299523 241451
rect 250177 234617 250211 234651
rect 323409 249781 323443 249815
rect 310713 241485 310747 241519
rect 306757 240057 306791 240091
rect 372721 251209 372755 251243
rect 375849 260797 375883 260831
rect 375849 251209 375883 251243
rect 377137 260797 377171 260831
rect 377137 251209 377171 251243
rect 463709 260797 463743 260831
rect 463709 251209 463743 251243
rect 460029 251141 460063 251175
rect 367017 251073 367051 251107
rect 367017 241485 367051 241519
rect 460029 241485 460063 241519
rect 331413 236657 331447 236691
rect 375849 241417 375883 241451
rect 299489 231829 299523 231863
rect 463801 241417 463835 241451
rect 463801 234617 463835 234651
rect 375849 231829 375883 231863
rect 250177 230469 250211 230503
rect 310805 231761 310839 231795
rect 367017 231761 367051 231795
rect 337301 225301 337335 225335
rect 310805 222173 310839 222207
rect 331413 222173 331447 222207
rect 337301 222173 337335 222207
rect 367017 222173 367051 222207
rect 270693 222105 270727 222139
rect 244381 220745 244415 220779
rect 331413 220813 331447 220847
rect 375849 222105 375883 222139
rect 341165 220745 341199 220779
rect 270693 212517 270727 212551
rect 290197 219385 290231 219419
rect 244381 212449 244415 212483
rect 286057 212449 286091 212483
rect 290197 211089 290231 211123
rect 291669 219385 291703 219419
rect 341165 215237 341199 215271
rect 375849 212517 375883 212551
rect 291669 204289 291703 204323
rect 310805 212449 310839 212483
rect 286057 202861 286091 202895
rect 367017 212449 367051 212483
rect 310805 202861 310839 202895
rect 330125 211089 330159 211123
rect 367017 202861 367051 202895
rect 393513 204901 393547 204935
rect 330125 202793 330159 202827
rect 375849 202793 375883 202827
rect 324605 201433 324639 201467
rect 290013 200073 290047 200107
rect 245853 191845 245887 191879
rect 324605 193137 324639 193171
rect 327181 201433 327215 201467
rect 327181 193137 327215 193171
rect 331413 200073 331447 200107
rect 375849 193205 375883 193239
rect 367017 193137 367051 193171
rect 331413 191777 331447 191811
rect 337117 191777 337151 191811
rect 290013 190485 290047 190519
rect 245853 189057 245887 189091
rect 337117 186269 337151 186303
rect 393513 193069 393547 193103
rect 367017 183549 367051 183583
rect 393513 191777 393547 191811
rect 393513 183481 393547 183515
rect 460121 183481 460155 183515
rect 273545 182121 273579 182155
rect 245761 180897 245795 180931
rect 245761 179401 245795 179435
rect 267841 179333 267875 179367
rect 247141 171037 247175 171071
rect 235089 164169 235123 164203
rect 247141 161449 247175 161483
rect 266645 171037 266679 171071
rect 273545 172533 273579 172567
rect 290013 182121 290047 182155
rect 291669 182121 291703 182155
rect 301053 180761 301087 180795
rect 291669 173689 291703 173723
rect 299857 176749 299891 176783
rect 290013 172533 290047 172567
rect 299857 171105 299891 171139
rect 301053 171105 301087 171139
rect 306849 180761 306883 180795
rect 460121 176477 460155 176511
rect 306849 171105 306883 171139
rect 267841 169745 267875 169779
rect 331597 171037 331631 171071
rect 266645 161449 266679 161483
rect 330217 162741 330251 162775
rect 285965 161381 285999 161415
rect 235089 154581 235123 154615
rect 265357 160021 265391 160055
rect 232329 154513 232363 154547
rect 259745 154513 259779 154547
rect 265357 150433 265391 150467
rect 272349 160021 272383 160055
rect 272349 148257 272383 148291
rect 273545 153153 273579 153187
rect 259745 147577 259779 147611
rect 232329 144993 232363 145027
rect 285965 151793 285999 151827
rect 310805 153153 310839 153187
rect 273545 144857 273579 144891
rect 281733 148325 281767 148359
rect 310805 147577 310839 147611
rect 331597 161449 331631 161483
rect 337117 171037 337151 171071
rect 337117 161449 337151 161483
rect 367017 164169 367051 164203
rect 367017 154649 367051 154683
rect 375849 164169 375883 164203
rect 375849 154581 375883 154615
rect 393605 162809 393639 162843
rect 393605 153221 393639 153255
rect 393605 148461 393639 148495
rect 330217 144925 330251 144959
rect 331413 146013 331447 146047
rect 281733 143565 281767 143599
rect 230857 143497 230891 143531
rect 230857 133909 230891 133943
rect 232329 143497 232363 143531
rect 245853 143497 245887 143531
rect 245853 137921 245887 137955
rect 250177 143497 250211 143531
rect 250177 137921 250211 137955
rect 251373 142069 251407 142103
rect 232329 133909 232363 133943
rect 324789 139893 324823 139927
rect 251373 132481 251407 132515
rect 296913 139349 296947 139383
rect 259653 132413 259687 132447
rect 235089 125545 235123 125579
rect 232329 124117 232363 124151
rect 247325 124117 247359 124151
rect 235089 115957 235123 115991
rect 245945 115957 245979 115991
rect 232329 114529 232363 114563
rect 245945 114529 245979 114563
rect 259653 122825 259687 122859
rect 262597 132413 262631 132447
rect 291393 129897 291427 129931
rect 291393 129625 291427 129659
rect 262597 122825 262631 122859
rect 247325 114529 247359 114563
rect 251373 122757 251407 122791
rect 251373 113169 251407 113203
rect 270785 122757 270819 122791
rect 294429 122757 294463 122791
rect 270785 113169 270819 113203
rect 291485 120037 291519 120071
rect 244381 113101 244415 113135
rect 235089 106233 235123 106267
rect 232329 104805 232363 104839
rect 285965 113101 285999 113135
rect 262505 109701 262539 109735
rect 244381 103513 244415 103547
rect 245945 106233 245979 106267
rect 235089 96645 235123 96679
rect 262505 104873 262539 104907
rect 290013 111741 290047 111775
rect 295717 122757 295751 122791
rect 324789 133909 324823 133943
rect 326077 137717 326111 137751
rect 326077 133909 326111 133943
rect 357633 144857 357667 144891
rect 341349 138669 341383 138703
rect 331413 133909 331447 133943
rect 339785 135201 339819 135235
rect 299765 133841 299799 133875
rect 299765 124185 299799 124219
rect 301053 133841 301087 133875
rect 301053 124185 301087 124219
rect 310805 125749 310839 125783
rect 296913 122689 296947 122723
rect 303905 122757 303939 122791
rect 295717 116569 295751 116603
rect 294429 113169 294463 113203
rect 357633 137921 357667 137955
rect 367017 144857 367051 144891
rect 463709 147713 463743 147747
rect 463709 144925 463743 144959
rect 393605 142137 393639 142171
rect 367017 135337 367051 135371
rect 367017 135201 367051 135235
rect 341349 128265 341383 128299
rect 357541 133841 357575 133875
rect 339785 124253 339819 124287
rect 367017 125613 367051 125647
rect 357541 124185 357575 124219
rect 375757 125545 375791 125579
rect 310805 121465 310839 121499
rect 324605 122757 324639 122791
rect 303905 113169 303939 113203
rect 325893 122757 325927 122791
rect 339785 122757 339819 122791
rect 339785 117997 339819 118031
rect 372813 122757 372847 122791
rect 341165 115889 341199 115923
rect 325893 114393 325927 114427
rect 337025 114461 337059 114495
rect 324605 113169 324639 113203
rect 291485 110449 291519 110483
rect 295717 111741 295751 111775
rect 290013 104193 290047 104227
rect 285965 103513 285999 103547
rect 245945 96645 245979 96679
rect 247141 103445 247175 103479
rect 232329 95217 232363 95251
rect 323409 108001 323443 108035
rect 295717 102153 295751 102187
rect 317705 103377 317739 103411
rect 310805 98685 310839 98719
rect 290013 97937 290047 97971
rect 265265 95285 265299 95319
rect 247141 93857 247175 93891
rect 259745 95149 259779 95183
rect 235089 86921 235123 86955
rect 232329 85493 232363 85527
rect 235089 77265 235123 77299
rect 236285 86921 236319 86955
rect 236285 77265 236319 77299
rect 247141 80053 247175 80087
rect 232329 75905 232363 75939
rect 262597 93789 262631 93823
rect 290013 93789 290047 93823
rect 265265 92497 265299 92531
rect 262597 84269 262631 84303
rect 270693 90389 270727 90423
rect 259745 77265 259779 77299
rect 267841 82773 267875 82807
rect 247141 73185 247175 73219
rect 251373 77197 251407 77231
rect 235089 67541 235123 67575
rect 232329 66045 232363 66079
rect 230765 60605 230799 60639
rect 235089 62713 235123 62747
rect 236285 67541 236319 67575
rect 236285 57953 236319 57987
rect 244381 66181 244415 66215
rect 232329 56593 232363 56627
rect 270693 77265 270727 77299
rect 272165 90389 272199 90423
rect 317705 95217 317739 95251
rect 375757 115957 375791 115991
rect 377045 124117 377079 124151
rect 377045 114529 377079 114563
rect 389373 121397 389407 121431
rect 372813 113169 372847 113203
rect 341165 106301 341199 106335
rect 357633 109701 357667 109735
rect 337025 104873 337059 104907
rect 323409 95217 323443 95251
rect 324605 104805 324639 104839
rect 337209 104737 337243 104771
rect 327181 103445 327215 103479
rect 331413 103445 331447 103479
rect 330125 103377 330159 103411
rect 330125 98685 330159 98719
rect 327181 96577 327215 96611
rect 324605 95217 324639 95251
rect 357633 99297 357667 99331
rect 367017 106233 367051 106267
rect 393605 120037 393639 120071
rect 393605 110449 393639 110483
rect 463893 114461 463927 114495
rect 463893 104873 463927 104907
rect 389373 103513 389407 103547
rect 367017 96713 367051 96747
rect 372721 103377 372755 103411
rect 337209 95217 337243 95251
rect 331413 93857 331447 93891
rect 310805 89641 310839 89675
rect 329941 93789 329975 93823
rect 281825 88961 281859 88995
rect 272165 77265 272199 77299
rect 273545 79985 273579 80019
rect 273545 75905 273579 75939
rect 310805 85493 310839 85527
rect 281825 75905 281859 75939
rect 286057 84949 286091 84983
rect 286057 75905 286091 75939
rect 366925 87193 366959 87227
rect 366925 87057 366959 87091
rect 329941 84201 329975 84235
rect 341073 86921 341107 86955
rect 341073 77265 341107 77299
rect 357633 86921 357667 86955
rect 357633 77265 357667 77299
rect 367017 85493 367051 85527
rect 310805 75905 310839 75939
rect 341073 77129 341107 77163
rect 267841 73185 267875 73219
rect 294245 74477 294279 74511
rect 272165 70533 272199 70567
rect 272165 67609 272199 67643
rect 251373 64889 251407 64923
rect 265265 66181 265299 66215
rect 244381 56593 244415 56627
rect 250177 56593 250211 56627
rect 230765 48297 230799 48331
rect 247233 55165 247267 55199
rect 236285 48229 236319 48263
rect 230765 38709 230799 38743
rect 250177 53805 250211 53839
rect 259929 56525 259963 56559
rect 273545 66181 273579 66215
rect 393605 100657 393639 100691
rect 389281 98685 389315 98719
rect 389281 89641 389315 89675
rect 372721 77265 372755 77299
rect 375849 86921 375883 86955
rect 375849 77265 375883 77299
rect 377137 86921 377171 86955
rect 463709 94129 463743 94163
rect 393605 86853 393639 86887
rect 431325 86921 431359 86955
rect 377137 77265 377171 77299
rect 463709 85561 463743 85595
rect 431325 77265 431359 77299
rect 367017 75905 367051 75939
rect 431325 77129 431359 77163
rect 389373 75837 389407 75871
rect 341073 70261 341107 70295
rect 377137 70465 377171 70499
rect 377137 67609 377171 67643
rect 389373 66249 389407 66283
rect 393697 74477 393731 74511
rect 294245 64889 294279 64923
rect 310805 66181 310839 66215
rect 303905 63461 303939 63495
rect 273545 56593 273579 56627
rect 281733 61421 281767 61455
rect 265265 50881 265299 50915
rect 278881 51153 278915 51187
rect 278881 48297 278915 48331
rect 295533 61421 295567 61455
rect 281733 48297 281767 48331
rect 288725 57001 288759 57035
rect 288725 48297 288759 48331
rect 310805 60673 310839 60707
rect 323409 66181 323443 66215
rect 323409 56593 323443 56627
rect 327181 66181 327215 66215
rect 367017 66181 367051 66215
rect 330125 61421 330159 61455
rect 330125 57817 330159 57851
rect 339785 60809 339819 60843
rect 327181 56593 327215 56627
rect 339785 56593 339819 56627
rect 357633 57885 357667 57919
rect 303905 53805 303939 53839
rect 341349 56525 341383 56559
rect 337117 51085 337151 51119
rect 341349 50609 341383 50643
rect 295533 48297 295567 48331
rect 327365 48297 327399 48331
rect 337117 48297 337151 48331
rect 431325 67609 431359 67643
rect 393697 64889 393731 64923
rect 460029 57885 460063 57919
rect 367017 48365 367051 48399
rect 389189 57545 389223 57579
rect 357633 48297 357667 48331
rect 389189 48297 389223 48331
rect 460029 48297 460063 48331
rect 327365 46937 327399 46971
rect 460029 48161 460063 48195
rect 259929 45645 259963 45679
rect 265173 46869 265207 46903
rect 247233 45577 247267 45611
rect 251373 45509 251407 45543
rect 236285 38641 236319 38675
rect 245761 44081 245795 44115
rect 230765 37281 230799 37315
rect 232237 37145 232271 37179
rect 265173 37281 265207 37315
rect 266737 46869 266771 46903
rect 284769 46869 284803 46903
rect 266737 37281 266771 37315
rect 281733 38573 281767 38607
rect 251373 35921 251407 35955
rect 245761 34493 245795 34527
rect 247233 35853 247267 35887
rect 232237 27625 232271 27659
rect 230765 27557 230799 27591
rect 259561 35853 259595 35887
rect 247233 26333 247267 26367
rect 250085 35785 250119 35819
rect 270785 35853 270819 35887
rect 259561 26333 259595 26367
rect 265265 27557 265299 27591
rect 250085 26265 250119 26299
rect 245853 26197 245887 26231
rect 230765 17969 230799 18003
rect 232145 22729 232179 22763
rect 244197 22117 244231 22151
rect 244197 16609 244231 16643
rect 245853 16609 245887 16643
rect 247141 26197 247175 26231
rect 232145 14093 232179 14127
rect 230673 12461 230707 12495
rect 230673 11169 230707 11203
rect 259561 26197 259595 26231
rect 249993 22117 250027 22151
rect 284769 37281 284803 37315
rect 291485 46869 291519 46903
rect 323317 46869 323351 46903
rect 291485 35921 291519 35955
rect 299765 45509 299799 45543
rect 299765 35921 299799 35955
rect 306941 40749 306975 40783
rect 339785 46869 339819 46903
rect 339785 42041 339819 42075
rect 366833 46869 366867 46903
rect 323317 37281 323351 37315
rect 460029 41361 460063 41395
rect 366833 37281 366867 37315
rect 460121 38573 460155 38607
rect 306941 35921 306975 35955
rect 393605 37213 393639 37247
rect 339693 31773 339727 31807
rect 281733 28985 281767 29019
rect 306665 31093 306699 31127
rect 339693 28985 339727 29019
rect 460121 31705 460155 31739
rect 393605 27625 393639 27659
rect 306665 26333 306699 26367
rect 366833 27557 366867 27591
rect 270785 26265 270819 26299
rect 303997 26265 304031 26299
rect 272073 26197 272107 26231
rect 265265 18037 265299 18071
rect 267749 22593 267783 22627
rect 259561 17901 259595 17935
rect 249993 16609 250027 16643
rect 291577 26197 291611 26231
rect 273453 17901 273487 17935
rect 303997 24837 304031 24871
rect 310897 26197 310931 26231
rect 291577 16609 291611 16643
rect 295533 19261 295567 19295
rect 331413 26197 331447 26231
rect 310897 16609 310931 16643
rect 330217 25857 330251 25891
rect 295533 12189 295567 12223
rect 273453 10897 273487 10931
rect 272073 10829 272107 10863
rect 267749 10625 267783 10659
rect 330217 9673 330251 9707
rect 331413 9673 331447 9707
rect 339693 19193 339727 19227
rect 339693 9673 339727 9707
rect 375849 27557 375883 27591
rect 375849 20825 375883 20859
rect 389373 26197 389407 26231
rect 389373 16609 389407 16643
rect 366833 9673 366867 9707
rect 247141 9129 247175 9163
rect 227545 7633 227579 7667
rect 227545 6953 227579 6987
rect 466101 5253 466135 5287
rect 461225 5117 461259 5151
rect 321569 5049 321603 5083
rect 327181 5049 327215 5083
rect 376861 4981 376895 5015
rect 224233 4913 224267 4947
rect 321753 4913 321787 4947
rect 326997 4913 327031 4947
rect 376769 4913 376803 4947
rect 224141 4777 224175 4811
rect 224233 4777 224267 4811
rect 350549 4505 350583 4539
rect 350181 4437 350215 4471
rect 224141 4233 224175 4267
rect 269129 4233 269163 4267
rect 278697 4233 278731 4267
rect 264621 4029 264655 4063
rect 269129 4029 269163 4063
rect 273453 4097 273487 4131
rect 82829 3213 82863 3247
rect 82829 3009 82863 3043
rect 95249 3009 95283 3043
rect 94973 2941 95007 2975
rect 287621 4165 287655 4199
rect 278697 4029 278731 4063
rect 282929 4029 282963 4063
rect 273453 3825 273487 3859
rect 332333 4097 332367 4131
rect 287621 3961 287655 3995
rect 287713 3961 287747 3995
rect 282929 3689 282963 3723
rect 320833 3893 320867 3927
rect 287713 3689 287747 3723
rect 288633 3825 288667 3859
rect 282837 3349 282871 3383
rect 273269 3213 273303 3247
rect 273269 3009 273303 3043
rect 288633 3281 288667 3315
rect 292497 3689 292531 3723
rect 320649 3621 320683 3655
rect 326353 3893 326387 3927
rect 332241 3893 332275 3927
rect 332333 3893 332367 3927
rect 335369 4097 335403 4131
rect 326353 3689 326387 3723
rect 332149 3757 332183 3791
rect 332241 3757 332275 3791
rect 320833 3553 320867 3587
rect 322765 3553 322799 3587
rect 332149 3553 332183 3587
rect 340889 4097 340923 4131
rect 349169 4097 349203 4131
rect 335921 3893 335955 3927
rect 335921 3689 335955 3723
rect 335369 3553 335403 3587
rect 335737 3553 335771 3587
rect 320649 3417 320683 3451
rect 292497 3281 292531 3315
rect 322765 3077 322799 3111
rect 282837 3009 282871 3043
rect 335737 3009 335771 3043
rect 335829 3145 335863 3179
rect 340613 3145 340647 3179
rect 335645 2941 335679 2975
rect 335829 2941 335863 2975
rect 340705 2873 340739 2907
rect 335645 2805 335679 2839
rect 345489 3349 345523 3383
rect 345949 3349 345983 3383
rect 340797 2805 340831 2839
rect 345581 3213 345615 3247
rect 345673 3213 345707 3247
rect 345949 3145 345983 3179
rect 350549 4369 350583 4403
rect 352389 4097 352423 4131
rect 350549 4029 350583 4063
rect 352389 3961 352423 3995
rect 352481 3961 352515 3995
rect 350181 3213 350215 3247
rect 350549 3621 350583 3655
rect 350641 3621 350675 3655
rect 349169 2941 349203 2975
rect 352941 3961 352975 3995
rect 355425 3961 355459 3995
rect 376769 3893 376803 3927
rect 355057 3621 355091 3655
rect 355425 3621 355459 3655
rect 355425 3417 355459 3451
rect 355517 3621 355551 3655
rect 454693 4913 454727 4947
rect 425253 3961 425287 3995
rect 422309 3689 422343 3723
rect 376769 3485 376803 3519
rect 389465 3485 389499 3519
rect 352941 3349 352975 3383
rect 370329 3417 370363 3451
rect 352481 3213 352515 3247
rect 364993 3281 365027 3315
rect 369869 3281 369903 3315
rect 356069 3213 356103 3247
rect 354873 2941 354907 2975
rect 355517 3077 355551 3111
rect 350825 2873 350859 2907
rect 345581 2805 345615 2839
rect 355609 3077 355643 3111
rect 364993 3077 365027 3111
rect 356069 2941 356103 2975
rect 360301 3009 360335 3043
rect 360485 2941 360519 2975
rect 355609 2873 355643 2907
rect 355701 2805 355735 2839
rect 355977 2805 356011 2839
rect 355517 2737 355551 2771
rect 264621 1105 264655 1139
rect 427001 3961 427035 3995
rect 449081 3961 449115 3995
rect 427001 3621 427035 3655
rect 428105 3689 428139 3723
rect 425253 3417 425287 3451
rect 427001 3213 427035 3247
rect 427185 3213 427219 3247
rect 431877 3689 431911 3723
rect 428105 3009 428139 3043
rect 428197 3009 428231 3043
rect 422309 2873 422343 2907
rect 428197 2805 428231 2839
rect 432521 3281 432555 3315
rect 433901 3213 433935 3247
rect 434821 3213 434855 3247
rect 436017 3213 436051 3247
rect 432521 2873 432555 2907
rect 435925 3009 435959 3043
rect 435925 2873 435959 2907
rect 436017 2873 436051 2907
rect 449081 2873 449115 2907
rect 431877 2737 431911 2771
rect 466101 4913 466135 4947
rect 469505 5049 469539 5083
rect 461225 4845 461259 4879
rect 468861 4777 468895 4811
rect 466377 3825 466411 3859
rect 460213 3689 460247 3723
rect 460213 3485 460247 3519
rect 461593 3621 461627 3655
rect 466193 3485 466227 3519
rect 518173 3213 518207 3247
rect 518173 3009 518207 3043
rect 461593 2941 461627 2975
rect 454693 2737 454727 2771
rect 389465 561 389499 595
rect 394249 1037 394283 1071
rect 394249 561 394283 595
<< metal1 >>
rect 202782 700952 202788 701004
rect 202840 700992 202846 701004
rect 358814 700992 358820 701004
rect 202840 700964 358820 700992
rect 202840 700952 202846 700964
rect 358814 700952 358820 700964
rect 358872 700952 358878 701004
rect 170306 700884 170312 700936
rect 170364 700924 170370 700936
rect 362954 700924 362960 700936
rect 170364 700896 362960 700924
rect 170364 700884 170370 700896
rect 362954 700884 362960 700896
rect 363012 700884 363018 700936
rect 328362 700816 328368 700868
rect 328420 700856 328426 700868
rect 527174 700856 527180 700868
rect 328420 700828 527180 700856
rect 328420 700816 328426 700828
rect 527174 700816 527180 700828
rect 527232 700816 527238 700868
rect 329742 700748 329748 700800
rect 329800 700788 329806 700800
rect 543458 700788 543464 700800
rect 329800 700760 543464 700788
rect 329800 700748 329806 700760
rect 543458 700748 543464 700760
rect 543516 700748 543522 700800
rect 154114 700680 154120 700732
rect 154172 700720 154178 700732
rect 367094 700720 367100 700732
rect 154172 700692 367100 700720
rect 154172 700680 154178 700692
rect 367094 700680 367100 700692
rect 367152 700680 367158 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 364334 700652 364340 700664
rect 137888 700624 364340 700652
rect 137888 700612 137894 700624
rect 364334 700612 364340 700624
rect 364392 700612 364398 700664
rect 105446 700544 105452 700596
rect 105504 700584 105510 700596
rect 368474 700584 368480 700596
rect 105504 700556 368480 700584
rect 105504 700544 105510 700556
rect 368474 700544 368480 700556
rect 368532 700544 368538 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 373994 700516 374000 700528
rect 89220 700488 374000 700516
rect 89220 700476 89226 700488
rect 373994 700476 374000 700488
rect 374052 700476 374058 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 371234 700448 371240 700460
rect 73028 700420 371240 700448
rect 73028 700408 73034 700420
rect 371234 700408 371240 700420
rect 371292 700408 371298 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 375374 700380 375380 700392
rect 40552 700352 375380 700380
rect 40552 700340 40558 700352
rect 375374 700340 375380 700352
rect 375432 700340 375438 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 379514 700312 379520 700324
rect 24360 700284 379520 700312
rect 24360 700272 24366 700284
rect 379514 700272 379520 700284
rect 379572 700272 379578 700324
rect 218974 700204 218980 700256
rect 219032 700244 219038 700256
rect 360194 700244 360200 700256
rect 219032 700216 360200 700244
rect 219032 700204 219038 700216
rect 360194 700204 360200 700216
rect 360252 700204 360258 700256
rect 336642 700136 336648 700188
rect 336700 700176 336706 700188
rect 478506 700176 478512 700188
rect 336700 700148 478512 700176
rect 336700 700136 336706 700148
rect 478506 700136 478512 700148
rect 478564 700136 478570 700188
rect 335262 700068 335268 700120
rect 335320 700108 335326 700120
rect 462314 700108 462320 700120
rect 335320 700080 462320 700108
rect 335320 700068 335326 700080
rect 462314 700068 462320 700080
rect 462372 700068 462378 700120
rect 235166 700000 235172 700052
rect 235224 700040 235230 700052
rect 356054 700040 356060 700052
rect 235224 700012 356060 700040
rect 235224 700000 235230 700012
rect 356054 700000 356060 700012
rect 356112 700000 356118 700052
rect 267642 699932 267648 699984
rect 267700 699972 267706 699984
rect 351914 699972 351920 699984
rect 267700 699944 351920 699972
rect 267700 699932 267706 699944
rect 351914 699932 351920 699944
rect 351972 699932 351978 699984
rect 283834 699864 283840 699916
rect 283892 699904 283898 699916
rect 354674 699904 354680 699916
rect 283892 699876 354680 699904
rect 283892 699864 283898 699876
rect 354674 699864 354680 699876
rect 354732 699864 354738 699916
rect 343542 699796 343548 699848
rect 343600 699836 343606 699848
rect 413646 699836 413652 699848
rect 343600 699808 413652 699836
rect 343600 699796 343606 699808
rect 413646 699796 413652 699808
rect 413704 699796 413710 699848
rect 340782 699728 340788 699780
rect 340840 699768 340846 699780
rect 397454 699768 397460 699780
rect 340840 699740 397460 699768
rect 340840 699728 340846 699740
rect 397454 699728 397460 699740
rect 397512 699728 397518 699780
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 332502 699660 332508 699712
rect 332560 699700 332566 699712
rect 346394 699700 346400 699712
rect 332560 699672 346400 699700
rect 332560 699660 332566 699672
rect 346394 699660 346400 699672
rect 346452 699660 346458 699712
rect 347774 699660 347780 699712
rect 347832 699700 347838 699712
rect 348786 699700 348792 699712
rect 347832 699672 348792 699700
rect 347832 699660 347838 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 321462 696940 321468 696992
rect 321520 696980 321526 696992
rect 580166 696980 580172 696992
rect 321520 696952 580172 696980
rect 321520 696940 321526 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 364610 687760 364616 687812
rect 364668 687800 364674 687812
rect 365162 687800 365168 687812
rect 364668 687772 365168 687800
rect 364668 687760 364674 687772
rect 365162 687760 365168 687772
rect 365220 687760 365226 687812
rect 429212 685936 429976 685964
rect 324222 685856 324228 685908
rect 324280 685896 324286 685908
rect 429212 685896 429240 685936
rect 324280 685868 429240 685896
rect 429948 685896 429976 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 429948 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 324280 685856 324286 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 364521 685831 364579 685837
rect 364521 685797 364533 685831
rect 364567 685828 364579 685831
rect 364610 685828 364616 685840
rect 364567 685800 364616 685828
rect 364567 685797 364579 685800
rect 364521 685791 364579 685797
rect 364610 685788 364616 685800
rect 364668 685788 364674 685840
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429565 684471 429623 684477
rect 429565 684468 429577 684471
rect 429344 684440 429577 684468
rect 429344 684428 429350 684440
rect 429565 684437 429577 684440
rect 429611 684437 429623 684471
rect 429565 684431 429623 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 382274 681748 382280 681760
rect 3568 681720 382280 681748
rect 3568 681708 3574 681720
rect 382274 681708 382280 681720
rect 382332 681708 382338 681760
rect 364518 676240 364524 676252
rect 364479 676212 364524 676240
rect 364518 676200 364524 676212
rect 364576 676200 364582 676252
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 320082 673480 320088 673532
rect 320140 673520 320146 673532
rect 580166 673520 580172 673532
rect 320140 673492 580172 673520
rect 320140 673480 320146 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 386414 667944 386420 667956
rect 3476 667916 386420 667944
rect 3476 667904 3482 667916
rect 386414 667904 386420 667916
rect 386472 667904 386478 667956
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 383654 652780 383660 652792
rect 3108 652752 383660 652780
rect 3108 652740 3114 652752
rect 383654 652740 383660 652752
rect 383712 652740 383718 652792
rect 315942 650020 315948 650072
rect 316000 650060 316006 650072
rect 580166 650060 580172 650072
rect 316000 650032 580172 650060
rect 316000 650020 316006 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 317322 638936 317328 638988
rect 317380 638976 317386 638988
rect 580166 638976 580172 638988
rect 317380 638948 580172 638976
rect 317380 638936 317386 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 313182 626560 313188 626612
rect 313240 626600 313246 626612
rect 580166 626600 580172 626612
rect 313240 626572 580172 626600
rect 313240 626560 313246 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 387794 623812 387800 623824
rect 3476 623784 387800 623812
rect 3476 623772 3482 623784
rect 387794 623772 387800 623784
rect 387852 623772 387858 623824
rect 364521 618239 364579 618245
rect 364521 618205 364533 618239
rect 364567 618236 364579 618239
rect 364610 618236 364616 618248
rect 364567 618208 364616 618236
rect 364567 618205 364579 618208
rect 364521 618199 364579 618205
rect 364610 618196 364616 618208
rect 364668 618196 364674 618248
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 391934 610008 391940 610020
rect 3476 609980 391940 610008
rect 3476 609968 3482 609980
rect 391934 609968 391940 609980
rect 391992 609968 391998 610020
rect 364518 608648 364524 608660
rect 364479 608620 364524 608648
rect 364518 608608 364524 608620
rect 364576 608608 364582 608660
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 309042 603100 309048 603152
rect 309100 603140 309106 603152
rect 580166 603140 580172 603152
rect 309100 603112 580172 603140
rect 309100 603100 309106 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 364610 598924 364616 598936
rect 364571 598896 364616 598924
rect 364610 598884 364616 598896
rect 364668 598884 364674 598936
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 390554 594844 390560 594856
rect 3292 594816 390560 594844
rect 3292 594804 3298 594816
rect 390554 594804 390560 594816
rect 390612 594804 390618 594856
rect 311802 592016 311808 592068
rect 311860 592056 311866 592068
rect 580166 592056 580172 592068
rect 311860 592028 580172 592056
rect 311860 592016 311866 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 364613 589339 364671 589345
rect 364613 589305 364625 589339
rect 364659 589336 364671 589339
rect 364702 589336 364708 589348
rect 364659 589308 364708 589336
rect 364659 589305 364671 589308
rect 364613 589299 364671 589305
rect 364702 589296 364708 589308
rect 364760 589296 364766 589348
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 344462 584672 344468 584724
rect 344520 584712 344526 584724
rect 364702 584712 364708 584724
rect 344520 584684 364708 584712
rect 344520 584672 344526 584684
rect 364702 584672 364708 584684
rect 364760 584672 364766 584724
rect 300762 584604 300768 584656
rect 300820 584644 300826 584656
rect 350810 584644 350816 584656
rect 300820 584616 350816 584644
rect 300820 584604 300826 584616
rect 350810 584604 350816 584616
rect 350868 584604 350874 584656
rect 338206 584536 338212 584588
rect 338264 584576 338270 584588
rect 429654 584576 429660 584588
rect 338264 584548 429660 584576
rect 338264 584536 338270 584548
rect 429654 584536 429660 584548
rect 429712 584536 429718 584588
rect 331858 584468 331864 584520
rect 331916 584508 331922 584520
rect 494238 584508 494244 584520
rect 331916 584480 494244 584508
rect 331916 584468 331922 584480
rect 494238 584468 494244 584480
rect 494296 584468 494302 584520
rect 325510 584400 325516 584452
rect 325568 584440 325574 584452
rect 559374 584440 559380 584452
rect 325568 584412 559380 584440
rect 325568 584400 325574 584412
rect 559374 584400 559380 584412
rect 559432 584400 559438 584452
rect 304534 583652 304540 583704
rect 304592 583692 304598 583704
rect 471238 583692 471244 583704
rect 304592 583664 471244 583692
rect 304592 583652 304598 583664
rect 471238 583652 471244 583664
rect 471296 583652 471302 583704
rect 298186 583584 298192 583636
rect 298244 583624 298250 583636
rect 469766 583624 469772 583636
rect 298244 583596 469772 583624
rect 298244 583584 298250 583596
rect 469766 583584 469772 583596
rect 469824 583584 469830 583636
rect 262398 583516 262404 583568
rect 262456 583556 262462 583568
rect 580718 583556 580724 583568
rect 262456 583528 580724 583556
rect 262456 583516 262462 583528
rect 580718 583516 580724 583528
rect 580776 583516 580782 583568
rect 256050 583448 256056 583500
rect 256108 583488 256114 583500
rect 580442 583488 580448 583500
rect 256108 583460 580448 583488
rect 256108 583448 256114 583460
rect 580442 583448 580448 583460
rect 580500 583448 580506 583500
rect 251818 583380 251824 583432
rect 251876 583420 251882 583432
rect 580350 583420 580356 583432
rect 251876 583392 580356 583420
rect 251876 583380 251882 583392
rect 580350 583380 580356 583392
rect 580408 583380 580414 583432
rect 6638 583312 6644 583364
rect 6696 583352 6702 583364
rect 399202 583352 399208 583364
rect 6696 583324 399208 583352
rect 6696 583312 6702 583324
rect 399202 583312 399208 583324
rect 399260 583312 399266 583364
rect 6362 583244 6368 583296
rect 6420 583284 6426 583296
rect 403434 583284 403440 583296
rect 6420 583256 403440 583284
rect 6420 583244 6426 583256
rect 403434 583244 403440 583256
rect 403492 583244 403498 583296
rect 4706 583176 4712 583228
rect 4764 583216 4770 583228
rect 405550 583216 405556 583228
rect 4764 583188 405556 583216
rect 4764 583176 4770 583188
rect 405550 583176 405556 583188
rect 405608 583176 405614 583228
rect 5350 583108 5356 583160
rect 5408 583148 5414 583160
rect 409782 583148 409788 583160
rect 5408 583120 409788 583148
rect 5408 583108 5414 583120
rect 409782 583108 409788 583120
rect 409840 583108 409846 583160
rect 3234 583040 3240 583092
rect 3292 583080 3298 583092
rect 407666 583080 407672 583092
rect 3292 583052 407672 583080
rect 3292 583040 3298 583052
rect 407666 583040 407672 583052
rect 407724 583040 407730 583092
rect 5442 582972 5448 583024
rect 5500 583012 5506 583024
rect 411898 583012 411904 583024
rect 5500 582984 411904 583012
rect 5500 582972 5506 582984
rect 411898 582972 411904 582984
rect 411956 582972 411962 583024
rect 14458 582904 14464 582956
rect 14516 582944 14522 582956
rect 424502 582944 424508 582956
rect 14516 582916 424508 582944
rect 14516 582904 14522 582916
rect 424502 582904 424508 582916
rect 424560 582904 424566 582956
rect 5258 582836 5264 582888
rect 5316 582876 5322 582888
rect 418154 582876 418160 582888
rect 5316 582848 418160 582876
rect 5316 582836 5322 582848
rect 418154 582836 418160 582848
rect 418212 582836 418218 582888
rect 15838 582768 15844 582820
rect 15896 582808 15902 582820
rect 430850 582808 430856 582820
rect 15896 582780 430856 582808
rect 15896 582768 15902 582780
rect 430850 582768 430856 582780
rect 430908 582768 430914 582820
rect 4062 582700 4068 582752
rect 4120 582740 4126 582752
rect 422386 582740 422392 582752
rect 4120 582712 422392 582740
rect 4120 582700 4126 582712
rect 422386 582700 422392 582712
rect 422444 582700 422450 582752
rect 17218 582632 17224 582684
rect 17276 582672 17282 582684
rect 437106 582672 437112 582684
rect 17276 582644 437112 582672
rect 17276 582632 17282 582644
rect 437106 582632 437112 582644
rect 437164 582632 437170 582684
rect 24118 582564 24124 582616
rect 24176 582604 24182 582616
rect 449802 582604 449808 582616
rect 24176 582576 449808 582604
rect 24176 582564 24182 582576
rect 449802 582564 449808 582576
rect 449860 582564 449866 582616
rect 5166 582496 5172 582548
rect 5224 582536 5230 582548
rect 434990 582536 434996 582548
rect 5224 582508 434996 582536
rect 5224 582496 5230 582508
rect 434990 582496 434996 582508
rect 435048 582496 435054 582548
rect 3694 582428 3700 582480
rect 3752 582468 3758 582480
rect 443454 582468 443460 582480
rect 3752 582440 443460 582468
rect 3752 582428 3758 582440
rect 443454 582428 443460 582440
rect 443512 582428 443518 582480
rect 5074 582360 5080 582412
rect 5132 582400 5138 582412
rect 447686 582400 447692 582412
rect 5132 582372 447692 582400
rect 5132 582360 5138 582372
rect 447686 582360 447692 582372
rect 447744 582360 447750 582412
rect 302418 581544 302424 581596
rect 302476 581584 302482 581596
rect 469582 581584 469588 581596
rect 302476 581556 469588 581584
rect 302476 581544 302482 581556
rect 469582 581544 469588 581556
rect 469640 581544 469646 581596
rect 296070 581476 296076 581528
rect 296128 581516 296134 581528
rect 469674 581516 469680 581528
rect 296128 581488 469680 581516
rect 296128 581476 296134 581488
rect 469674 581476 469680 581488
rect 469732 581476 469738 581528
rect 289722 581408 289728 581460
rect 289780 581448 289786 581460
rect 470502 581448 470508 581460
rect 289780 581420 470508 581448
rect 289780 581408 289786 581420
rect 470502 581408 470508 581420
rect 470560 581408 470566 581460
rect 287606 581340 287612 581392
rect 287664 581380 287670 581392
rect 470410 581380 470416 581392
rect 287664 581352 470416 581380
rect 287664 581340 287670 581352
rect 470410 581340 470416 581352
rect 470468 581340 470474 581392
rect 283466 581272 283472 581324
rect 283524 581312 283530 581324
rect 470318 581312 470324 581324
rect 283524 581284 470324 581312
rect 283524 581272 283530 581284
rect 470318 581272 470324 581284
rect 470376 581272 470382 581324
rect 281350 581204 281356 581256
rect 281408 581244 281414 581256
rect 470134 581244 470140 581256
rect 281408 581216 470140 581244
rect 281408 581204 281414 581216
rect 470134 581204 470140 581216
rect 470192 581204 470198 581256
rect 275002 581136 275008 581188
rect 275060 581176 275066 581188
rect 470042 581176 470048 581188
rect 275060 581148 470048 581176
rect 275060 581136 275066 581148
rect 470042 581136 470048 581148
rect 470100 581136 470106 581188
rect 264514 581068 264520 581120
rect 264572 581108 264578 581120
rect 580902 581108 580908 581120
rect 264572 581080 580908 581108
rect 264572 581068 264578 581080
rect 580902 581068 580908 581080
rect 580960 581068 580966 581120
rect 258166 581000 258172 581052
rect 258224 581040 258230 581052
rect 580626 581040 580632 581052
rect 258224 581012 580632 581040
rect 258224 581000 258230 581012
rect 580626 581000 580632 581012
rect 580684 581000 580690 581052
rect 268654 580252 268660 580304
rect 268712 580292 268718 580304
rect 469858 580292 469864 580304
rect 268712 580264 469864 580292
rect 268712 580252 268718 580264
rect 469858 580252 469864 580264
rect 469916 580252 469922 580304
rect 306558 580184 306564 580236
rect 306616 580224 306622 580236
rect 580166 580224 580172 580236
rect 306616 580196 580172 580224
rect 306616 580184 306622 580196
rect 580166 580184 580172 580196
rect 580224 580184 580230 580236
rect 6730 580116 6736 580168
rect 6788 580156 6794 580168
rect 395062 580156 395068 580168
rect 6788 580128 395068 580156
rect 6788 580116 6794 580128
rect 395062 580116 395068 580128
rect 395120 580116 395126 580168
rect 6454 580048 6460 580100
rect 6512 580088 6518 580100
rect 401318 580088 401324 580100
rect 6512 580060 401324 580088
rect 6512 580048 6518 580060
rect 401318 580048 401324 580060
rect 401376 580048 401382 580100
rect 6270 579980 6276 580032
rect 6328 580020 6334 580032
rect 414106 580020 414112 580032
rect 6328 579992 414112 580020
rect 6328 579980 6334 579992
rect 414106 579980 414112 579992
rect 414164 579980 414170 580032
rect 3970 579912 3976 579964
rect 4028 579952 4034 579964
rect 426434 579952 426440 579964
rect 4028 579924 426440 579952
rect 4028 579912 4034 579924
rect 426434 579912 426440 579924
rect 426492 579912 426498 579964
rect 3786 579844 3792 579896
rect 3844 579884 3850 579896
rect 438854 579884 438860 579896
rect 3844 579856 438860 579884
rect 3844 579844 3850 579856
rect 438854 579844 438860 579856
rect 438912 579844 438918 579896
rect 4982 579776 4988 579828
rect 5040 579816 5046 579828
rect 451550 579816 451556 579828
rect 5040 579788 451556 579816
rect 5040 579776 5046 579788
rect 451550 579776 451556 579788
rect 451608 579776 451614 579828
rect 4890 579708 4896 579760
rect 4948 579748 4954 579760
rect 458266 579748 458272 579760
rect 4948 579720 458272 579748
rect 4948 579708 4954 579720
rect 458266 579708 458272 579720
rect 458324 579708 458330 579760
rect 6178 579640 6184 579692
rect 6236 579680 6242 579692
rect 464246 579680 464252 579692
rect 6236 579652 464252 579680
rect 6236 579640 6242 579652
rect 464246 579640 464252 579652
rect 464304 579640 464310 579692
rect 271138 579368 271144 579420
rect 271196 579408 271202 579420
rect 271196 579380 282224 579408
rect 271196 579368 271202 579380
rect 254118 579300 254124 579352
rect 254176 579300 254182 579352
rect 260650 579300 260656 579352
rect 260708 579300 260714 579352
rect 266814 579300 266820 579352
rect 266872 579300 266878 579352
rect 273162 579300 273168 579352
rect 273220 579300 273226 579352
rect 277302 579300 277308 579352
rect 277360 579300 277366 579352
rect 279602 579300 279608 579352
rect 279660 579300 279666 579352
rect 254136 578660 254164 579300
rect 260668 578728 260696 579300
rect 266832 578796 266860 579300
rect 273180 578864 273208 579300
rect 277320 578932 277348 579300
rect 279620 579000 279648 579300
rect 282196 579136 282224 579380
rect 285766 579300 285772 579352
rect 285824 579300 285830 579352
rect 292114 579340 292120 579352
rect 292075 579312 292120 579340
rect 292114 579300 292120 579312
rect 292172 579300 292178 579352
rect 396718 579340 396724 579352
rect 396679 579312 396724 579340
rect 396718 579300 396724 579312
rect 396776 579300 396782 579352
rect 415670 579340 415676 579352
rect 415631 579312 415676 579340
rect 415670 579300 415676 579312
rect 415728 579300 415734 579352
rect 428366 579340 428372 579352
rect 428327 579312 428372 579340
rect 428366 579300 428372 579312
rect 428424 579300 428430 579352
rect 441062 579340 441068 579352
rect 441023 579312 441068 579340
rect 441062 579300 441068 579312
rect 441120 579300 441126 579352
rect 453574 579340 453580 579352
rect 453535 579312 453580 579340
rect 453574 579300 453580 579312
rect 453632 579300 453638 579352
rect 455782 579340 455788 579352
rect 455743 579312 455788 579340
rect 455782 579300 455788 579312
rect 455840 579300 455846 579352
rect 285784 579204 285812 579300
rect 470226 579204 470232 579216
rect 285784 579176 470232 579204
rect 470226 579164 470232 579176
rect 470284 579164 470290 579216
rect 469950 579136 469956 579148
rect 282196 579108 469956 579136
rect 469950 579096 469956 579108
rect 470008 579096 470014 579148
rect 292117 579071 292175 579077
rect 292117 579037 292129 579071
rect 292163 579068 292175 579071
rect 579890 579068 579896 579080
rect 292163 579040 579896 579068
rect 292163 579037 292175 579040
rect 292117 579031 292175 579037
rect 579890 579028 579896 579040
rect 579948 579028 579954 579080
rect 580074 579000 580080 579012
rect 279620 578972 580080 579000
rect 580074 578960 580080 578972
rect 580132 578960 580138 579012
rect 579982 578932 579988 578944
rect 277320 578904 579988 578932
rect 579982 578892 579988 578904
rect 580040 578892 580046 578944
rect 580166 578864 580172 578876
rect 273180 578836 580172 578864
rect 580166 578824 580172 578836
rect 580224 578824 580230 578876
rect 580810 578796 580816 578808
rect 266832 578768 580816 578796
rect 580810 578756 580816 578768
rect 580868 578756 580874 578808
rect 580534 578728 580540 578740
rect 260668 578700 580540 578728
rect 580534 578688 580540 578700
rect 580592 578688 580598 578740
rect 580258 578660 580264 578672
rect 254136 578632 580264 578660
rect 580258 578620 580264 578632
rect 580316 578620 580322 578672
rect 6546 578552 6552 578604
rect 6604 578592 6610 578604
rect 396721 578595 396779 578601
rect 396721 578592 396733 578595
rect 6604 578564 396733 578592
rect 6604 578552 6610 578564
rect 396721 578561 396733 578564
rect 396767 578561 396779 578595
rect 396721 578555 396779 578561
rect 3326 578484 3332 578536
rect 3384 578524 3390 578536
rect 415673 578527 415731 578533
rect 415673 578524 415685 578527
rect 3384 578496 415685 578524
rect 3384 578484 3390 578496
rect 415673 578493 415685 578496
rect 415719 578493 415731 578527
rect 415673 578487 415731 578493
rect 3878 578416 3884 578468
rect 3936 578456 3942 578468
rect 428369 578459 428427 578465
rect 428369 578456 428381 578459
rect 3936 578428 428381 578456
rect 3936 578416 3942 578428
rect 428369 578425 428381 578428
rect 428415 578425 428427 578459
rect 428369 578419 428427 578425
rect 3602 578348 3608 578400
rect 3660 578388 3666 578400
rect 441065 578391 441123 578397
rect 441065 578388 441077 578391
rect 3660 578360 441077 578388
rect 3660 578348 3666 578360
rect 441065 578357 441077 578360
rect 441111 578357 441123 578391
rect 441065 578351 441123 578357
rect 3418 578280 3424 578332
rect 3476 578320 3482 578332
rect 453577 578323 453635 578329
rect 453577 578320 453589 578323
rect 3476 578292 453589 578320
rect 3476 578280 3482 578292
rect 453577 578289 453589 578292
rect 453623 578289 453635 578323
rect 453577 578283 453635 578289
rect 3510 578212 3516 578264
rect 3568 578252 3574 578264
rect 455785 578255 455843 578261
rect 455785 578252 455797 578255
rect 3568 578224 455797 578252
rect 3568 578212 3574 578224
rect 455785 578221 455797 578224
rect 455831 578221 455843 578255
rect 455785 578215 455843 578221
rect 3142 568284 3148 568336
rect 3200 568324 3206 568336
rect 6730 568324 6736 568336
rect 3200 568296 6736 568324
rect 3200 568284 3206 568296
rect 6730 568284 6736 568296
rect 6788 568284 6794 568336
rect 579798 567128 579804 567180
rect 579856 567168 579862 567180
rect 580902 567168 580908 567180
rect 579856 567140 580908 567168
rect 579856 567128 579862 567140
rect 580902 567128 580908 567140
rect 580960 567128 580966 567180
rect 579798 557608 579804 557660
rect 579856 557648 579862 557660
rect 579856 557620 580948 557648
rect 579856 557608 579862 557620
rect 580920 557592 580948 557620
rect 580902 557540 580908 557592
rect 580960 557540 580966 557592
rect 469582 557472 469588 557524
rect 469640 557512 469646 557524
rect 579798 557512 579804 557524
rect 469640 557484 579804 557512
rect 469640 557472 469646 557484
rect 579798 557472 579804 557484
rect 579856 557472 579862 557524
rect 3142 553324 3148 553376
rect 3200 553364 3206 553376
rect 6638 553364 6644 553376
rect 3200 553336 6644 553364
rect 3200 553324 3206 553336
rect 6638 553324 6644 553336
rect 6696 553324 6702 553376
rect 579706 547816 579712 547868
rect 579764 547856 579770 547868
rect 580902 547856 580908 547868
rect 579764 547828 580908 547856
rect 579764 547816 579770 547828
rect 580902 547816 580908 547828
rect 580960 547816 580966 547868
rect 471238 546388 471244 546440
rect 471296 546428 471302 546440
rect 579798 546428 579804 546440
rect 471296 546400 579804 546428
rect 471296 546388 471302 546400
rect 579798 546388 579804 546400
rect 579856 546388 579862 546440
rect 3050 539044 3056 539096
rect 3108 539084 3114 539096
rect 6546 539084 6552 539096
rect 3108 539056 6552 539084
rect 3108 539044 3114 539056
rect 6546 539044 6552 539056
rect 6604 539044 6610 539096
rect 579706 538228 579712 538280
rect 579764 538268 579770 538280
rect 580902 538268 580908 538280
rect 579764 538240 580908 538268
rect 579764 538228 579770 538240
rect 580902 538228 580908 538240
rect 580960 538228 580966 538280
rect 579798 528504 579804 528556
rect 579856 528544 579862 528556
rect 580902 528544 580908 528556
rect 579856 528516 580908 528544
rect 579856 528504 579862 528516
rect 580902 528504 580908 528516
rect 580960 528504 580966 528556
rect 579798 518916 579804 518968
rect 579856 518956 579862 518968
rect 580902 518956 580908 518968
rect 579856 518928 580908 518956
rect 579856 518916 579862 518928
rect 580902 518916 580908 518928
rect 580960 518916 580966 518968
rect 469674 510552 469680 510604
rect 469732 510592 469738 510604
rect 579798 510592 579804 510604
rect 469732 510564 579804 510592
rect 469732 510552 469738 510564
rect 579798 510552 579804 510564
rect 579856 510552 579862 510604
rect 3142 510212 3148 510264
rect 3200 510252 3206 510264
rect 6454 510252 6460 510264
rect 3200 510224 6460 510252
rect 3200 510212 3206 510224
rect 6454 510212 6460 510224
rect 6512 510212 6518 510264
rect 579798 509192 579804 509244
rect 579856 509232 579862 509244
rect 580902 509232 580908 509244
rect 579856 509204 580908 509232
rect 579856 509192 579862 509204
rect 580902 509192 580908 509204
rect 580960 509192 580966 509244
rect 579798 499604 579804 499656
rect 579856 499644 579862 499656
rect 579856 499616 580948 499644
rect 579856 499604 579862 499616
rect 580920 499588 580948 499616
rect 580902 499536 580908 499588
rect 580960 499536 580966 499588
rect 469766 499468 469772 499520
rect 469824 499508 469830 499520
rect 579798 499508 579804 499520
rect 469824 499480 579804 499508
rect 469824 499468 469830 499480
rect 579798 499468 579804 499480
rect 579856 499468 579862 499520
rect 2774 495728 2780 495780
rect 2832 495768 2838 495780
rect 4706 495768 4712 495780
rect 2832 495740 4712 495768
rect 2832 495728 2838 495740
rect 4706 495728 4712 495740
rect 4764 495728 4770 495780
rect 579798 489812 579804 489864
rect 579856 489852 579862 489864
rect 580902 489852 580908 489864
rect 579856 489824 580908 489852
rect 579856 489812 579862 489824
rect 580902 489812 580908 489824
rect 580960 489812 580966 489864
rect 3142 481244 3148 481296
rect 3200 481284 3206 481296
rect 6362 481284 6368 481296
rect 3200 481256 6368 481284
rect 3200 481244 3206 481256
rect 6362 481244 6368 481256
rect 6420 481244 6426 481296
rect 579798 480224 579804 480276
rect 579856 480264 579862 480276
rect 580902 480264 580908 480276
rect 579856 480236 580908 480264
rect 579856 480224 579862 480236
rect 580902 480224 580908 480236
rect 580960 480224 580966 480276
rect 579706 470500 579712 470552
rect 579764 470540 579770 470552
rect 580902 470540 580908 470552
rect 579764 470512 580908 470540
rect 579764 470500 579770 470512
rect 580902 470500 580908 470512
rect 580960 470500 580966 470552
rect 470502 463632 470508 463684
rect 470560 463672 470566 463684
rect 579798 463672 579804 463684
rect 470560 463644 579804 463672
rect 470560 463632 470566 463644
rect 579798 463632 579804 463644
rect 579856 463632 579862 463684
rect 579706 460912 579712 460964
rect 579764 460952 579770 460964
rect 580902 460952 580908 460964
rect 579764 460924 580908 460952
rect 579764 460912 579770 460924
rect 580902 460912 580908 460924
rect 580960 460912 580966 460964
rect 470410 440172 470416 440224
rect 470468 440212 470474 440224
rect 579890 440212 579896 440224
rect 470468 440184 579896 440212
rect 470468 440172 470474 440184
rect 579890 440172 579896 440184
rect 579948 440172 579954 440224
rect 2774 438540 2780 438592
rect 2832 438580 2838 438592
rect 5442 438580 5448 438592
rect 2832 438552 5448 438580
rect 2832 438540 2838 438552
rect 5442 438540 5448 438552
rect 5500 438540 5506 438592
rect 2774 424804 2780 424856
rect 2832 424844 2838 424856
rect 5350 424844 5356 424856
rect 2832 424816 5356 424844
rect 2832 424804 2838 424816
rect 5350 424804 5356 424816
rect 5408 424804 5414 424856
rect 470318 416712 470324 416764
rect 470376 416752 470382 416764
rect 579890 416752 579896 416764
rect 470376 416724 579896 416752
rect 470376 416712 470382 416724
rect 579890 416712 579896 416724
rect 579948 416712 579954 416764
rect 579798 412564 579804 412616
rect 579856 412604 579862 412616
rect 580902 412604 580908 412616
rect 579856 412576 580908 412604
rect 579856 412564 579862 412576
rect 580902 412564 580908 412576
rect 580960 412564 580966 412616
rect 470226 405628 470232 405680
rect 470284 405668 470290 405680
rect 579890 405668 579896 405680
rect 470284 405640 579896 405668
rect 470284 405628 470290 405640
rect 579890 405628 579896 405640
rect 579948 405628 579954 405680
rect 579798 402976 579804 403028
rect 579856 403016 579862 403028
rect 580902 403016 580908 403028
rect 579856 402988 580908 403016
rect 579856 402976 579862 402988
rect 580902 402976 580908 402988
rect 580960 402976 580966 403028
rect 3234 395836 3240 395888
rect 3292 395876 3298 395888
rect 6270 395876 6276 395888
rect 3292 395848 6276 395876
rect 3292 395836 3298 395848
rect 6270 395836 6276 395848
rect 6328 395836 6334 395888
rect 470134 393252 470140 393304
rect 470192 393292 470198 393304
rect 579890 393292 579896 393304
rect 470192 393264 579896 393292
rect 470192 393252 470198 393264
rect 579890 393252 579896 393264
rect 579948 393252 579954 393304
rect 580902 393292 580908 393304
rect 580000 393264 580908 393292
rect 579798 393184 579804 393236
rect 579856 393224 579862 393236
rect 580000 393224 580028 393264
rect 580902 393252 580908 393264
rect 580960 393252 580966 393304
rect 579856 393196 580028 393224
rect 579856 393184 579862 393196
rect 579798 384276 579804 384328
rect 579856 384316 579862 384328
rect 580902 384316 580908 384328
rect 579856 384288 580908 384316
rect 579856 384276 579862 384288
rect 580902 384276 580908 384288
rect 580960 384276 580966 384328
rect 2774 380740 2780 380792
rect 2832 380780 2838 380792
rect 5258 380780 5264 380792
rect 2832 380752 5264 380780
rect 2832 380740 2838 380752
rect 5258 380740 5264 380752
rect 5316 380740 5322 380792
rect 579982 361224 579988 361276
rect 580040 361264 580046 361276
rect 580902 361264 580908 361276
rect 580040 361236 580908 361264
rect 580040 361224 580046 361236
rect 580902 361224 580908 361236
rect 580960 361224 580966 361276
rect 579798 360136 579804 360188
rect 579856 360176 579862 360188
rect 579982 360176 579988 360188
rect 579856 360148 579988 360176
rect 579856 360136 579862 360148
rect 579982 360136 579988 360148
rect 580040 360136 580046 360188
rect 470042 346332 470048 346384
rect 470100 346372 470106 346384
rect 579798 346372 579804 346384
rect 470100 346344 579804 346372
rect 470100 346332 470106 346344
rect 579798 346332 579804 346344
rect 579856 346332 579862 346384
rect 580074 345040 580080 345092
rect 580132 345080 580138 345092
rect 580902 345080 580908 345092
rect 580132 345052 580908 345080
rect 580132 345040 580138 345052
rect 580902 345040 580908 345052
rect 580960 345040 580966 345092
rect 580074 344904 580080 344956
rect 580132 344944 580138 344956
rect 580902 344944 580908 344956
rect 580132 344916 580908 344944
rect 580132 344904 580138 344916
rect 580902 344904 580908 344916
rect 580960 344904 580966 344956
rect 336737 338827 336795 338833
rect 336737 338793 336749 338827
rect 336783 338824 336795 338827
rect 341610 338824 341616 338836
rect 336783 338796 341616 338824
rect 336783 338793 336795 338796
rect 336737 338787 336795 338793
rect 341610 338784 341616 338796
rect 341668 338784 341674 338836
rect 346397 338691 346455 338697
rect 346397 338657 346409 338691
rect 346443 338688 346455 338691
rect 348510 338688 348516 338700
rect 346443 338660 348516 338688
rect 346443 338657 346455 338660
rect 346397 338651 346455 338657
rect 348510 338648 348516 338660
rect 348568 338648 348574 338700
rect 327350 338376 327356 338428
rect 327408 338416 327414 338428
rect 327902 338416 327908 338428
rect 327408 338388 327908 338416
rect 327408 338376 327414 338388
rect 327902 338376 327908 338388
rect 327960 338376 327966 338428
rect 287057 338147 287115 338153
rect 287057 338113 287069 338147
rect 287103 338144 287115 338147
rect 296625 338147 296683 338153
rect 296625 338144 296637 338147
rect 287103 338116 296637 338144
rect 287103 338113 287115 338116
rect 287057 338107 287115 338113
rect 296625 338113 296637 338116
rect 296671 338113 296683 338147
rect 296625 338107 296683 338113
rect 306377 338147 306435 338153
rect 306377 338113 306389 338147
rect 306423 338144 306435 338147
rect 315945 338147 316003 338153
rect 315945 338144 315957 338147
rect 306423 338116 315957 338144
rect 306423 338113 306435 338116
rect 306377 338107 306435 338113
rect 315945 338113 315957 338116
rect 315991 338113 316003 338147
rect 315945 338107 316003 338113
rect 342809 338147 342867 338153
rect 342809 338113 342821 338147
rect 342855 338144 342867 338147
rect 344649 338147 344707 338153
rect 344649 338144 344661 338147
rect 342855 338116 344661 338144
rect 342855 338113 342867 338116
rect 342809 338107 342867 338113
rect 344649 338113 344661 338116
rect 344695 338113 344707 338147
rect 344649 338107 344707 338113
rect 79318 338036 79324 338088
rect 79376 338076 79382 338088
rect 257890 338076 257896 338088
rect 79376 338048 257896 338076
rect 79376 338036 79382 338048
rect 257890 338036 257896 338048
rect 257948 338036 257954 338088
rect 309778 338036 309784 338088
rect 309836 338076 309842 338088
rect 354398 338076 354404 338088
rect 309836 338048 354404 338076
rect 309836 338036 309842 338048
rect 354398 338036 354404 338048
rect 354456 338036 354462 338088
rect 358078 338036 358084 338088
rect 358136 338076 358142 338088
rect 371510 338076 371516 338088
rect 358136 338048 371516 338076
rect 358136 338036 358142 338048
rect 371510 338036 371516 338048
rect 371568 338036 371574 338088
rect 372249 338079 372307 338085
rect 372249 338045 372261 338079
rect 372295 338076 372307 338079
rect 378870 338076 378876 338088
rect 372295 338048 378876 338076
rect 372295 338045 372307 338048
rect 372249 338039 372307 338045
rect 378870 338036 378876 338048
rect 378928 338036 378934 338088
rect 411254 338036 411260 338088
rect 411312 338076 411318 338088
rect 412450 338076 412456 338088
rect 411312 338048 412456 338076
rect 411312 338036 411318 338048
rect 412450 338036 412456 338048
rect 412508 338036 412514 338088
rect 414658 338036 414664 338088
rect 414716 338076 414722 338088
rect 429838 338076 429844 338088
rect 414716 338048 429844 338076
rect 414716 338036 414722 338048
rect 429838 338036 429844 338048
rect 429896 338036 429902 338088
rect 435726 338036 435732 338088
rect 435784 338076 435790 338088
rect 499574 338076 499580 338088
rect 435784 338048 499580 338076
rect 435784 338036 435790 338048
rect 499574 338036 499580 338048
rect 499632 338036 499638 338088
rect 71038 337968 71044 338020
rect 71096 338008 71102 338020
rect 252002 338008 252008 338020
rect 71096 337980 252008 338008
rect 71096 337968 71102 337980
rect 252002 337968 252008 337980
rect 252060 337968 252066 338020
rect 278777 338011 278835 338017
rect 278777 337977 278789 338011
rect 278823 338008 278835 338011
rect 287057 338011 287115 338017
rect 287057 338008 287069 338011
rect 278823 337980 287069 338008
rect 278823 337977 278835 337980
rect 278777 337971 278835 337977
rect 287057 337977 287069 337980
rect 287103 337977 287115 338011
rect 287057 337971 287115 337977
rect 306190 337968 306196 338020
rect 306248 338008 306254 338020
rect 355870 338008 355876 338020
rect 306248 337980 355876 338008
rect 306248 337968 306254 337980
rect 355870 337968 355876 337980
rect 355928 337968 355934 338020
rect 364242 337968 364248 338020
rect 364300 338008 364306 338020
rect 379330 338008 379336 338020
rect 364300 337980 379336 338008
rect 364300 337968 364306 337980
rect 379330 337968 379336 337980
rect 379388 337968 379394 338020
rect 399478 337968 399484 338020
rect 399536 338008 399542 338020
rect 400122 338008 400128 338020
rect 399536 337980 400128 338008
rect 399536 337968 399542 337980
rect 400122 337968 400128 337980
rect 400180 337968 400186 338020
rect 403342 337968 403348 338020
rect 403400 338008 403406 338020
rect 412545 338011 412603 338017
rect 412545 338008 412557 338011
rect 403400 337980 412557 338008
rect 403400 337968 403406 337980
rect 412545 337977 412557 337980
rect 412591 337977 412603 338011
rect 412545 337971 412603 337977
rect 415118 337968 415124 338020
rect 415176 338008 415182 338020
rect 420270 338008 420276 338020
rect 415176 337980 420276 338008
rect 415176 337968 415182 337980
rect 420270 337968 420276 337980
rect 420328 337968 420334 338020
rect 420546 337968 420552 338020
rect 420604 338008 420610 338020
rect 422297 338011 422355 338017
rect 422297 338008 422309 338011
rect 420604 337980 422309 338008
rect 420604 337968 420610 337980
rect 422297 337977 422309 337980
rect 422343 337977 422355 338011
rect 440142 338008 440148 338020
rect 440103 337980 440148 338008
rect 422297 337971 422355 337977
rect 440142 337968 440148 337980
rect 440200 337968 440206 338020
rect 451093 338011 451151 338017
rect 451093 337977 451105 338011
rect 451139 338008 451151 338011
rect 454681 338011 454739 338017
rect 454681 338008 454693 338011
rect 451139 337980 454693 338008
rect 451139 337977 451151 337980
rect 451093 337971 451151 337977
rect 454681 337977 454693 337980
rect 454727 337977 454739 338011
rect 454681 337971 454739 337977
rect 454770 337968 454776 338020
rect 454828 338008 454834 338020
rect 469125 338011 469183 338017
rect 469125 338008 469137 338011
rect 454828 337980 469137 338008
rect 454828 337968 454834 337980
rect 469125 337977 469137 337980
rect 469171 337977 469183 338011
rect 469125 337971 469183 337977
rect 469217 338011 469275 338017
rect 469217 337977 469229 338011
rect 469263 338008 469275 338011
rect 527818 338008 527824 338020
rect 469263 337980 527824 338008
rect 469263 337977 469275 337980
rect 469217 337971 469275 337977
rect 527818 337968 527824 337980
rect 527876 337968 527882 338020
rect 66898 337900 66904 337952
rect 66956 337940 66962 337952
rect 247126 337940 247132 337952
rect 66956 337912 247132 337940
rect 66956 337900 66962 337912
rect 247126 337900 247132 337912
rect 247184 337900 247190 337952
rect 303154 337900 303160 337952
rect 303212 337940 303218 337952
rect 327169 337943 327227 337949
rect 327169 337940 327181 337943
rect 303212 337912 327181 337940
rect 303212 337900 303218 337912
rect 327169 337909 327181 337912
rect 327215 337909 327227 337943
rect 327169 337903 327227 337909
rect 327261 337943 327319 337949
rect 327261 337909 327273 337943
rect 327307 337940 327319 337943
rect 352926 337940 352932 337952
rect 327307 337912 352932 337940
rect 327307 337909 327319 337912
rect 327261 337903 327319 337909
rect 352926 337900 352932 337912
rect 352984 337900 352990 337952
rect 355318 337900 355324 337952
rect 355376 337940 355382 337952
rect 370038 337940 370044 337952
rect 355376 337912 370044 337940
rect 355376 337900 355382 337912
rect 370038 337900 370044 337912
rect 370096 337900 370102 337952
rect 371142 337900 371148 337952
rect 371200 337940 371206 337952
rect 382274 337940 382280 337952
rect 371200 337912 382280 337940
rect 371200 337900 371206 337912
rect 382274 337900 382280 337912
rect 382332 337900 382338 337952
rect 409230 337900 409236 337952
rect 409288 337940 409294 337952
rect 416038 337940 416044 337952
rect 409288 337912 416044 337940
rect 409288 337900 409294 337912
rect 416038 337900 416044 337912
rect 416096 337900 416102 337952
rect 416590 337900 416596 337952
rect 416648 337940 416654 337952
rect 421558 337940 421564 337952
rect 416648 337912 421564 337940
rect 416648 337900 416654 337912
rect 421558 337900 421564 337912
rect 421616 337900 421622 337952
rect 422018 337900 422024 337952
rect 422076 337940 422082 337952
rect 438118 337940 438124 337952
rect 422076 337912 438124 337940
rect 422076 337900 422082 337912
rect 438118 337900 438124 337912
rect 438176 337900 438182 337952
rect 438670 337900 438676 337952
rect 438728 337940 438734 337952
rect 440237 337943 440295 337949
rect 440237 337940 440249 337943
rect 438728 337912 440249 337940
rect 438728 337900 438734 337912
rect 440237 337909 440249 337912
rect 440283 337909 440295 337943
rect 440237 337903 440295 337909
rect 440329 337943 440387 337949
rect 440329 337909 440341 337943
rect 440375 337940 440387 337943
rect 441893 337943 441951 337949
rect 441893 337940 441905 337943
rect 440375 337912 441905 337940
rect 440375 337909 440387 337912
rect 440329 337903 440387 337909
rect 441893 337909 441905 337912
rect 441939 337909 441951 337943
rect 441893 337903 441951 337909
rect 441985 337943 442043 337949
rect 441985 337909 441997 337943
rect 442031 337940 442043 337943
rect 449158 337940 449164 337952
rect 442031 337912 449164 337940
rect 442031 337909 442043 337912
rect 441985 337903 442043 337909
rect 449158 337900 449164 337912
rect 449216 337900 449222 337952
rect 450446 337900 450452 337952
rect 450504 337940 450510 337952
rect 451182 337940 451188 337952
rect 450504 337912 451188 337940
rect 450504 337900 450510 337912
rect 451182 337900 451188 337912
rect 451240 337900 451246 337952
rect 451826 337900 451832 337952
rect 451884 337940 451890 337952
rect 461581 337943 461639 337949
rect 461581 337940 461593 337943
rect 451884 337912 461593 337940
rect 451884 337900 451890 337912
rect 461581 337909 461593 337912
rect 461627 337909 461639 337943
rect 461581 337903 461639 337909
rect 461673 337943 461731 337949
rect 461673 337909 461685 337943
rect 461719 337940 461731 337943
rect 463421 337943 463479 337949
rect 463421 337940 463433 337943
rect 461719 337912 463433 337940
rect 461719 337909 461731 337912
rect 461673 337903 461731 337909
rect 463421 337909 463433 337912
rect 463467 337909 463479 337943
rect 525058 337940 525064 337952
rect 463421 337903 463479 337909
rect 463528 337912 525064 337940
rect 61378 337832 61384 337884
rect 61436 337872 61442 337884
rect 247586 337872 247592 337884
rect 61436 337844 247592 337872
rect 61436 337832 61442 337844
rect 247586 337832 247592 337844
rect 247644 337832 247650 337884
rect 258810 337832 258816 337884
rect 258868 337872 258874 337884
rect 272610 337872 272616 337884
rect 258868 337844 272616 337872
rect 258868 337832 258874 337844
rect 272610 337832 272616 337844
rect 272668 337832 272674 337884
rect 296625 337875 296683 337881
rect 296625 337841 296637 337875
rect 296671 337872 296683 337875
rect 306377 337875 306435 337881
rect 306377 337872 306389 337875
rect 296671 337844 306389 337872
rect 296671 337841 296683 337844
rect 296625 337835 296683 337841
rect 306377 337841 306389 337844
rect 306423 337841 306435 337875
rect 306377 337835 306435 337841
rect 315945 337875 316003 337881
rect 315945 337841 315957 337875
rect 315991 337872 316003 337875
rect 317414 337872 317420 337884
rect 315991 337844 317420 337872
rect 315991 337841 316003 337844
rect 315945 337835 316003 337841
rect 317414 337832 317420 337844
rect 317472 337832 317478 337884
rect 326982 337832 326988 337884
rect 327040 337872 327046 337884
rect 327077 337875 327135 337881
rect 327077 337872 327089 337875
rect 327040 337844 327089 337872
rect 327040 337832 327046 337844
rect 327077 337841 327089 337844
rect 327123 337841 327135 337875
rect 327077 337835 327135 337841
rect 336090 337832 336096 337884
rect 336148 337872 336154 337884
rect 344554 337872 344560 337884
rect 336148 337844 344560 337872
rect 336148 337832 336154 337844
rect 344554 337832 344560 337844
rect 344612 337832 344618 337884
rect 344649 337875 344707 337881
rect 344649 337841 344661 337875
rect 344695 337872 344707 337875
rect 349982 337872 349988 337884
rect 344695 337844 349988 337872
rect 344695 337841 344707 337844
rect 344649 337835 344707 337841
rect 349982 337832 349988 337844
rect 350040 337832 350046 337884
rect 365622 337872 365628 337884
rect 355336 337844 365628 337872
rect 57238 337764 57244 337816
rect 57296 337804 57302 337816
rect 244182 337804 244188 337816
rect 57296 337776 244188 337804
rect 57296 337764 57302 337776
rect 244182 337764 244188 337776
rect 244240 337764 244246 337816
rect 259638 337764 259644 337816
rect 259696 337804 259702 337816
rect 260098 337804 260104 337816
rect 259696 337776 260104 337804
rect 259696 337764 259702 337776
rect 260098 337764 260104 337776
rect 260156 337764 260162 337816
rect 275281 337807 275339 337813
rect 275281 337773 275293 337807
rect 275327 337804 275339 337807
rect 278777 337807 278835 337813
rect 278777 337804 278789 337807
rect 275327 337776 278789 337804
rect 275327 337773 275339 337776
rect 275281 337767 275339 337773
rect 278777 337773 278789 337776
rect 278823 337773 278835 337807
rect 278777 337767 278835 337773
rect 288250 337764 288256 337816
rect 288308 337804 288314 337816
rect 307021 337807 307079 337813
rect 288308 337776 302096 337804
rect 288308 337764 288314 337776
rect 35158 337696 35164 337748
rect 35216 337736 35222 337748
rect 238294 337736 238300 337748
rect 35216 337708 238300 337736
rect 35216 337696 35222 337708
rect 238294 337696 238300 337708
rect 238352 337696 238358 337748
rect 254578 337696 254584 337748
rect 254636 337736 254642 337748
rect 262306 337736 262312 337748
rect 254636 337708 262312 337736
rect 254636 337696 254642 337708
rect 262306 337696 262312 337708
rect 262364 337696 262370 337748
rect 302068 337736 302096 337776
rect 307021 337773 307033 337807
rect 307067 337804 307079 337807
rect 351914 337804 351920 337816
rect 307067 337776 351920 337804
rect 307067 337773 307079 337776
rect 307021 337767 307079 337773
rect 351914 337764 351920 337776
rect 351972 337764 351978 337816
rect 327166 337736 327172 337748
rect 302068 337708 327172 337736
rect 327166 337696 327172 337708
rect 327224 337696 327230 337748
rect 336182 337696 336188 337748
rect 336240 337736 336246 337748
rect 346397 337739 346455 337745
rect 346397 337736 346409 337739
rect 336240 337708 346409 337736
rect 336240 337696 336246 337708
rect 346397 337705 346409 337708
rect 346443 337705 346455 337739
rect 346397 337699 346455 337705
rect 39298 337628 39304 337680
rect 39356 337668 39362 337680
rect 244642 337668 244648 337680
rect 39356 337640 244648 337668
rect 39356 337628 39362 337640
rect 244642 337628 244648 337640
rect 244700 337628 244706 337680
rect 260098 337628 260104 337680
rect 260156 337668 260162 337680
rect 277026 337668 277032 337680
rect 260156 337640 277032 337668
rect 260156 337628 260162 337640
rect 277026 337628 277032 337640
rect 277084 337628 277090 337680
rect 285582 337628 285588 337680
rect 285640 337668 285646 337680
rect 347038 337668 347044 337680
rect 285640 337640 347044 337668
rect 285640 337628 285646 337640
rect 347038 337628 347044 337640
rect 347096 337628 347102 337680
rect 348418 337628 348424 337680
rect 348476 337668 348482 337680
rect 355336 337668 355364 337844
rect 365622 337832 365628 337844
rect 365680 337832 365686 337884
rect 366913 337875 366971 337881
rect 366913 337841 366925 337875
rect 366959 337872 366971 337875
rect 380802 337872 380808 337884
rect 366959 337844 380808 337872
rect 366959 337841 366971 337844
rect 366913 337835 366971 337841
rect 380802 337832 380808 337844
rect 380860 337832 380866 337884
rect 388438 337832 388444 337884
rect 388496 337872 388502 337884
rect 389174 337872 389180 337884
rect 388496 337844 389180 337872
rect 388496 337832 388502 337844
rect 389174 337832 389180 337844
rect 389232 337832 389238 337884
rect 397454 337832 397460 337884
rect 397512 337872 397518 337884
rect 399478 337872 399484 337884
rect 397512 337844 399484 337872
rect 397512 337832 397518 337844
rect 399478 337832 399484 337844
rect 399536 337832 399542 337884
rect 399938 337832 399944 337884
rect 399996 337872 400002 337884
rect 412818 337872 412824 337884
rect 399996 337844 412824 337872
rect 399996 337832 400002 337844
rect 412818 337832 412824 337844
rect 412876 337832 412882 337884
rect 413646 337832 413652 337884
rect 413704 337872 413710 337884
rect 417418 337872 417424 337884
rect 413704 337844 417424 337872
rect 413704 337832 413710 337844
rect 417418 337832 417424 337844
rect 417476 337832 417482 337884
rect 417602 337832 417608 337884
rect 417660 337872 417666 337884
rect 455598 337872 455604 337884
rect 417660 337844 455604 337872
rect 417660 337832 417666 337844
rect 455598 337832 455604 337844
rect 455656 337832 455662 337884
rect 458726 337832 458732 337884
rect 458784 337872 458790 337884
rect 459370 337872 459376 337884
rect 458784 337844 459376 337872
rect 458784 337832 458790 337844
rect 459370 337832 459376 337844
rect 459428 337832 459434 337884
rect 460658 337832 460664 337884
rect 460716 337872 460722 337884
rect 463528 337872 463556 337912
rect 525058 337900 525064 337912
rect 525116 337900 525122 337952
rect 460716 337844 463556 337872
rect 463605 337875 463663 337881
rect 460716 337832 460722 337844
rect 463605 337841 463617 337875
rect 463651 337872 463663 337875
rect 523678 337872 523684 337884
rect 463651 337844 523684 337872
rect 463651 337841 463663 337844
rect 463605 337835 463663 337841
rect 523678 337832 523684 337844
rect 523736 337832 523742 337884
rect 358722 337764 358728 337816
rect 358780 337804 358786 337816
rect 358780 337776 360884 337804
rect 358780 337764 358786 337776
rect 348476 337640 355364 337668
rect 348476 337628 348482 337640
rect 356698 337628 356704 337680
rect 356756 337668 356762 337680
rect 360746 337668 360752 337680
rect 356756 337640 360752 337668
rect 356756 337628 356762 337640
rect 360746 337628 360752 337640
rect 360804 337628 360810 337680
rect 360856 337668 360884 337776
rect 362862 337764 362868 337816
rect 362920 337804 362926 337816
rect 372249 337807 372307 337813
rect 372249 337804 372261 337807
rect 362920 337776 372261 337804
rect 362920 337764 362926 337776
rect 372249 337773 372261 337776
rect 372295 337773 372307 337807
rect 377398 337804 377404 337816
rect 372249 337767 372307 337773
rect 372356 337776 377404 337804
rect 361666 337696 361672 337748
rect 361724 337736 361730 337748
rect 362310 337736 362316 337748
rect 361724 337708 362316 337736
rect 361724 337696 361730 337708
rect 362310 337696 362316 337708
rect 362368 337696 362374 337748
rect 363046 337696 363052 337748
rect 363104 337736 363110 337748
rect 363782 337736 363788 337748
rect 363104 337708 363788 337736
rect 363104 337696 363110 337708
rect 363782 337696 363788 337708
rect 363840 337696 363846 337748
rect 372356 337736 372384 337776
rect 377398 337764 377404 337776
rect 377456 337764 377462 337816
rect 398006 337764 398012 337816
rect 398064 337804 398070 337816
rect 399570 337804 399576 337816
rect 398064 337776 399576 337804
rect 398064 337764 398070 337776
rect 399570 337764 399576 337776
rect 399628 337764 399634 337816
rect 401870 337764 401876 337816
rect 401928 337804 401934 337816
rect 416958 337804 416964 337816
rect 401928 337776 416964 337804
rect 401928 337764 401934 337776
rect 416958 337764 416964 337776
rect 417016 337764 417022 337816
rect 419994 337764 420000 337816
rect 420052 337804 420058 337816
rect 420730 337804 420736 337816
rect 420052 337776 420736 337804
rect 420052 337764 420058 337776
rect 420730 337764 420736 337776
rect 420788 337764 420794 337816
rect 424962 337764 424968 337816
rect 425020 337804 425026 337816
rect 442258 337804 442264 337816
rect 425020 337776 442264 337804
rect 425020 337764 425026 337776
rect 442258 337764 442264 337776
rect 442316 337764 442322 337816
rect 444558 337764 444564 337816
rect 444616 337804 444622 337816
rect 445662 337804 445668 337816
rect 444616 337776 445668 337804
rect 444616 337764 444622 337776
rect 445662 337764 445668 337776
rect 445720 337764 445726 337816
rect 446030 337764 446036 337816
rect 446088 337804 446094 337816
rect 453209 337807 453267 337813
rect 453209 337804 453221 337807
rect 446088 337776 453221 337804
rect 446088 337764 446094 337776
rect 453209 337773 453221 337776
rect 453255 337773 453267 337807
rect 453209 337767 453267 337773
rect 453298 337764 453304 337816
rect 453356 337804 453362 337816
rect 453942 337804 453948 337816
rect 453356 337776 453948 337804
rect 453356 337764 453362 337776
rect 453942 337764 453948 337776
rect 454000 337764 454006 337816
rect 459005 337807 459063 337813
rect 459005 337773 459017 337807
rect 459051 337804 459063 337807
rect 463786 337804 463792 337816
rect 459051 337776 463792 337804
rect 459051 337773 459063 337776
rect 459005 337767 459063 337773
rect 463786 337764 463792 337776
rect 463844 337764 463850 337816
rect 465626 337764 465632 337816
rect 465684 337804 465690 337816
rect 466178 337804 466184 337816
rect 465684 337776 466184 337804
rect 465684 337764 465690 337776
rect 466178 337764 466184 337776
rect 466236 337764 466242 337816
rect 467098 337764 467104 337816
rect 467156 337804 467162 337816
rect 467742 337804 467748 337816
rect 467156 337776 467748 337804
rect 467156 337764 467162 337776
rect 467742 337764 467748 337776
rect 467800 337764 467806 337816
rect 468018 337764 468024 337816
rect 468076 337804 468082 337816
rect 469030 337804 469036 337816
rect 468076 337776 469036 337804
rect 468076 337764 468082 337776
rect 469030 337764 469036 337776
rect 469088 337764 469094 337816
rect 469125 337807 469183 337813
rect 469125 337773 469137 337807
rect 469171 337804 469183 337807
rect 521010 337804 521016 337816
rect 469171 337776 521016 337804
rect 469171 337773 469183 337776
rect 469125 337767 469183 337773
rect 521010 337764 521016 337776
rect 521068 337764 521074 337816
rect 375926 337736 375932 337748
rect 363892 337708 372384 337736
rect 372448 337708 375932 337736
rect 363892 337668 363920 337708
rect 360856 337640 363920 337668
rect 363969 337671 364027 337677
rect 363969 337637 363981 337671
rect 364015 337668 364027 337671
rect 372448 337668 372476 337708
rect 375926 337696 375932 337708
rect 375984 337696 375990 337748
rect 380158 337696 380164 337748
rect 380216 337736 380222 337748
rect 381354 337736 381360 337748
rect 380216 337708 381360 337736
rect 380216 337696 380222 337708
rect 381354 337696 381360 337708
rect 381412 337696 381418 337748
rect 381538 337696 381544 337748
rect 381596 337736 381602 337748
rect 382826 337736 382832 337748
rect 381596 337708 382832 337736
rect 381596 337696 381602 337708
rect 382826 337696 382832 337708
rect 382884 337696 382890 337748
rect 384942 337696 384948 337748
rect 385000 337736 385006 337748
rect 388162 337736 388168 337748
rect 385000 337708 388168 337736
rect 385000 337696 385006 337708
rect 388162 337696 388168 337708
rect 388220 337696 388226 337748
rect 408770 337696 408776 337748
rect 408828 337736 408834 337748
rect 409782 337736 409788 337748
rect 408828 337708 409788 337736
rect 408828 337696 408834 337708
rect 409782 337696 409788 337708
rect 409840 337696 409846 337748
rect 412468 337708 413600 337736
rect 381814 337668 381820 337680
rect 364015 337640 372476 337668
rect 373828 337640 381820 337668
rect 364015 337637 364027 337640
rect 363969 337631 364027 337637
rect 32398 337560 32404 337612
rect 32456 337600 32462 337612
rect 241698 337600 241704 337612
rect 32456 337572 241704 337600
rect 32456 337560 32462 337572
rect 241698 337560 241704 337572
rect 241756 337560 241762 337612
rect 252186 337560 252192 337612
rect 252244 337600 252250 337612
rect 256418 337600 256424 337612
rect 252244 337572 256424 337600
rect 252244 337560 252250 337572
rect 256418 337560 256424 337572
rect 256476 337560 256482 337612
rect 261386 337560 261392 337612
rect 261444 337600 261450 337612
rect 279970 337600 279976 337612
rect 261444 337572 279976 337600
rect 261444 337560 261450 337572
rect 279970 337560 279976 337572
rect 280028 337560 280034 337612
rect 281442 337560 281448 337612
rect 281500 337600 281506 337612
rect 345290 337600 345296 337612
rect 281500 337572 345296 337600
rect 281500 337560 281506 337572
rect 345290 337560 345296 337572
rect 345348 337560 345354 337612
rect 345569 337603 345627 337609
rect 345569 337569 345581 337603
rect 345615 337600 345627 337603
rect 351454 337600 351460 337612
rect 345615 337572 351460 337600
rect 345615 337569 345627 337572
rect 345569 337563 345627 337569
rect 351454 337560 351460 337572
rect 351512 337560 351518 337612
rect 351638 337560 351644 337612
rect 351696 337600 351702 337612
rect 368201 337603 368259 337609
rect 368201 337600 368213 337603
rect 351696 337572 368213 337600
rect 351696 337560 351702 337572
rect 368201 337569 368213 337572
rect 368247 337569 368259 337603
rect 368201 337563 368259 337569
rect 369118 337560 369124 337612
rect 369176 337600 369182 337612
rect 371050 337600 371056 337612
rect 369176 337572 371056 337600
rect 369176 337560 369182 337572
rect 371050 337560 371056 337572
rect 371108 337560 371114 337612
rect 28258 337492 28264 337544
rect 28316 337532 28322 337544
rect 28316 337504 234476 337532
rect 28316 337492 28322 337504
rect 19978 337424 19984 337476
rect 20036 337464 20042 337476
rect 234338 337464 234344 337476
rect 20036 337436 234344 337464
rect 20036 337424 20042 337436
rect 234338 337424 234344 337436
rect 234396 337424 234402 337476
rect 234448 337464 234476 337504
rect 253198 337492 253204 337544
rect 253256 337532 253262 337544
rect 259362 337532 259368 337544
rect 253256 337504 259368 337532
rect 253256 337492 253262 337504
rect 259362 337492 259368 337504
rect 259420 337492 259426 337544
rect 275554 337532 275560 337544
rect 260300 337504 275560 337532
rect 237834 337464 237840 337476
rect 234448 337436 237840 337464
rect 237834 337424 237840 337436
rect 237892 337424 237898 337476
rect 258718 337424 258724 337476
rect 258776 337464 258782 337476
rect 260300 337464 260328 337504
rect 275554 337492 275560 337504
rect 275612 337492 275618 337544
rect 275922 337492 275928 337544
rect 275980 337532 275986 337544
rect 327169 337535 327227 337541
rect 327169 337532 327181 337535
rect 275980 337504 327181 337532
rect 275980 337492 275986 337504
rect 327169 337501 327181 337504
rect 327215 337501 327227 337535
rect 327169 337495 327227 337501
rect 341705 337535 341763 337541
rect 341705 337501 341717 337535
rect 341751 337532 341763 337535
rect 342809 337535 342867 337541
rect 342809 337532 342821 337535
rect 341751 337504 342821 337532
rect 341751 337501 341763 337504
rect 341705 337495 341763 337501
rect 342809 337501 342821 337504
rect 342855 337501 342867 337535
rect 342809 337495 342867 337501
rect 342898 337492 342904 337544
rect 342956 337532 342962 337544
rect 353386 337532 353392 337544
rect 342956 337504 353392 337532
rect 342956 337492 342962 337504
rect 353386 337492 353392 337504
rect 353444 337492 353450 337544
rect 353941 337535 353999 337541
rect 353941 337501 353953 337535
rect 353987 337532 353999 337535
rect 357342 337532 357348 337544
rect 353987 337504 357348 337532
rect 353987 337501 353999 337504
rect 353941 337495 353999 337501
rect 357342 337492 357348 337504
rect 357400 337492 357406 337544
rect 359458 337492 359464 337544
rect 359516 337532 359522 337544
rect 363690 337532 363696 337544
rect 359516 337504 363696 337532
rect 359516 337492 359522 337504
rect 363690 337492 363696 337504
rect 363748 337492 363754 337544
rect 269666 337464 269672 337476
rect 258776 337436 260328 337464
rect 260392 337436 269672 337464
rect 258776 337424 258782 337436
rect 13078 337356 13084 337408
rect 13136 337396 13142 337408
rect 233510 337396 233516 337408
rect 13136 337368 233516 337396
rect 13136 337356 13142 337368
rect 233510 337356 233516 337368
rect 233568 337356 233574 337408
rect 233878 337356 233884 337408
rect 233936 337396 233942 337408
rect 241238 337396 241244 337408
rect 233936 337368 241244 337396
rect 233936 337356 233942 337368
rect 241238 337356 241244 337368
rect 241296 337356 241302 337408
rect 247678 337356 247684 337408
rect 247736 337396 247742 337408
rect 248598 337396 248604 337408
rect 247736 337368 248604 337396
rect 247736 337356 247742 337368
rect 248598 337356 248604 337368
rect 248656 337356 248662 337408
rect 249058 337356 249064 337408
rect 249116 337396 249122 337408
rect 250530 337396 250536 337408
rect 249116 337368 250536 337396
rect 249116 337356 249122 337368
rect 250530 337356 250536 337368
rect 250588 337356 250594 337408
rect 250714 337356 250720 337408
rect 250772 337396 250778 337408
rect 253474 337396 253480 337408
rect 250772 337368 253480 337396
rect 250772 337356 250778 337368
rect 253474 337356 253480 337368
rect 253532 337356 253538 337408
rect 257338 337356 257344 337408
rect 257396 337396 257402 337408
rect 260392 337396 260420 337436
rect 269666 337424 269672 337436
rect 269724 337424 269730 337476
rect 297910 337424 297916 337476
rect 297968 337464 297974 337476
rect 307021 337467 307079 337473
rect 307021 337464 307033 337467
rect 297968 337436 307033 337464
rect 297968 337424 297974 337436
rect 307021 337433 307033 337436
rect 307067 337433 307079 337467
rect 307021 337427 307079 337433
rect 314654 337424 314660 337476
rect 314712 337464 314718 337476
rect 315390 337464 315396 337476
rect 314712 337436 315396 337464
rect 314712 337424 314718 337436
rect 315390 337424 315396 337436
rect 315448 337424 315454 337476
rect 316126 337424 316132 337476
rect 316184 337464 316190 337476
rect 316310 337464 316316 337476
rect 316184 337436 316316 337464
rect 316184 337424 316190 337436
rect 316310 337424 316316 337436
rect 316368 337424 316374 337476
rect 317414 337424 317420 337476
rect 317472 337464 317478 337476
rect 318334 337464 318340 337476
rect 317472 337436 318340 337464
rect 317472 337424 317478 337436
rect 318334 337424 318340 337436
rect 318392 337424 318398 337476
rect 318886 337424 318892 337476
rect 318944 337464 318950 337476
rect 319254 337464 319260 337476
rect 318944 337436 319260 337464
rect 318944 337424 318950 337436
rect 319254 337424 319260 337436
rect 319312 337424 319318 337476
rect 320174 337424 320180 337476
rect 320232 337464 320238 337476
rect 320726 337464 320732 337476
rect 320232 337436 320732 337464
rect 320232 337424 320238 337436
rect 320726 337424 320732 337436
rect 320784 337424 320790 337476
rect 327077 337467 327135 337473
rect 327077 337433 327089 337467
rect 327123 337464 327135 337467
rect 336737 337467 336795 337473
rect 336737 337464 336749 337467
rect 327123 337436 336749 337464
rect 327123 337433 327135 337436
rect 327077 337427 327135 337433
rect 336737 337433 336749 337436
rect 336783 337433 336795 337467
rect 336737 337427 336795 337433
rect 338758 337424 338764 337476
rect 338816 337464 338822 337476
rect 347498 337464 347504 337476
rect 338816 337436 347504 337464
rect 338816 337424 338822 337436
rect 347498 337424 347504 337436
rect 347556 337424 347562 337476
rect 349062 337424 349068 337476
rect 349120 337464 349126 337476
rect 372982 337464 372988 337476
rect 349120 337436 372988 337464
rect 349120 337424 349126 337436
rect 372982 337424 372988 337436
rect 373040 337424 373046 337476
rect 266722 337396 266728 337408
rect 257396 337368 260420 337396
rect 260944 337368 266728 337396
rect 257396 337356 257402 337368
rect 77938 337288 77944 337340
rect 77996 337328 78002 337340
rect 77996 337300 84700 337328
rect 77996 337288 78002 337300
rect 84672 337192 84700 337300
rect 84838 337288 84844 337340
rect 84896 337328 84902 337340
rect 260834 337328 260840 337340
rect 84896 337300 260840 337328
rect 84896 337288 84902 337300
rect 260834 337288 260840 337300
rect 260892 337288 260898 337340
rect 108945 337263 109003 337269
rect 108945 337229 108957 337263
rect 108991 337260 109003 337263
rect 113177 337263 113235 337269
rect 113177 337260 113189 337263
rect 108991 337232 113189 337260
rect 108991 337229 109003 337232
rect 108945 337223 109003 337229
rect 113177 337229 113189 337232
rect 113223 337229 113235 337263
rect 113177 337223 113235 337229
rect 122745 337263 122803 337269
rect 122745 337229 122757 337263
rect 122791 337260 122803 337263
rect 132494 337260 132500 337272
rect 122791 337232 132500 337260
rect 122791 337229 122803 337232
rect 122745 337223 122803 337229
rect 132494 337220 132500 337232
rect 132552 337220 132558 337272
rect 142062 337220 142068 337272
rect 142120 337260 142126 337272
rect 151814 337260 151820 337272
rect 142120 337232 151820 337260
rect 142120 337220 142126 337232
rect 151814 337220 151820 337232
rect 151872 337220 151878 337272
rect 161382 337220 161388 337272
rect 161440 337260 161446 337272
rect 171134 337260 171140 337272
rect 161440 337232 171140 337260
rect 161440 337220 161446 337232
rect 171134 337220 171140 337232
rect 171192 337220 171198 337272
rect 180702 337220 180708 337272
rect 180760 337260 180766 337272
rect 190454 337260 190460 337272
rect 180760 337232 190460 337260
rect 180760 337220 180766 337232
rect 190454 337220 190460 337232
rect 190512 337220 190518 337272
rect 200022 337220 200028 337272
rect 200080 337260 200086 337272
rect 209774 337260 209780 337272
rect 200080 337232 209780 337260
rect 200080 337220 200086 337232
rect 209774 337220 209780 337232
rect 209832 337220 209838 337272
rect 219342 337220 219348 337272
rect 219400 337260 219406 337272
rect 229186 337260 229192 337272
rect 219400 337232 229192 337260
rect 219400 337220 219406 337232
rect 229186 337220 229192 337232
rect 229244 337220 229250 337272
rect 234614 337220 234620 337272
rect 234672 337260 234678 337272
rect 254946 337260 254952 337272
rect 234672 337232 254952 337260
rect 234672 337220 234678 337232
rect 254946 337220 254952 337232
rect 255004 337220 255010 337272
rect 255958 337220 255964 337272
rect 256016 337260 256022 337272
rect 260944 337260 260972 337368
rect 266722 337356 266728 337368
rect 266780 337356 266786 337408
rect 269022 337356 269028 337408
rect 269080 337396 269086 337408
rect 340230 337396 340236 337408
rect 269080 337368 340236 337396
rect 269080 337356 269086 337368
rect 340230 337356 340236 337368
rect 340288 337356 340294 337408
rect 340782 337356 340788 337408
rect 340840 337396 340846 337408
rect 369578 337396 369584 337408
rect 340840 337368 369584 337396
rect 340840 337356 340846 337368
rect 369578 337356 369584 337368
rect 369636 337356 369642 337408
rect 369762 337356 369768 337408
rect 369820 337396 369826 337408
rect 373828 337396 373856 337640
rect 381814 337628 381820 337640
rect 381872 337628 381878 337680
rect 384298 337628 384304 337680
rect 384356 337668 384362 337680
rect 387702 337668 387708 337680
rect 384356 337640 387708 337668
rect 384356 337628 384362 337640
rect 387702 337628 387708 337640
rect 387760 337628 387766 337680
rect 404354 337628 404360 337680
rect 404412 337668 404418 337680
rect 412468 337668 412496 337708
rect 404412 337640 412496 337668
rect 412545 337671 412603 337677
rect 404412 337628 404418 337640
rect 412545 337637 412557 337671
rect 412591 337668 412603 337671
rect 413465 337671 413523 337677
rect 413465 337668 413477 337671
rect 412591 337640 413477 337668
rect 412591 337637 412603 337640
rect 412545 337631 412603 337637
rect 413465 337637 413477 337640
rect 413511 337637 413523 337671
rect 413572 337668 413600 337708
rect 419534 337696 419540 337748
rect 419592 337736 419598 337748
rect 420822 337736 420828 337748
rect 419592 337708 420828 337736
rect 419592 337696 419598 337708
rect 420822 337696 420828 337708
rect 420880 337696 420886 337748
rect 421466 337696 421472 337748
rect 421524 337736 421530 337748
rect 422202 337736 422208 337748
rect 421524 337708 422208 337736
rect 421524 337696 421530 337708
rect 422202 337696 422208 337708
rect 422260 337696 422266 337748
rect 422478 337696 422484 337748
rect 422536 337736 422542 337748
rect 424410 337736 424416 337748
rect 422536 337708 424416 337736
rect 422536 337696 422542 337708
rect 424410 337696 424416 337708
rect 424468 337696 424474 337748
rect 425422 337696 425428 337748
rect 425480 337736 425486 337748
rect 428458 337736 428464 337748
rect 425480 337708 428464 337736
rect 425480 337696 425486 337708
rect 428458 337696 428464 337708
rect 428516 337696 428522 337748
rect 439130 337696 439136 337748
rect 439188 337736 439194 337748
rect 440142 337736 440148 337748
rect 439188 337708 440148 337736
rect 439188 337696 439194 337708
rect 440142 337696 440148 337708
rect 440200 337696 440206 337748
rect 440237 337739 440295 337745
rect 440237 337705 440249 337739
rect 440283 337736 440295 337739
rect 506474 337736 506480 337748
rect 440283 337708 506480 337736
rect 440283 337705 440295 337708
rect 440237 337699 440295 337705
rect 506474 337696 506480 337708
rect 506532 337696 506538 337748
rect 420178 337668 420184 337680
rect 413572 337640 420184 337668
rect 413465 337631 413523 337637
rect 420178 337628 420184 337640
rect 420236 337628 420242 337680
rect 427906 337628 427912 337680
rect 427964 337668 427970 337680
rect 441985 337671 442043 337677
rect 441985 337668 441997 337671
rect 427964 337640 441997 337668
rect 427964 337628 427970 337640
rect 441985 337637 441997 337640
rect 442031 337637 442043 337671
rect 441985 337631 442043 337637
rect 442074 337628 442080 337680
rect 442132 337668 442138 337680
rect 442902 337668 442908 337680
rect 442132 337640 442908 337668
rect 442132 337628 442138 337640
rect 442902 337628 442908 337640
rect 442960 337628 442966 337680
rect 443546 337628 443552 337680
rect 443604 337668 443610 337680
rect 444282 337668 444288 337680
rect 443604 337640 444288 337668
rect 443604 337628 443610 337640
rect 444282 337628 444288 337640
rect 444340 337628 444346 337680
rect 445018 337628 445024 337680
rect 445076 337668 445082 337680
rect 445570 337668 445576 337680
rect 445076 337640 445576 337668
rect 445076 337628 445082 337640
rect 445570 337628 445576 337640
rect 445628 337628 445634 337680
rect 446490 337628 446496 337680
rect 446548 337668 446554 337680
rect 447042 337668 447048 337680
rect 446548 337640 447048 337668
rect 446548 337628 446554 337640
rect 447042 337628 447048 337640
rect 447100 337628 447106 337680
rect 448238 337628 448244 337680
rect 448296 337668 448302 337680
rect 448422 337668 448428 337680
rect 448296 337640 448428 337668
rect 448296 337628 448302 337640
rect 448422 337628 448428 337640
rect 448480 337628 448486 337680
rect 449894 337628 449900 337680
rect 449952 337668 449958 337680
rect 450998 337668 451004 337680
rect 449952 337640 451004 337668
rect 449952 337628 449958 337640
rect 450998 337628 451004 337640
rect 451056 337628 451062 337680
rect 451366 337628 451372 337680
rect 451424 337668 451430 337680
rect 452470 337668 452476 337680
rect 451424 337640 452476 337668
rect 451424 337628 451430 337640
rect 452470 337628 452476 337640
rect 452528 337628 452534 337680
rect 452838 337628 452844 337680
rect 452896 337668 452902 337680
rect 453758 337668 453764 337680
rect 452896 337640 453764 337668
rect 452896 337628 452902 337640
rect 453758 337628 453764 337640
rect 453816 337628 453822 337680
rect 454310 337628 454316 337680
rect 454368 337668 454374 337680
rect 455230 337668 455236 337680
rect 454368 337640 455236 337668
rect 454368 337628 454374 337640
rect 455230 337628 455236 337640
rect 455288 337628 455294 337680
rect 455782 337628 455788 337680
rect 455840 337668 455846 337680
rect 456610 337668 456616 337680
rect 455840 337640 456616 337668
rect 455840 337628 455846 337640
rect 456610 337628 456616 337640
rect 456668 337628 456674 337680
rect 456794 337628 456800 337680
rect 456852 337668 456858 337680
rect 458082 337668 458088 337680
rect 456852 337640 458088 337668
rect 456852 337628 456858 337640
rect 458082 337628 458088 337640
rect 458140 337628 458146 337680
rect 458174 337628 458180 337680
rect 458232 337668 458238 337680
rect 461489 337671 461547 337677
rect 461489 337668 461501 337671
rect 458232 337640 461501 337668
rect 458232 337628 458238 337640
rect 461489 337637 461501 337640
rect 461535 337637 461547 337671
rect 461489 337631 461547 337637
rect 461581 337671 461639 337677
rect 461581 337637 461593 337671
rect 461627 337668 461639 337671
rect 520918 337668 520924 337680
rect 461627 337640 520924 337668
rect 461627 337637 461639 337640
rect 461581 337631 461639 337637
rect 520918 337628 520924 337640
rect 520976 337628 520982 337680
rect 373902 337560 373908 337612
rect 373960 337600 373966 337612
rect 383286 337600 383292 337612
rect 373960 337572 383292 337600
rect 373960 337560 373966 337572
rect 383286 337560 383292 337572
rect 383344 337560 383350 337612
rect 404814 337560 404820 337612
rect 404872 337600 404878 337612
rect 415489 337603 415547 337609
rect 415489 337600 415501 337603
rect 404872 337572 415501 337600
rect 404872 337560 404878 337572
rect 415489 337569 415501 337572
rect 415535 337569 415547 337603
rect 415489 337563 415547 337569
rect 415578 337560 415584 337612
rect 415636 337600 415642 337612
rect 416590 337600 416596 337612
rect 415636 337572 416596 337600
rect 415636 337560 415642 337572
rect 416590 337560 416596 337572
rect 416648 337560 416654 337612
rect 422297 337603 422355 337609
rect 422297 337569 422309 337603
rect 422343 337600 422355 337603
rect 422343 337572 426572 337600
rect 422343 337569 422355 337572
rect 422297 337563 422355 337569
rect 400398 337492 400404 337544
rect 400456 337532 400462 337544
rect 406378 337532 406384 337544
rect 400456 337504 406384 337532
rect 400456 337492 400462 337504
rect 406378 337492 406384 337504
rect 406436 337492 406442 337544
rect 407298 337492 407304 337544
rect 407356 337532 407362 337544
rect 426069 337535 426127 337541
rect 426069 337532 426081 337535
rect 407356 337504 426081 337532
rect 407356 337492 407362 337504
rect 426069 337501 426081 337504
rect 426115 337501 426127 337535
rect 426069 337495 426127 337501
rect 375282 337424 375288 337476
rect 375340 337464 375346 337476
rect 383746 337464 383752 337476
rect 375340 337436 383752 337464
rect 375340 337424 375346 337436
rect 383746 337424 383752 337436
rect 383804 337424 383810 337476
rect 387058 337424 387064 337476
rect 387116 337464 387122 337476
rect 388714 337464 388720 337476
rect 387116 337436 388720 337464
rect 387116 337424 387122 337436
rect 388714 337424 388720 337436
rect 388772 337424 388778 337476
rect 398466 337424 398472 337476
rect 398524 337464 398530 337476
rect 398524 337436 402376 337464
rect 398524 337424 398530 337436
rect 369820 337368 373856 337396
rect 369820 337356 369826 337368
rect 382182 337356 382188 337408
rect 382240 337396 382246 337408
rect 386690 337396 386696 337408
rect 382240 337368 386696 337396
rect 382240 337356 382246 337368
rect 386690 337356 386696 337368
rect 386748 337356 386754 337408
rect 400950 337356 400956 337408
rect 401008 337396 401014 337408
rect 402238 337396 402244 337408
rect 401008 337368 402244 337396
rect 401008 337356 401014 337368
rect 402238 337356 402244 337368
rect 402296 337356 402302 337408
rect 402348 337396 402376 337436
rect 405826 337424 405832 337476
rect 405884 337464 405890 337476
rect 426434 337464 426440 337476
rect 405884 337436 426440 337464
rect 405884 337424 405890 337436
rect 426434 337424 426440 337436
rect 426492 337424 426498 337476
rect 426544 337464 426572 337572
rect 430114 337560 430120 337612
rect 430172 337600 430178 337612
rect 435177 337603 435235 337609
rect 435177 337600 435189 337603
rect 430172 337572 435189 337600
rect 430172 337560 430178 337572
rect 435177 337569 435189 337572
rect 435223 337569 435235 337603
rect 435177 337563 435235 337569
rect 436646 337560 436652 337612
rect 436704 337600 436710 337612
rect 437290 337600 437296 337612
rect 436704 337572 437296 337600
rect 436704 337560 436710 337572
rect 437290 337560 437296 337572
rect 437348 337560 437354 337612
rect 437658 337560 437664 337612
rect 437716 337600 437722 337612
rect 438670 337600 438676 337612
rect 437716 337572 438676 337600
rect 437716 337560 437722 337572
rect 438670 337560 438676 337572
rect 438728 337560 438734 337612
rect 440602 337560 440608 337612
rect 440660 337600 440666 337612
rect 441522 337600 441528 337612
rect 440660 337572 441528 337600
rect 440660 337560 440666 337572
rect 441522 337560 441528 337572
rect 441580 337560 441586 337612
rect 441614 337560 441620 337612
rect 441672 337600 441678 337612
rect 443638 337600 443644 337612
rect 441672 337572 443644 337600
rect 441672 337560 441678 337572
rect 443638 337560 443644 337572
rect 443696 337560 443702 337612
rect 443748 337572 448652 337600
rect 427170 337492 427176 337544
rect 427228 337532 427234 337544
rect 432601 337535 432659 337541
rect 432601 337532 432613 337535
rect 427228 337504 432613 337532
rect 427228 337492 427234 337504
rect 432601 337501 432613 337504
rect 432647 337501 432659 337535
rect 432601 337495 432659 337501
rect 432693 337535 432751 337541
rect 432693 337501 432705 337535
rect 432739 337532 432751 337535
rect 437109 337535 437167 337541
rect 437109 337532 437121 337535
rect 432739 337504 437121 337532
rect 432739 337501 432751 337504
rect 432693 337495 432751 337501
rect 437109 337501 437121 337504
rect 437155 337501 437167 337535
rect 437109 337495 437167 337501
rect 437198 337492 437204 337544
rect 437256 337532 437262 337544
rect 442350 337532 442356 337544
rect 437256 337504 442356 337532
rect 437256 337492 437262 337504
rect 442350 337492 442356 337504
rect 442408 337492 442414 337544
rect 443748 337532 443776 337572
rect 442460 337504 443776 337532
rect 426544 337436 432644 337464
rect 408678 337396 408684 337408
rect 402348 337368 408684 337396
rect 408678 337356 408684 337368
rect 408736 337356 408742 337408
rect 411714 337356 411720 337408
rect 411772 337396 411778 337408
rect 431589 337399 431647 337405
rect 431589 337396 431601 337399
rect 411772 337368 431601 337396
rect 411772 337356 411778 337368
rect 431589 337365 431601 337368
rect 431635 337365 431647 337399
rect 432616 337396 432644 337436
rect 434254 337424 434260 337476
rect 434312 337464 434318 337476
rect 439498 337464 439504 337476
rect 434312 337436 439504 337464
rect 434312 337424 434318 337436
rect 439498 337424 439504 337436
rect 439556 337424 439562 337476
rect 441893 337467 441951 337473
rect 441893 337433 441905 337467
rect 441939 337464 441951 337467
rect 442460 337464 442488 337504
rect 447502 337492 447508 337544
rect 447560 337532 447566 337544
rect 448422 337532 448428 337544
rect 447560 337504 448428 337532
rect 447560 337492 447566 337504
rect 448422 337492 448428 337504
rect 448480 337492 448486 337544
rect 441939 337436 442488 337464
rect 441939 337433 441951 337436
rect 441893 337427 441951 337433
rect 443086 337424 443092 337476
rect 443144 337464 443150 337476
rect 448517 337467 448575 337473
rect 448517 337464 448529 337467
rect 443144 337436 448529 337464
rect 443144 337424 443150 337436
rect 448517 337433 448529 337436
rect 448563 337433 448575 337467
rect 448624 337464 448652 337572
rect 448974 337560 448980 337612
rect 449032 337600 449038 337612
rect 518158 337600 518164 337612
rect 449032 337572 518164 337600
rect 449032 337560 449038 337572
rect 518158 337560 518164 337572
rect 518216 337560 518222 337612
rect 448701 337535 448759 337541
rect 448701 337501 448713 337535
rect 448747 337532 448759 337535
rect 514018 337532 514024 337544
rect 448747 337504 514024 337532
rect 448747 337501 448759 337504
rect 448701 337495 448759 337501
rect 514018 337492 514024 337504
rect 514076 337492 514082 337544
rect 451093 337467 451151 337473
rect 451093 337464 451105 337467
rect 448624 337436 451105 337464
rect 448517 337427 448575 337433
rect 451093 337433 451105 337436
rect 451139 337433 451151 337467
rect 451093 337427 451151 337433
rect 453209 337467 453267 337473
rect 453209 337433 453221 337467
rect 453255 337464 453267 337467
rect 516778 337464 516784 337476
rect 453255 337436 516784 337464
rect 453255 337433 453267 337436
rect 453209 337427 453267 337433
rect 516778 337424 516784 337436
rect 516836 337424 516842 337476
rect 440329 337399 440387 337405
rect 440329 337396 440341 337399
rect 432616 337368 440341 337396
rect 431589 337359 431647 337365
rect 440329 337365 440341 337368
rect 440375 337365 440387 337399
rect 440329 337359 440387 337365
rect 446953 337399 447011 337405
rect 446953 337365 446965 337399
rect 446999 337396 447011 337399
rect 510614 337396 510620 337408
rect 446999 337368 510620 337396
rect 446999 337365 447011 337368
rect 446953 337359 447011 337365
rect 510614 337356 510620 337368
rect 510672 337356 510678 337408
rect 272794 337288 272800 337340
rect 272852 337328 272858 337340
rect 314194 337328 314200 337340
rect 272852 337300 314200 337328
rect 272852 337288 272858 337300
rect 314194 337288 314200 337300
rect 314252 337288 314258 337340
rect 316034 337288 316040 337340
rect 316092 337328 316098 337340
rect 316862 337328 316868 337340
rect 316092 337300 316868 337328
rect 316092 337288 316098 337300
rect 316862 337288 316868 337300
rect 316920 337288 316926 337340
rect 318794 337288 318800 337340
rect 318852 337328 318858 337340
rect 319806 337328 319812 337340
rect 318852 337300 319812 337328
rect 318852 337288 318858 337300
rect 319806 337288 319812 337300
rect 319864 337288 319870 337340
rect 321462 337288 321468 337340
rect 321520 337328 321526 337340
rect 361758 337328 361764 337340
rect 321520 337300 361764 337328
rect 321520 337288 321526 337300
rect 361758 337288 361764 337300
rect 361816 337288 361822 337340
rect 366910 337288 366916 337340
rect 366968 337328 366974 337340
rect 380342 337328 380348 337340
rect 366968 337300 380348 337328
rect 366968 337288 366974 337300
rect 380342 337288 380348 337300
rect 380400 337288 380406 337340
rect 396994 337288 397000 337340
rect 397052 337328 397058 337340
rect 405918 337328 405924 337340
rect 397052 337300 405924 337328
rect 397052 337288 397058 337300
rect 405918 337288 405924 337300
rect 405976 337288 405982 337340
rect 412726 337288 412732 337340
rect 412784 337328 412790 337340
rect 413830 337328 413836 337340
rect 412784 337300 413836 337328
rect 412784 337288 412790 337300
rect 413830 337288 413836 337300
rect 413888 337288 413894 337340
rect 418522 337288 418528 337340
rect 418580 337328 418586 337340
rect 419442 337328 419448 337340
rect 418580 337300 419448 337328
rect 418580 337288 418586 337300
rect 419442 337288 419448 337300
rect 419500 337288 419506 337340
rect 421006 337288 421012 337340
rect 421064 337328 421070 337340
rect 459005 337331 459063 337337
rect 459005 337328 459017 337331
rect 421064 337300 459017 337328
rect 421064 337288 421070 337300
rect 459005 337297 459017 337300
rect 459051 337297 459063 337331
rect 459005 337291 459063 337297
rect 459097 337331 459155 337337
rect 459097 337297 459109 337331
rect 459143 337328 459155 337331
rect 470594 337328 470600 337340
rect 459143 337300 470600 337328
rect 459143 337297 459155 337300
rect 459097 337291 459155 337297
rect 470594 337288 470600 337300
rect 470652 337288 470658 337340
rect 470686 337288 470692 337340
rect 470744 337328 470750 337340
rect 529198 337328 529204 337340
rect 470744 337300 529204 337328
rect 470744 337288 470750 337300
rect 529198 337288 529204 337300
rect 529256 337288 529262 337340
rect 256016 337232 260972 337260
rect 256016 337220 256022 337232
rect 271322 337220 271328 337272
rect 271380 337260 271386 337272
rect 312446 337260 312452 337272
rect 271380 337232 312452 337260
rect 271380 337220 271386 337232
rect 312446 337220 312452 337232
rect 312504 337220 312510 337272
rect 312538 337220 312544 337272
rect 312596 337260 312602 337272
rect 350442 337260 350448 337272
rect 312596 337232 350448 337260
rect 312596 337220 312602 337232
rect 350442 337220 350448 337232
rect 350500 337220 350506 337272
rect 350537 337263 350595 337269
rect 350537 337229 350549 337263
rect 350583 337260 350595 337263
rect 353941 337263 353999 337269
rect 353941 337260 353953 337263
rect 350583 337232 353953 337260
rect 350583 337229 350595 337232
rect 350537 337223 350595 337229
rect 353941 337229 353953 337232
rect 353987 337229 353999 337263
rect 353941 337223 353999 337229
rect 355962 337220 355968 337272
rect 356020 337260 356026 337272
rect 363969 337263 364027 337269
rect 363969 337260 363981 337263
rect 356020 337232 363981 337260
rect 356020 337220 356026 337232
rect 363969 337229 363981 337232
rect 364015 337229 364027 337263
rect 363969 337223 364027 337229
rect 414198 337220 414204 337272
rect 414256 337260 414262 337272
rect 415302 337260 415308 337272
rect 414256 337232 415308 337260
rect 414256 337220 414262 337232
rect 415302 337220 415308 337232
rect 415360 337220 415366 337272
rect 423490 337220 423496 337272
rect 423548 337260 423554 337272
rect 461581 337263 461639 337269
rect 461581 337260 461593 337263
rect 423548 337232 461593 337260
rect 423548 337220 423554 337232
rect 461581 337229 461593 337232
rect 461627 337229 461639 337263
rect 461581 337223 461639 337229
rect 463602 337220 463608 337272
rect 463660 337260 463666 337272
rect 469217 337263 469275 337269
rect 469217 337260 469229 337263
rect 463660 337232 469229 337260
rect 463660 337220 463666 337232
rect 469217 337229 469229 337232
rect 469263 337229 469275 337263
rect 469217 337223 469275 337229
rect 469490 337220 469496 337272
rect 469548 337260 469554 337272
rect 530578 337260 530584 337272
rect 469548 337232 530584 337260
rect 469548 337220 469554 337232
rect 530578 337220 530584 337232
rect 530636 337220 530642 337272
rect 84672 337164 94544 337192
rect 94516 337124 94544 337164
rect 97258 337152 97264 337204
rect 97316 337192 97322 337204
rect 268194 337192 268200 337204
rect 97316 337164 268200 337192
rect 97316 337152 97322 337164
rect 268194 337152 268200 337164
rect 268252 337152 268258 337204
rect 271782 337152 271788 337204
rect 271840 337192 271846 337204
rect 275281 337195 275339 337201
rect 275281 337192 275293 337195
rect 271840 337164 275293 337192
rect 271840 337152 271846 337164
rect 275281 337161 275293 337164
rect 275327 337161 275339 337195
rect 275281 337155 275339 337161
rect 333238 337152 333244 337204
rect 333296 337192 333302 337204
rect 366634 337192 366640 337204
rect 333296 337164 366640 337192
rect 333296 337152 333302 337164
rect 366634 337152 366640 337164
rect 366692 337152 366698 337204
rect 368201 337195 368259 337201
rect 368201 337161 368213 337195
rect 368247 337192 368259 337195
rect 372062 337192 372068 337204
rect 368247 337164 372068 337192
rect 368247 337161 368259 337164
rect 368201 337155 368259 337161
rect 372062 337152 372068 337164
rect 372120 337152 372126 337204
rect 415489 337195 415547 337201
rect 415489 337161 415501 337195
rect 415535 337192 415547 337195
rect 424318 337192 424324 337204
rect 415535 337164 424324 337192
rect 415535 337161 415547 337164
rect 415489 337155 415547 337161
rect 424318 337152 424324 337164
rect 424376 337152 424382 337204
rect 431494 337192 431500 337204
rect 425992 337164 431500 337192
rect 99377 337127 99435 337133
rect 99377 337124 99389 337127
rect 94516 337096 99389 337124
rect 99377 337093 99389 337096
rect 99423 337093 99435 337127
rect 99377 337087 99435 337093
rect 100662 337084 100668 337136
rect 100720 337124 100726 337136
rect 271138 337124 271144 337136
rect 100720 337096 271144 337124
rect 100720 337084 100726 337096
rect 271138 337084 271144 337096
rect 271196 337084 271202 337136
rect 316678 337084 316684 337136
rect 316736 337124 316742 337136
rect 341705 337127 341763 337133
rect 341705 337124 341717 337127
rect 316736 337096 341717 337124
rect 316736 337084 316742 337096
rect 341705 337093 341717 337096
rect 341751 337093 341763 337127
rect 341705 337087 341763 337093
rect 341886 337084 341892 337136
rect 341944 337124 341950 337136
rect 348970 337124 348976 337136
rect 341944 337096 348976 337124
rect 341944 337084 341950 337096
rect 348970 337084 348976 337096
rect 349028 337084 349034 337136
rect 351822 337084 351828 337136
rect 351880 337124 351886 337136
rect 374454 337124 374460 337136
rect 351880 337096 374460 337124
rect 351880 337084 351886 337096
rect 374454 337084 374460 337096
rect 374512 337084 374518 337136
rect 406286 337084 406292 337136
rect 406344 337124 406350 337136
rect 411898 337124 411904 337136
rect 406344 337096 411904 337124
rect 406344 337084 406350 337096
rect 411898 337084 411904 337096
rect 411956 337084 411962 337136
rect 417050 337084 417056 337136
rect 417108 337124 417114 337136
rect 417970 337124 417976 337136
rect 417108 337096 417976 337124
rect 417108 337084 417114 337096
rect 417970 337084 417976 337096
rect 418028 337084 418034 337136
rect 419074 337084 419080 337136
rect 419132 337124 419138 337136
rect 425992 337124 426020 337164
rect 431494 337152 431500 337164
rect 431552 337152 431558 337204
rect 431589 337195 431647 337201
rect 431589 337161 431601 337195
rect 431635 337192 431647 337195
rect 434070 337192 434076 337204
rect 431635 337164 434076 337192
rect 431635 337161 431647 337164
rect 431589 337155 431647 337161
rect 434070 337152 434076 337164
rect 434128 337152 434134 337204
rect 444377 337195 444435 337201
rect 444377 337192 444389 337195
rect 435100 337164 444389 337192
rect 419132 337096 426020 337124
rect 426069 337127 426127 337133
rect 419132 337084 419138 337096
rect 426069 337093 426081 337127
rect 426115 337124 426127 337127
rect 427078 337124 427084 337136
rect 426115 337096 427084 337124
rect 426115 337093 426127 337096
rect 426069 337087 426127 337093
rect 427078 337084 427084 337096
rect 427136 337084 427142 337136
rect 427817 337127 427875 337133
rect 427817 337093 427829 337127
rect 427863 337124 427875 337127
rect 432693 337127 432751 337133
rect 432693 337124 432705 337127
rect 427863 337096 432705 337124
rect 427863 337093 427875 337096
rect 427817 337087 427875 337093
rect 432693 337093 432705 337096
rect 432739 337093 432751 337127
rect 432693 337087 432751 337093
rect 432782 337084 432788 337136
rect 432840 337124 432846 337136
rect 435100 337124 435128 337164
rect 444377 337161 444389 337164
rect 444423 337161 444435 337195
rect 444377 337155 444435 337161
rect 444561 337195 444619 337201
rect 444561 337161 444573 337195
rect 444607 337192 444619 337195
rect 492674 337192 492680 337204
rect 444607 337164 492680 337192
rect 444607 337161 444619 337164
rect 444561 337155 444619 337161
rect 492674 337152 492680 337164
rect 492732 337152 492738 337204
rect 432840 337096 435128 337124
rect 435177 337127 435235 337133
rect 432840 337084 432846 337096
rect 435177 337093 435189 337127
rect 435223 337124 435235 337127
rect 444469 337127 444527 337133
rect 444469 337124 444481 337127
rect 435223 337096 444481 337124
rect 435223 337093 435235 337096
rect 435177 337087 435235 337093
rect 444469 337093 444481 337096
rect 444515 337093 444527 337127
rect 444469 337087 444527 337093
rect 444653 337127 444711 337133
rect 444653 337093 444665 337127
rect 444699 337124 444711 337127
rect 485774 337124 485780 337136
rect 444699 337096 485780 337124
rect 444699 337093 444711 337096
rect 444653 337087 444711 337093
rect 485774 337084 485780 337096
rect 485832 337084 485838 337136
rect 95878 337016 95884 337068
rect 95936 337056 95942 337068
rect 263778 337056 263784 337068
rect 95936 337028 263784 337056
rect 95936 337016 95942 337028
rect 263778 337016 263784 337028
rect 263836 337016 263842 337068
rect 335262 337016 335268 337068
rect 335320 337056 335326 337068
rect 367646 337056 367652 337068
rect 335320 337028 367652 337056
rect 335320 337016 335326 337028
rect 367646 337016 367652 337028
rect 367704 337016 367710 337068
rect 393590 337016 393596 337068
rect 393648 337056 393654 337068
rect 397454 337056 397460 337068
rect 393648 337028 397460 337056
rect 393648 337016 393654 337028
rect 397454 337016 397460 337028
rect 397512 337016 397518 337068
rect 401410 337016 401416 337068
rect 401468 337056 401474 337068
rect 404998 337056 405004 337068
rect 401468 337028 405004 337056
rect 401468 337016 401474 337028
rect 404998 337016 405004 337028
rect 405056 337016 405062 337068
rect 413465 337059 413523 337065
rect 413465 337025 413477 337059
rect 413511 337056 413523 337059
rect 421098 337056 421104 337068
rect 413511 337028 421104 337056
rect 413511 337025 413523 337028
rect 413465 337019 413523 337025
rect 421098 337016 421104 337028
rect 421156 337016 421162 337068
rect 432601 337059 432659 337065
rect 432601 337025 432613 337059
rect 432647 337056 432659 337059
rect 444374 337056 444380 337068
rect 432647 337028 444380 337056
rect 432647 337025 432659 337028
rect 432601 337019 432659 337025
rect 444374 337016 444380 337028
rect 444432 337016 444438 337068
rect 444742 337016 444748 337068
rect 444800 337056 444806 337068
rect 477586 337056 477592 337068
rect 444800 337028 477592 337056
rect 444800 337016 444806 337028
rect 477586 337016 477592 337028
rect 477644 337016 477650 337068
rect 107562 336948 107568 337000
rect 107620 336988 107626 337000
rect 274082 336988 274088 337000
rect 107620 336960 274088 336988
rect 107620 336948 107626 336960
rect 274082 336948 274088 336960
rect 274140 336948 274146 337000
rect 319438 336948 319444 337000
rect 319496 336988 319502 337000
rect 345569 336991 345627 336997
rect 345569 336988 345581 336991
rect 319496 336960 345581 336988
rect 319496 336948 319502 336960
rect 345569 336957 345581 336960
rect 345615 336957 345627 336991
rect 345569 336951 345627 336957
rect 378042 336948 378048 337000
rect 378100 336988 378106 337000
rect 385218 336988 385224 337000
rect 378100 336960 385224 336988
rect 378100 336948 378106 336960
rect 385218 336948 385224 336960
rect 385276 336948 385282 337000
rect 398926 336948 398932 337000
rect 398984 336988 398990 337000
rect 403618 336988 403624 337000
rect 398984 336960 403624 336988
rect 398984 336948 398990 336960
rect 403618 336948 403624 336960
rect 403676 336948 403682 337000
rect 407758 336948 407764 337000
rect 407816 336988 407822 337000
rect 407816 336960 411300 336988
rect 407816 336948 407822 336960
rect 102778 336880 102784 336932
rect 102836 336920 102842 336932
rect 265250 336920 265256 336932
rect 102836 336892 265256 336920
rect 102836 336880 102842 336892
rect 265250 336880 265256 336892
rect 265308 336880 265314 336932
rect 284294 336880 284300 336932
rect 284352 336920 284358 336932
rect 284846 336920 284852 336932
rect 284352 336892 284852 336920
rect 284352 336880 284358 336892
rect 284846 336880 284852 336892
rect 284904 336880 284910 336932
rect 327718 336880 327724 336932
rect 327776 336920 327782 336932
rect 345474 336920 345480 336932
rect 327776 336892 345480 336920
rect 327776 336880 327782 336892
rect 345474 336880 345480 336892
rect 345532 336880 345538 336932
rect 345658 336880 345664 336932
rect 345716 336920 345722 336932
rect 360286 336920 360292 336932
rect 345716 336892 360292 336920
rect 345716 336880 345722 336892
rect 360286 336880 360292 336892
rect 360344 336880 360350 336932
rect 380802 336880 380808 336932
rect 380860 336920 380866 336932
rect 386230 336920 386236 336932
rect 380860 336892 386236 336920
rect 380860 336880 380866 336892
rect 386230 336880 386236 336892
rect 386288 336880 386294 336932
rect 392118 336880 392124 336932
rect 392176 336920 392182 336932
rect 393590 336920 393596 336932
rect 392176 336892 393596 336920
rect 392176 336880 392182 336892
rect 393590 336880 393596 336892
rect 393648 336880 393654 336932
rect 410242 336880 410248 336932
rect 410300 336920 410306 336932
rect 411162 336920 411168 336932
rect 410300 336892 411168 336920
rect 410300 336880 410306 336892
rect 411162 336880 411168 336892
rect 411220 336880 411226 336932
rect 411272 336920 411300 336960
rect 426802 336948 426808 337000
rect 426860 336988 426866 337000
rect 444469 336991 444527 336997
rect 444469 336988 444481 336991
rect 426860 336960 444481 336988
rect 426860 336948 426866 336960
rect 444469 336957 444481 336960
rect 444515 336957 444527 336991
rect 444469 336951 444527 336957
rect 444561 336991 444619 336997
rect 444561 336957 444573 336991
rect 444607 336988 444619 336991
rect 475378 336988 475384 337000
rect 444607 336960 475384 336988
rect 444607 336957 444619 336960
rect 444561 336951 444619 336957
rect 475378 336948 475384 336960
rect 475436 336948 475442 337000
rect 413278 336920 413284 336932
rect 411272 336892 413284 336920
rect 413278 336880 413284 336892
rect 413336 336880 413342 336932
rect 444285 336923 444343 336929
rect 444285 336889 444297 336923
rect 444331 336920 444343 336923
rect 444374 336920 444380 336932
rect 444331 336892 444380 336920
rect 444331 336889 444343 336892
rect 444285 336883 444343 336889
rect 444374 336880 444380 336892
rect 444432 336880 444438 336932
rect 459097 336923 459155 336929
rect 459097 336920 459109 336923
rect 447060 336892 459109 336920
rect 99377 336855 99435 336861
rect 99377 336821 99389 336855
rect 99423 336852 99435 336855
rect 108945 336855 109003 336861
rect 108945 336852 108957 336855
rect 99423 336824 108957 336852
rect 99423 336821 99435 336824
rect 99377 336815 99435 336821
rect 108945 336821 108957 336824
rect 108991 336821 109003 336855
rect 108945 336815 109003 336821
rect 118602 336812 118608 336864
rect 118660 336852 118666 336864
rect 278498 336852 278504 336864
rect 118660 336824 278504 336852
rect 118660 336812 118666 336824
rect 278498 336812 278504 336824
rect 278556 336812 278562 336864
rect 327169 336855 327227 336861
rect 327169 336821 327181 336855
rect 327215 336852 327227 336855
rect 343082 336852 343088 336864
rect 327215 336824 343088 336852
rect 327215 336821 327227 336824
rect 327169 336815 327227 336821
rect 343082 336812 343088 336824
rect 343140 336812 343146 336864
rect 344278 336812 344284 336864
rect 344336 336852 344342 336864
rect 350537 336855 350595 336861
rect 350537 336852 350549 336855
rect 344336 336824 350549 336852
rect 344336 336812 344342 336824
rect 350537 336821 350549 336824
rect 350583 336821 350595 336855
rect 350537 336815 350595 336821
rect 351178 336812 351184 336864
rect 351236 336852 351242 336864
rect 351638 336852 351644 336864
rect 351236 336824 351644 336852
rect 351236 336812 351242 336824
rect 351638 336812 351644 336824
rect 351696 336812 351702 336864
rect 354858 336852 354864 336864
rect 352484 336824 354864 336852
rect 113177 336787 113235 336793
rect 113177 336753 113189 336787
rect 113223 336784 113235 336787
rect 122745 336787 122803 336793
rect 122745 336784 122757 336787
rect 113223 336756 122757 336784
rect 113223 336753 113235 336756
rect 113177 336747 113235 336753
rect 122745 336753 122757 336756
rect 122791 336753 122803 336787
rect 122745 336747 122803 336753
rect 125502 336744 125508 336796
rect 125560 336784 125566 336796
rect 281166 336784 281172 336796
rect 125560 336756 281172 336784
rect 125560 336744 125566 336756
rect 281166 336744 281172 336756
rect 281224 336744 281230 336796
rect 290458 336744 290464 336796
rect 290516 336784 290522 336796
rect 344094 336784 344100 336796
rect 290516 336756 344100 336784
rect 290516 336744 290522 336756
rect 344094 336744 344100 336756
rect 344152 336744 344158 336796
rect 344370 336744 344376 336796
rect 344428 336784 344434 336796
rect 352484 336784 352512 336824
rect 354858 336812 354864 336824
rect 354916 336812 354922 336864
rect 362218 336812 362224 336864
rect 362276 336852 362282 336864
rect 365162 336852 365168 336864
rect 362276 336824 365168 336852
rect 362276 336812 362282 336824
rect 365162 336812 365168 336824
rect 365220 336812 365226 336864
rect 381630 336812 381636 336864
rect 381688 336852 381694 336864
rect 384758 336852 384764 336864
rect 381688 336824 384764 336852
rect 381688 336812 381694 336824
rect 384758 336812 384764 336824
rect 384816 336812 384822 336864
rect 396074 336812 396080 336864
rect 396132 336852 396138 336864
rect 398098 336852 398104 336864
rect 396132 336824 398104 336852
rect 396132 336812 396138 336824
rect 398098 336812 398104 336824
rect 398156 336812 398162 336864
rect 423950 336812 423956 336864
rect 424008 336852 424014 336864
rect 427817 336855 427875 336861
rect 427817 336852 427829 336855
rect 424008 336824 427829 336852
rect 424008 336812 424014 336824
rect 427817 336821 427829 336824
rect 427863 336821 427875 336855
rect 427817 336815 427875 336821
rect 428366 336812 428372 336864
rect 428424 336852 428430 336864
rect 431218 336852 431224 336864
rect 428424 336824 431224 336852
rect 428424 336812 428430 336824
rect 431218 336812 431224 336824
rect 431276 336812 431282 336864
rect 431310 336812 431316 336864
rect 431368 336852 431374 336864
rect 433978 336852 433984 336864
rect 431368 336824 433984 336852
rect 431368 336812 431374 336824
rect 433978 336812 433984 336824
rect 434036 336812 434042 336864
rect 434714 336812 434720 336864
rect 434772 336852 434778 336864
rect 435910 336852 435916 336864
rect 434772 336824 435916 336852
rect 434772 336812 434778 336824
rect 435910 336812 435916 336824
rect 435968 336812 435974 336864
rect 440145 336855 440203 336861
rect 440145 336821 440157 336855
rect 440191 336852 440203 336855
rect 446953 336855 447011 336861
rect 446953 336852 446965 336855
rect 440191 336824 446965 336852
rect 440191 336821 440203 336824
rect 440145 336815 440203 336821
rect 446953 336821 446965 336824
rect 446999 336821 447011 336855
rect 446953 336815 447011 336821
rect 344428 336756 352512 336784
rect 344428 336744 344434 336756
rect 352558 336744 352564 336796
rect 352616 336784 352622 336796
rect 357802 336784 357808 336796
rect 352616 336756 357808 336784
rect 352616 336744 352622 336756
rect 357802 336744 357808 336756
rect 357860 336744 357866 336796
rect 363598 336744 363604 336796
rect 363656 336784 363662 336796
rect 364702 336784 364708 336796
rect 363656 336756 364708 336784
rect 363656 336744 363662 336756
rect 364702 336744 364708 336756
rect 364760 336744 364766 336796
rect 370498 336744 370504 336796
rect 370556 336784 370562 336796
rect 372522 336784 372528 336796
rect 370556 336756 372528 336784
rect 370556 336744 370562 336756
rect 372522 336744 372528 336756
rect 372580 336744 372586 336796
rect 376018 336744 376024 336796
rect 376076 336784 376082 336796
rect 376938 336784 376944 336796
rect 376076 336756 376944 336784
rect 376076 336744 376082 336756
rect 376938 336744 376944 336756
rect 376996 336744 377002 336796
rect 377674 336744 377680 336796
rect 377732 336784 377738 336796
rect 378410 336784 378416 336796
rect 377732 336756 378416 336784
rect 377732 336744 377738 336756
rect 378410 336744 378416 336756
rect 378468 336744 378474 336796
rect 392578 336744 392584 336796
rect 392636 336784 392642 336796
rect 393222 336784 393228 336796
rect 392636 336756 393228 336784
rect 392636 336744 392642 336756
rect 393222 336744 393228 336756
rect 393280 336744 393286 336796
rect 394050 336744 394056 336796
rect 394108 336784 394114 336796
rect 394602 336784 394608 336796
rect 394108 336756 394608 336784
rect 394108 336744 394114 336756
rect 394602 336744 394608 336756
rect 394660 336744 394666 336796
rect 395062 336744 395068 336796
rect 395120 336784 395126 336796
rect 395890 336784 395896 336796
rect 395120 336756 395896 336784
rect 395120 336744 395126 336756
rect 395890 336744 395896 336756
rect 395948 336744 395954 336796
rect 396534 336744 396540 336796
rect 396592 336784 396598 336796
rect 398190 336784 398196 336796
rect 396592 336756 398196 336784
rect 396592 336744 396598 336756
rect 398190 336744 398196 336756
rect 398248 336744 398254 336796
rect 429378 336744 429384 336796
rect 429436 336784 429442 336796
rect 430390 336784 430396 336796
rect 429436 336756 430396 336784
rect 429436 336744 429442 336756
rect 430390 336744 430396 336756
rect 430448 336744 430454 336796
rect 430850 336744 430856 336796
rect 430908 336784 430914 336796
rect 431770 336784 431776 336796
rect 430908 336756 431776 336784
rect 430908 336744 430914 336756
rect 431770 336744 431776 336756
rect 431828 336744 431834 336796
rect 432322 336744 432328 336796
rect 432380 336784 432386 336796
rect 433150 336784 433156 336796
rect 432380 336756 433156 336784
rect 432380 336744 432386 336756
rect 433150 336744 433156 336756
rect 433208 336744 433214 336796
rect 433702 336744 433708 336796
rect 433760 336784 433766 336796
rect 434622 336784 434628 336796
rect 433760 336756 434628 336784
rect 433760 336744 433766 336756
rect 434622 336744 434628 336756
rect 434680 336744 434686 336796
rect 435174 336744 435180 336796
rect 435232 336784 435238 336796
rect 436002 336784 436008 336796
rect 435232 336756 436008 336784
rect 435232 336744 435238 336756
rect 436002 336744 436008 336756
rect 436060 336744 436066 336796
rect 436186 336744 436192 336796
rect 436244 336784 436250 336796
rect 437382 336784 437388 336796
rect 436244 336756 437388 336784
rect 436244 336744 436250 336756
rect 437382 336744 437388 336756
rect 437440 336744 437446 336796
rect 444374 336744 444380 336796
rect 444432 336784 444438 336796
rect 447060 336784 447088 336892
rect 459097 336889 459109 336892
rect 459143 336889 459155 336923
rect 459097 336883 459155 336889
rect 459186 336880 459192 336932
rect 459244 336920 459250 336932
rect 460290 336920 460296 336932
rect 459244 336892 460296 336920
rect 459244 336880 459250 336892
rect 460290 336880 460296 336892
rect 460348 336880 460354 336932
rect 461670 336880 461676 336932
rect 461728 336920 461734 336932
rect 464985 336923 465043 336929
rect 464985 336920 464997 336923
rect 461728 336892 464997 336920
rect 461728 336880 461734 336892
rect 464985 336889 464997 336892
rect 465031 336889 465043 336923
rect 464985 336883 465043 336889
rect 465074 336880 465080 336932
rect 465132 336920 465138 336932
rect 466362 336920 466368 336932
rect 465132 336892 466368 336920
rect 465132 336880 465138 336892
rect 466362 336880 466368 336892
rect 466420 336880 466426 336932
rect 466546 336880 466552 336932
rect 466604 336920 466610 336932
rect 470502 336920 470508 336932
rect 466604 336892 470508 336920
rect 466604 336880 466610 336892
rect 470502 336880 470508 336892
rect 470560 336880 470566 336932
rect 454681 336855 454739 336861
rect 454681 336821 454693 336855
rect 454727 336852 454739 336855
rect 459646 336852 459652 336864
rect 454727 336824 459652 336852
rect 454727 336821 454739 336824
rect 454681 336815 454739 336821
rect 459646 336812 459652 336824
rect 459704 336812 459710 336864
rect 460198 336812 460204 336864
rect 460256 336852 460262 336864
rect 460750 336852 460756 336864
rect 460256 336824 460756 336852
rect 460256 336812 460262 336824
rect 460750 336812 460756 336824
rect 460808 336812 460814 336864
rect 461581 336855 461639 336861
rect 461581 336821 461593 336855
rect 461627 336852 461639 336855
rect 469214 336852 469220 336864
rect 461627 336824 469220 336852
rect 461627 336821 461639 336824
rect 461581 336815 461639 336821
rect 469214 336812 469220 336824
rect 469272 336812 469278 336864
rect 509878 336852 509884 336864
rect 469324 336824 509884 336852
rect 444432 336756 447088 336784
rect 444432 336744 444438 336756
rect 457254 336744 457260 336796
rect 457312 336784 457318 336796
rect 457990 336784 457996 336796
rect 457312 336756 457996 336784
rect 457312 336744 457318 336756
rect 457990 336744 457996 336756
rect 458048 336744 458054 336796
rect 458266 336744 458272 336796
rect 458324 336784 458330 336796
rect 459462 336784 459468 336796
rect 458324 336756 459468 336784
rect 458324 336744 458330 336756
rect 459462 336744 459468 336756
rect 459520 336744 459526 336796
rect 459738 336744 459744 336796
rect 459796 336784 459802 336796
rect 460842 336784 460848 336796
rect 459796 336756 460848 336784
rect 459796 336744 459802 336756
rect 460842 336744 460848 336756
rect 460900 336744 460906 336796
rect 461210 336744 461216 336796
rect 461268 336784 461274 336796
rect 462130 336784 462136 336796
rect 461268 336756 462136 336784
rect 461268 336744 461274 336756
rect 462130 336744 462136 336756
rect 462188 336744 462194 336796
rect 462682 336744 462688 336796
rect 462740 336784 462746 336796
rect 463510 336784 463516 336796
rect 462740 336756 463516 336784
rect 462740 336744 462746 336756
rect 463510 336744 463516 336756
rect 463568 336744 463574 336796
rect 464154 336744 464160 336796
rect 464212 336784 464218 336796
rect 464982 336784 464988 336796
rect 464212 336756 464988 336784
rect 464212 336744 464218 336756
rect 464982 336744 464988 336756
rect 465040 336744 465046 336796
rect 469324 336784 469352 336824
rect 509878 336812 509884 336824
rect 509936 336812 509942 336864
rect 505738 336784 505744 336796
rect 465092 336756 469352 336784
rect 469416 336756 505744 336784
rect 323305 336719 323363 336725
rect 323305 336685 323317 336719
rect 323351 336716 323363 336719
rect 323670 336716 323676 336728
rect 323351 336688 323676 336716
rect 323351 336685 323363 336688
rect 323305 336679 323363 336685
rect 323670 336676 323676 336688
rect 323728 336676 323734 336728
rect 464890 336676 464896 336728
rect 464948 336716 464954 336728
rect 465092 336716 465120 336756
rect 464948 336688 465120 336716
rect 465169 336719 465227 336725
rect 464948 336676 464954 336688
rect 465169 336685 465181 336719
rect 465215 336716 465227 336719
rect 469416 336716 469444 336756
rect 505738 336744 505744 336756
rect 505796 336744 505802 336796
rect 465215 336688 469444 336716
rect 465215 336685 465227 336688
rect 465169 336679 465227 336685
rect 437109 336651 437167 336657
rect 437109 336617 437121 336651
rect 437155 336648 437167 336651
rect 444285 336651 444343 336657
rect 444285 336648 444297 336651
rect 437155 336620 444297 336648
rect 437155 336617 437167 336620
rect 437109 336611 437167 336617
rect 444285 336617 444297 336620
rect 444331 336617 444343 336651
rect 444285 336611 444343 336617
rect 236178 335656 236184 335708
rect 236236 335696 236242 335708
rect 237006 335696 237012 335708
rect 236236 335668 237012 335696
rect 236236 335656 236242 335668
rect 237006 335656 237012 335668
rect 237064 335656 237070 335708
rect 302234 335656 302240 335708
rect 302292 335696 302298 335708
rect 302694 335696 302700 335708
rect 302292 335668 302700 335696
rect 302292 335656 302298 335668
rect 302694 335656 302700 335668
rect 302752 335656 302758 335708
rect 331306 335656 331312 335708
rect 331364 335696 331370 335708
rect 331950 335696 331956 335708
rect 331364 335668 331956 335696
rect 331364 335656 331370 335668
rect 331950 335656 331956 335668
rect 332008 335656 332014 335708
rect 334066 335656 334072 335708
rect 334124 335696 334130 335708
rect 334894 335696 334900 335708
rect 334124 335668 334900 335696
rect 334124 335656 334130 335668
rect 334894 335656 334900 335668
rect 334952 335656 334958 335708
rect 236086 335588 236092 335640
rect 236144 335628 236150 335640
rect 236546 335628 236552 335640
rect 236144 335600 236552 335628
rect 236144 335588 236150 335600
rect 236546 335588 236552 335600
rect 236604 335588 236610 335640
rect 241606 335588 241612 335640
rect 241664 335628 241670 335640
rect 242342 335628 242348 335640
rect 241664 335600 242348 335628
rect 241664 335588 241670 335600
rect 242342 335588 242348 335600
rect 242400 335588 242406 335640
rect 260926 335588 260932 335640
rect 260984 335628 260990 335640
rect 261478 335628 261484 335640
rect 260984 335600 261484 335628
rect 260984 335588 260990 335600
rect 261478 335588 261484 335600
rect 261536 335588 261542 335640
rect 262582 335588 262588 335640
rect 262640 335628 262646 335640
rect 263042 335628 263048 335640
rect 262640 335600 263048 335628
rect 262640 335588 262646 335600
rect 263042 335588 263048 335600
rect 263100 335588 263106 335640
rect 263686 335588 263692 335640
rect 263744 335628 263750 335640
rect 264422 335628 264428 335640
rect 263744 335600 264428 335628
rect 263744 335588 263750 335600
rect 264422 335588 264428 335600
rect 264480 335588 264486 335640
rect 265066 335588 265072 335640
rect 265124 335628 265130 335640
rect 265894 335628 265900 335640
rect 265124 335600 265900 335628
rect 265124 335588 265130 335600
rect 265894 335588 265900 335600
rect 265952 335588 265958 335640
rect 266446 335588 266452 335640
rect 266504 335628 266510 335640
rect 267366 335628 267372 335640
rect 266504 335600 267372 335628
rect 266504 335588 266510 335600
rect 267366 335588 267372 335600
rect 267424 335588 267430 335640
rect 280246 335588 280252 335640
rect 280304 335628 280310 335640
rect 280614 335628 280620 335640
rect 280304 335600 280620 335628
rect 280304 335588 280310 335600
rect 280614 335588 280620 335600
rect 280672 335588 280678 335640
rect 283006 335588 283012 335640
rect 283064 335628 283070 335640
rect 283558 335628 283564 335640
rect 283064 335600 283564 335628
rect 283064 335588 283070 335600
rect 283558 335588 283564 335600
rect 283616 335588 283622 335640
rect 285674 335588 285680 335640
rect 285732 335628 285738 335640
rect 285950 335628 285956 335640
rect 285732 335600 285956 335628
rect 285732 335588 285738 335600
rect 285950 335588 285956 335600
rect 286008 335588 286014 335640
rect 287054 335588 287060 335640
rect 287112 335628 287118 335640
rect 287974 335628 287980 335640
rect 287112 335600 287980 335628
rect 287112 335588 287118 335600
rect 287974 335588 287980 335600
rect 288032 335588 288038 335640
rect 288434 335588 288440 335640
rect 288492 335628 288498 335640
rect 289446 335628 289452 335640
rect 288492 335600 289452 335628
rect 288492 335588 288498 335600
rect 289446 335588 289452 335600
rect 289504 335588 289510 335640
rect 292758 335588 292764 335640
rect 292816 335628 292822 335640
rect 293310 335628 293316 335640
rect 292816 335600 293316 335628
rect 292816 335588 292822 335600
rect 293310 335588 293316 335600
rect 293368 335588 293374 335640
rect 298278 335588 298284 335640
rect 298336 335628 298342 335640
rect 298646 335628 298652 335640
rect 298336 335600 298652 335628
rect 298336 335588 298342 335600
rect 298646 335588 298652 335600
rect 298704 335588 298710 335640
rect 300854 335588 300860 335640
rect 300912 335628 300918 335640
rect 301222 335628 301228 335640
rect 300912 335600 301228 335628
rect 300912 335588 300918 335600
rect 301222 335588 301228 335600
rect 301280 335588 301286 335640
rect 303614 335588 303620 335640
rect 303672 335628 303678 335640
rect 304166 335628 304172 335640
rect 303672 335600 304172 335628
rect 303672 335588 303678 335600
rect 304166 335588 304172 335600
rect 304224 335588 304230 335640
rect 304994 335588 305000 335640
rect 305052 335628 305058 335640
rect 305638 335628 305644 335640
rect 305052 335600 305644 335628
rect 305052 335588 305058 335600
rect 305638 335588 305644 335600
rect 305696 335588 305702 335640
rect 307754 335588 307760 335640
rect 307812 335628 307818 335640
rect 308582 335628 308588 335640
rect 307812 335600 308588 335628
rect 307812 335588 307818 335600
rect 308582 335588 308588 335600
rect 308640 335588 308646 335640
rect 309134 335588 309140 335640
rect 309192 335628 309198 335640
rect 310054 335628 310060 335640
rect 309192 335600 310060 335628
rect 309192 335588 309198 335600
rect 310054 335588 310060 335600
rect 310112 335588 310118 335640
rect 310514 335588 310520 335640
rect 310572 335628 310578 335640
rect 311526 335628 311532 335640
rect 310572 335600 311532 335628
rect 310572 335588 310578 335600
rect 311526 335588 311532 335600
rect 311584 335588 311590 335640
rect 321646 335588 321652 335640
rect 321704 335628 321710 335640
rect 322198 335628 322204 335640
rect 321704 335600 322204 335628
rect 321704 335588 321710 335600
rect 322198 335588 322204 335600
rect 322256 335588 322262 335640
rect 329834 335588 329840 335640
rect 329892 335628 329898 335640
rect 330110 335628 330116 335640
rect 329892 335600 330116 335628
rect 329892 335588 329898 335600
rect 330110 335588 330116 335600
rect 330168 335588 330174 335640
rect 331214 335588 331220 335640
rect 331272 335628 331278 335640
rect 331582 335628 331588 335640
rect 331272 335600 331588 335628
rect 331272 335588 331278 335600
rect 331582 335588 331588 335600
rect 331640 335588 331646 335640
rect 332594 335588 332600 335640
rect 332652 335628 332658 335640
rect 333054 335628 333060 335640
rect 332652 335600 333060 335628
rect 332652 335588 332658 335600
rect 333054 335588 333060 335600
rect 333112 335588 333118 335640
rect 333974 335588 333980 335640
rect 334032 335628 334038 335640
rect 334526 335628 334532 335640
rect 334032 335600 334532 335628
rect 334032 335588 334038 335600
rect 334526 335588 334532 335600
rect 334584 335588 334590 335640
rect 338114 335588 338120 335640
rect 338172 335628 338178 335640
rect 338942 335628 338948 335640
rect 338172 335600 338948 335628
rect 338172 335588 338178 335600
rect 338942 335588 338948 335600
rect 339000 335588 339006 335640
rect 356146 335588 356152 335640
rect 356204 335628 356210 335640
rect 356606 335628 356612 335640
rect 356204 335600 356612 335628
rect 356204 335588 356210 335600
rect 356606 335588 356612 335600
rect 356664 335588 356670 335640
rect 358998 335588 359004 335640
rect 359056 335628 359062 335640
rect 359366 335628 359372 335640
rect 359056 335600 359372 335628
rect 359056 335588 359062 335600
rect 359366 335588 359372 335600
rect 359424 335588 359430 335640
rect 250165 335563 250223 335569
rect 250165 335529 250177 335563
rect 250211 335560 250223 335563
rect 250622 335560 250628 335572
rect 250211 335532 250628 335560
rect 250211 335529 250223 335532
rect 250165 335523 250223 335529
rect 250622 335520 250628 335532
rect 250680 335520 250686 335572
rect 248506 335452 248512 335504
rect 248564 335492 248570 335504
rect 249150 335492 249156 335504
rect 248564 335464 249156 335492
rect 248564 335452 248570 335464
rect 249150 335452 249156 335464
rect 249208 335452 249214 335504
rect 285950 335452 285956 335504
rect 286008 335492 286014 335504
rect 286594 335492 286600 335504
rect 286008 335464 286600 335492
rect 286008 335452 286014 335464
rect 286594 335452 286600 335464
rect 286652 335452 286658 335504
rect 278866 335384 278872 335436
rect 278924 335424 278930 335436
rect 278924 335396 279004 335424
rect 278924 335384 278930 335396
rect 278976 335232 279004 335396
rect 580074 335384 580080 335436
rect 580132 335424 580138 335436
rect 580994 335424 581000 335436
rect 580132 335396 581000 335424
rect 580132 335384 580138 335396
rect 580994 335384 581000 335396
rect 581052 335384 581058 335436
rect 367278 335316 367284 335368
rect 367336 335356 367342 335368
rect 367922 335356 367928 335368
rect 367336 335328 367928 335356
rect 367336 335316 367342 335328
rect 367922 335316 367928 335328
rect 367980 335316 367986 335368
rect 580074 335248 580080 335300
rect 580132 335288 580138 335300
rect 580994 335288 581000 335300
rect 580132 335260 581000 335288
rect 580132 335248 580138 335260
rect 580994 335248 581000 335260
rect 581052 335248 581058 335300
rect 278958 335180 278964 335232
rect 279016 335180 279022 335232
rect 332686 335044 332692 335096
rect 332744 335084 332750 335096
rect 333422 335084 333428 335096
rect 332744 335056 333428 335084
rect 332744 335044 332750 335056
rect 333422 335044 333428 335056
rect 333480 335044 333486 335096
rect 302510 334704 302516 334756
rect 302568 334744 302574 334756
rect 303062 334744 303068 334756
rect 302568 334716 303068 334744
rect 302568 334704 302574 334716
rect 303062 334704 303068 334716
rect 303120 334704 303126 334756
rect 258166 334568 258172 334620
rect 258224 334608 258230 334620
rect 258534 334608 258540 334620
rect 258224 334580 258540 334608
rect 258224 334568 258230 334580
rect 258534 334568 258540 334580
rect 258592 334568 258598 334620
rect 270770 334296 270776 334348
rect 270828 334336 270834 334348
rect 271230 334336 271236 334348
rect 270828 334308 271236 334336
rect 270828 334296 270834 334308
rect 271230 334296 271236 334308
rect 271288 334296 271294 334348
rect 272242 334296 272248 334348
rect 272300 334336 272306 334348
rect 272702 334336 272708 334348
rect 272300 334308 272708 334336
rect 272300 334296 272306 334308
rect 272702 334296 272708 334308
rect 272760 334296 272766 334348
rect 335354 333888 335360 333940
rect 335412 333928 335418 333940
rect 335998 333928 336004 333940
rect 335412 333900 336004 333928
rect 335412 333888 335418 333900
rect 335998 333888 336004 333900
rect 336056 333888 336062 333940
rect 278866 333276 278872 333328
rect 278924 333316 278930 333328
rect 279050 333316 279056 333328
rect 278924 333288 279056 333316
rect 278924 333276 278930 333288
rect 279050 333276 279056 333288
rect 279108 333276 279114 333328
rect 306466 333276 306472 333328
rect 306524 333316 306530 333328
rect 306650 333316 306656 333328
rect 306524 333288 306656 333316
rect 306524 333276 306530 333288
rect 306650 333276 306656 333288
rect 306708 333276 306714 333328
rect 242986 332052 242992 332104
rect 243044 332092 243050 332104
rect 243446 332092 243452 332104
rect 243044 332064 243452 332092
rect 243044 332052 243050 332064
rect 243446 332052 243452 332064
rect 243504 332052 243510 332104
rect 331398 331888 331404 331900
rect 331359 331860 331404 331888
rect 331398 331848 331404 331860
rect 331456 331848 331462 331900
rect 336734 331848 336740 331900
rect 336792 331888 336798 331900
rect 336918 331888 336924 331900
rect 336792 331860 336924 331888
rect 336792 331848 336798 331860
rect 336918 331848 336924 331860
rect 336976 331848 336982 331900
rect 328546 331644 328552 331696
rect 328604 331684 328610 331696
rect 329006 331684 329012 331696
rect 328604 331656 329012 331684
rect 328604 331644 328610 331656
rect 329006 331644 329012 331656
rect 329064 331644 329070 331696
rect 341426 331304 341432 331356
rect 341484 331344 341490 331356
rect 341702 331344 341708 331356
rect 341484 331316 341708 331344
rect 341484 331304 341490 331316
rect 341702 331304 341708 331316
rect 341760 331304 341766 331356
rect 299566 331236 299572 331288
rect 299624 331236 299630 331288
rect 259638 331168 259644 331220
rect 259696 331208 259702 331220
rect 259822 331208 259828 331220
rect 259696 331180 259828 331208
rect 259696 331168 259702 331180
rect 259822 331168 259828 331180
rect 259880 331168 259886 331220
rect 262582 331168 262588 331220
rect 262640 331208 262646 331220
rect 262766 331208 262772 331220
rect 262640 331180 262772 331208
rect 262640 331168 262646 331180
rect 262766 331168 262772 331180
rect 262824 331168 262830 331220
rect 299584 331152 299612 331236
rect 303890 331168 303896 331220
rect 303948 331208 303954 331220
rect 304626 331208 304632 331220
rect 303948 331180 304632 331208
rect 303948 331168 303954 331180
rect 304626 331168 304632 331180
rect 304684 331168 304690 331220
rect 389266 331168 389272 331220
rect 389324 331208 389330 331220
rect 389450 331208 389456 331220
rect 389324 331180 389456 331208
rect 389324 331168 389330 331180
rect 389450 331168 389456 331180
rect 389508 331168 389514 331220
rect 459646 331168 459652 331220
rect 459704 331208 459710 331220
rect 460106 331208 460112 331220
rect 459704 331180 460112 331208
rect 459704 331168 459710 331180
rect 460106 331168 460112 331180
rect 460164 331168 460170 331220
rect 299566 331100 299572 331152
rect 299624 331100 299630 331152
rect 299750 331100 299756 331152
rect 299808 331140 299814 331152
rect 300302 331140 300308 331152
rect 299808 331112 300308 331140
rect 299808 331100 299814 331112
rect 300302 331100 300308 331112
rect 300360 331100 300366 331152
rect 299474 331032 299480 331084
rect 299532 331072 299538 331084
rect 299658 331072 299664 331084
rect 299532 331044 299664 331072
rect 299532 331032 299538 331044
rect 299658 331032 299664 331044
rect 299716 331032 299722 331084
rect 301130 328448 301136 328500
rect 301188 328488 301194 328500
rect 301682 328488 301688 328500
rect 301188 328460 301688 328488
rect 301188 328448 301194 328460
rect 301682 328448 301688 328460
rect 301740 328448 301746 328500
rect 339770 328448 339776 328500
rect 339828 328488 339834 328500
rect 340322 328488 340328 328500
rect 339828 328460 340328 328488
rect 339828 328448 339834 328460
rect 340322 328448 340328 328460
rect 340380 328448 340386 328500
rect 366913 328491 366971 328497
rect 366913 328457 366925 328491
rect 366959 328488 366971 328491
rect 367002 328488 367008 328500
rect 366959 328460 367008 328488
rect 366959 328457 366971 328460
rect 366913 328451 366971 328457
rect 367002 328448 367008 328460
rect 367060 328448 367066 328500
rect 372706 328448 372712 328500
rect 372764 328488 372770 328500
rect 373074 328488 373080 328500
rect 372764 328460 373080 328488
rect 372764 328448 372770 328460
rect 373074 328448 373080 328460
rect 373132 328448 373138 328500
rect 259822 328420 259828 328432
rect 259783 328392 259828 328420
rect 259822 328380 259828 328392
rect 259880 328380 259886 328432
rect 265250 328380 265256 328432
rect 265308 328420 265314 328432
rect 265342 328420 265348 328432
rect 265308 328392 265348 328420
rect 265308 328380 265314 328392
rect 265342 328380 265348 328392
rect 265400 328380 265406 328432
rect 294230 328380 294236 328432
rect 294288 328420 294294 328432
rect 294414 328420 294420 328432
rect 294288 328392 294420 328420
rect 294288 328380 294294 328392
rect 294414 328380 294420 328392
rect 294472 328380 294478 328432
rect 295518 328380 295524 328432
rect 295576 328420 295582 328432
rect 295702 328420 295708 328432
rect 295576 328392 295708 328420
rect 295576 328380 295582 328392
rect 295702 328380 295708 328392
rect 295760 328380 295766 328432
rect 296806 328380 296812 328432
rect 296864 328420 296870 328432
rect 296990 328420 296996 328432
rect 296864 328392 296996 328420
rect 296864 328380 296870 328392
rect 296990 328380 296996 328392
rect 297048 328380 297054 328432
rect 341334 328420 341340 328432
rect 341295 328392 341340 328420
rect 341334 328380 341340 328392
rect 341392 328380 341398 328432
rect 389450 328420 389456 328432
rect 389411 328392 389456 328420
rect 389450 328380 389456 328392
rect 389508 328380 389514 328432
rect 393590 328380 393596 328432
rect 393648 328420 393654 328432
rect 393682 328420 393688 328432
rect 393648 328392 393688 328420
rect 393648 328380 393654 328392
rect 393682 328380 393688 328392
rect 393740 328380 393746 328432
rect 367002 328352 367008 328364
rect 366963 328324 367008 328352
rect 367002 328312 367008 328324
rect 367060 328312 367066 328364
rect 337010 327196 337016 327208
rect 336844 327168 337016 327196
rect 336844 327140 336872 327168
rect 337010 327156 337016 327168
rect 337068 327156 337074 327208
rect 250162 327128 250168 327140
rect 250123 327100 250168 327128
rect 250162 327088 250168 327100
rect 250220 327088 250226 327140
rect 323302 327128 323308 327140
rect 323263 327100 323308 327128
rect 323302 327088 323308 327100
rect 323360 327088 323366 327140
rect 324682 327088 324688 327140
rect 324740 327128 324746 327140
rect 325050 327128 325056 327140
rect 324740 327100 325056 327128
rect 324740 327088 324746 327100
rect 325050 327088 325056 327100
rect 325108 327088 325114 327140
rect 325970 327088 325976 327140
rect 326028 327128 326034 327140
rect 326614 327128 326620 327140
rect 326028 327100 326620 327128
rect 326028 327088 326034 327100
rect 326614 327088 326620 327100
rect 326672 327088 326678 327140
rect 336826 327088 336832 327140
rect 336884 327088 336890 327140
rect 265253 327063 265311 327069
rect 265253 327029 265265 327063
rect 265299 327060 265311 327063
rect 265342 327060 265348 327072
rect 265299 327032 265348 327060
rect 265299 327029 265311 327032
rect 265253 327023 265311 327029
rect 265342 327020 265348 327032
rect 265400 327020 265406 327072
rect 301041 327063 301099 327069
rect 301041 327029 301053 327063
rect 301087 327060 301099 327063
rect 301130 327060 301136 327072
rect 301087 327032 301136 327060
rect 301087 327029 301099 327032
rect 301041 327023 301099 327029
rect 301130 327020 301136 327032
rect 301188 327020 301194 327072
rect 327258 327060 327264 327072
rect 327219 327032 327264 327060
rect 327258 327020 327264 327032
rect 327316 327020 327322 327072
rect 288710 325660 288716 325712
rect 288768 325700 288774 325712
rect 288802 325700 288808 325712
rect 288768 325672 288808 325700
rect 288768 325660 288774 325672
rect 288802 325660 288808 325672
rect 288860 325660 288866 325712
rect 580074 325660 580080 325712
rect 580132 325700 580138 325712
rect 580902 325700 580908 325712
rect 580132 325672 580908 325700
rect 580132 325660 580138 325672
rect 580902 325660 580908 325672
rect 580960 325660 580966 325712
rect 3326 324232 3332 324284
rect 3384 324272 3390 324284
rect 14458 324272 14464 324284
rect 3384 324244 14464 324272
rect 3384 324232 3390 324244
rect 14458 324232 14464 324244
rect 14516 324232 14522 324284
rect 469950 322872 469956 322924
rect 470008 322912 470014 322924
rect 580074 322912 580080 322924
rect 470008 322884 580080 322912
rect 470008 322872 470014 322884
rect 580074 322872 580080 322884
rect 580132 322872 580138 322924
rect 273530 321756 273536 321768
rect 273491 321728 273536 321756
rect 273530 321716 273536 321728
rect 273588 321716 273594 321768
rect 262766 321580 262772 321632
rect 262824 321580 262830 321632
rect 266633 321623 266691 321629
rect 266633 321589 266645 321623
rect 266679 321620 266691 321623
rect 266722 321620 266728 321632
rect 266679 321592 266728 321620
rect 266679 321589 266691 321592
rect 266633 321583 266691 321589
rect 266722 321580 266728 321592
rect 266780 321580 266786 321632
rect 267737 321623 267795 321629
rect 267737 321589 267749 321623
rect 267783 321620 267795 321623
rect 267826 321620 267832 321632
rect 267783 321592 267832 321620
rect 267783 321589 267795 321592
rect 267737 321583 267795 321589
rect 267826 321580 267832 321592
rect 267884 321580 267890 321632
rect 281721 321623 281779 321629
rect 281721 321589 281733 321623
rect 281767 321620 281779 321623
rect 281810 321620 281816 321632
rect 281767 321592 281816 321620
rect 281767 321589 281779 321592
rect 281721 321583 281779 321589
rect 281810 321580 281816 321592
rect 281868 321580 281874 321632
rect 310790 321580 310796 321632
rect 310848 321580 310854 321632
rect 375834 321580 375840 321632
rect 375892 321580 375898 321632
rect 377122 321580 377128 321632
rect 377180 321580 377186 321632
rect 230750 321512 230756 321564
rect 230808 321552 230814 321564
rect 230934 321552 230940 321564
rect 230808 321524 230940 321552
rect 230808 321512 230814 321524
rect 230934 321512 230940 321524
rect 230992 321512 230998 321564
rect 232222 321512 232228 321564
rect 232280 321552 232286 321564
rect 232406 321552 232412 321564
rect 232280 321524 232412 321552
rect 232280 321512 232286 321524
rect 232406 321512 232412 321524
rect 232464 321512 232470 321564
rect 262784 321484 262812 321580
rect 262858 321484 262864 321496
rect 262784 321456 262864 321484
rect 262858 321444 262864 321456
rect 262916 321444 262922 321496
rect 310808 321484 310836 321580
rect 310882 321484 310888 321496
rect 310808 321456 310888 321484
rect 310882 321444 310888 321456
rect 310940 321444 310946 321496
rect 375852 321416 375880 321580
rect 375926 321416 375932 321428
rect 375852 321388 375932 321416
rect 375926 321376 375932 321388
rect 375984 321376 375990 321428
rect 377140 321416 377168 321580
rect 377214 321416 377220 321428
rect 377140 321388 377220 321416
rect 377214 321376 377220 321388
rect 377272 321376 377278 321428
rect 331398 318900 331404 318912
rect 331359 318872 331404 318900
rect 331398 318860 331404 318872
rect 331456 318860 331462 318912
rect 259825 318835 259883 318841
rect 259825 318801 259837 318835
rect 259871 318832 259883 318835
rect 259914 318832 259920 318844
rect 259871 318804 259920 318832
rect 259871 318801 259883 318804
rect 259825 318795 259883 318801
rect 259914 318792 259920 318804
rect 259972 318792 259978 318844
rect 266630 318832 266636 318844
rect 266591 318804 266636 318832
rect 266630 318792 266636 318804
rect 266688 318792 266694 318844
rect 267734 318832 267740 318844
rect 267695 318804 267740 318832
rect 267734 318792 267740 318804
rect 267792 318792 267798 318844
rect 299750 318792 299756 318844
rect 299808 318832 299814 318844
rect 299842 318832 299848 318844
rect 299808 318804 299848 318832
rect 299808 318792 299814 318804
rect 299842 318792 299848 318804
rect 299900 318792 299906 318844
rect 302510 318792 302516 318844
rect 302568 318832 302574 318844
rect 302602 318832 302608 318844
rect 302568 318804 302608 318832
rect 302568 318792 302574 318804
rect 302602 318792 302608 318804
rect 302660 318792 302666 318844
rect 306742 318792 306748 318844
rect 306800 318832 306806 318844
rect 306834 318832 306840 318844
rect 306800 318804 306840 318832
rect 306800 318792 306806 318804
rect 306834 318792 306840 318804
rect 306892 318792 306898 318844
rect 341337 318835 341395 318841
rect 341337 318801 341349 318835
rect 341383 318832 341395 318835
rect 341426 318832 341432 318844
rect 341383 318804 341432 318832
rect 341383 318801 341395 318804
rect 341337 318795 341395 318801
rect 341426 318792 341432 318804
rect 341484 318792 341490 318844
rect 357618 318792 357624 318844
rect 357676 318832 357682 318844
rect 357710 318832 357716 318844
rect 357676 318804 357716 318832
rect 357676 318792 357682 318804
rect 357710 318792 357716 318804
rect 357768 318792 357774 318844
rect 367002 318832 367008 318844
rect 366963 318804 367008 318832
rect 367002 318792 367008 318804
rect 367060 318792 367066 318844
rect 389453 318835 389511 318841
rect 389453 318801 389465 318835
rect 389499 318832 389511 318835
rect 389542 318832 389548 318844
rect 389499 318804 389548 318832
rect 389499 318801 389511 318804
rect 389453 318795 389511 318801
rect 389542 318792 389548 318804
rect 389600 318792 389606 318844
rect 431402 318792 431408 318844
rect 431460 318832 431466 318844
rect 431494 318832 431500 318844
rect 431460 318804 431500 318832
rect 431460 318792 431466 318804
rect 431494 318792 431500 318804
rect 431552 318792 431558 318844
rect 230845 318767 230903 318773
rect 230845 318733 230857 318767
rect 230891 318764 230903 318767
rect 230934 318764 230940 318776
rect 230891 318736 230940 318764
rect 230891 318733 230903 318736
rect 230845 318727 230903 318733
rect 230934 318724 230940 318736
rect 230992 318724 230998 318776
rect 235074 318764 235080 318776
rect 235035 318736 235080 318764
rect 235074 318724 235080 318736
rect 235132 318724 235138 318776
rect 236270 318764 236276 318776
rect 236231 318736 236276 318764
rect 236270 318724 236276 318736
rect 236328 318724 236334 318776
rect 372706 318764 372712 318776
rect 372667 318736 372712 318764
rect 372706 318724 372712 318736
rect 372764 318724 372770 318776
rect 273530 317540 273536 317552
rect 273491 317512 273536 317540
rect 273530 317500 273536 317512
rect 273588 317500 273594 317552
rect 265250 317472 265256 317484
rect 265211 317444 265256 317472
rect 265250 317432 265256 317444
rect 265308 317432 265314 317484
rect 301038 317472 301044 317484
rect 300999 317444 301044 317472
rect 301038 317432 301044 317444
rect 301096 317432 301102 317484
rect 327258 317472 327264 317484
rect 327219 317444 327264 317472
rect 327258 317432 327264 317444
rect 327316 317432 327322 317484
rect 250162 317404 250168 317416
rect 250123 317376 250168 317404
rect 250162 317364 250168 317376
rect 250220 317364 250226 317416
rect 251542 317404 251548 317416
rect 251503 317376 251548 317404
rect 251542 317364 251548 317376
rect 251600 317364 251606 317416
rect 270770 317404 270776 317416
rect 270731 317376 270776 317404
rect 270770 317364 270776 317376
rect 270828 317364 270834 317416
rect 272242 317404 272248 317416
rect 272203 317376 272248 317404
rect 272242 317364 272248 317376
rect 272300 317364 272306 317416
rect 273530 317364 273536 317416
rect 273588 317404 273594 317416
rect 273588 317376 273668 317404
rect 273588 317364 273594 317376
rect 273640 317348 273668 317376
rect 290090 317364 290096 317416
rect 290148 317404 290154 317416
rect 290182 317404 290188 317416
rect 290148 317376 290188 317404
rect 290148 317364 290154 317376
rect 290182 317364 290188 317376
rect 290240 317364 290246 317416
rect 291562 317364 291568 317416
rect 291620 317404 291626 317416
rect 291654 317404 291660 317416
rect 291620 317376 291660 317404
rect 291620 317364 291626 317376
rect 291654 317364 291660 317376
rect 291712 317364 291718 317416
rect 296898 317364 296904 317416
rect 296956 317404 296962 317416
rect 296990 317404 296996 317416
rect 296956 317376 296996 317404
rect 296956 317364 296962 317376
rect 296990 317364 296996 317376
rect 297048 317364 297054 317416
rect 306834 317404 306840 317416
rect 306795 317376 306840 317404
rect 306834 317364 306840 317376
rect 306892 317364 306898 317416
rect 330202 317404 330208 317416
rect 330163 317376 330208 317404
rect 330202 317364 330208 317376
rect 330260 317364 330266 317416
rect 331398 317404 331404 317416
rect 331359 317376 331404 317404
rect 331398 317364 331404 317376
rect 331456 317364 331462 317416
rect 393590 317404 393596 317416
rect 393551 317376 393596 317404
rect 393590 317364 393596 317376
rect 393648 317364 393654 317416
rect 460198 317404 460204 317416
rect 460159 317376 460204 317404
rect 460198 317364 460204 317376
rect 460256 317364 460262 317416
rect 273622 317296 273628 317348
rect 273680 317296 273686 317348
rect 579982 316072 579988 316124
rect 580040 316112 580046 316124
rect 580994 316112 581000 316124
rect 580040 316084 581000 316112
rect 580040 316072 580046 316084
rect 580994 316072 581000 316084
rect 581052 316072 581058 316124
rect 281718 316044 281724 316056
rect 281679 316016 281724 316044
rect 281718 316004 281724 316016
rect 281776 316004 281782 316056
rect 285766 316004 285772 316056
rect 285824 316044 285830 316056
rect 286042 316044 286048 316056
rect 285824 316016 286048 316044
rect 285824 316004 285830 316016
rect 286042 316004 286048 316016
rect 286100 316004 286106 316056
rect 267734 315936 267740 315988
rect 267792 315976 267798 315988
rect 267792 315948 267837 315976
rect 267792 315936 267798 315948
rect 580074 315936 580080 315988
rect 580132 315976 580138 315988
rect 580994 315976 581000 315988
rect 580132 315948 581000 315976
rect 580132 315936 580138 315948
rect 580994 315936 581000 315948
rect 581052 315936 581058 315988
rect 250162 312576 250168 312588
rect 250123 312548 250168 312576
rect 250162 312536 250168 312548
rect 250220 312536 250226 312588
rect 232406 311964 232412 311976
rect 232332 311936 232412 311964
rect 232332 311840 232360 311936
rect 232406 311924 232412 311936
rect 232464 311924 232470 311976
rect 244366 311924 244372 311976
rect 244424 311924 244430 311976
rect 245838 311924 245844 311976
rect 245896 311924 245902 311976
rect 284754 311924 284760 311976
rect 284812 311924 284818 311976
rect 299842 311964 299848 311976
rect 299768 311936 299848 311964
rect 232314 311788 232320 311840
rect 232372 311788 232378 311840
rect 235074 311828 235080 311840
rect 235035 311800 235080 311828
rect 235074 311788 235080 311800
rect 235132 311788 235138 311840
rect 244384 311760 244412 311924
rect 244458 311760 244464 311772
rect 244384 311732 244464 311760
rect 244458 311720 244464 311732
rect 244516 311720 244522 311772
rect 245856 311760 245884 311924
rect 259730 311856 259736 311908
rect 259788 311896 259794 311908
rect 259914 311896 259920 311908
rect 259788 311868 259920 311896
rect 259788 311856 259794 311868
rect 259914 311856 259920 311868
rect 259972 311856 259978 311908
rect 284772 311840 284800 311924
rect 299768 311840 299796 311936
rect 299842 311924 299848 311936
rect 299900 311924 299906 311976
rect 302602 311964 302608 311976
rect 302528 311936 302608 311964
rect 302528 311840 302556 311936
rect 302602 311924 302608 311936
rect 302660 311924 302666 311976
rect 310882 311964 310888 311976
rect 310843 311936 310888 311964
rect 310882 311924 310888 311936
rect 310940 311924 310946 311976
rect 323302 311964 323308 311976
rect 323228 311936 323308 311964
rect 323228 311908 323256 311936
rect 323302 311924 323308 311936
rect 323360 311924 323366 311976
rect 337102 311964 337108 311976
rect 337063 311936 337108 311964
rect 337102 311924 337108 311936
rect 337160 311924 337166 311976
rect 431402 311924 431408 311976
rect 431460 311964 431466 311976
rect 431494 311964 431500 311976
rect 431460 311936 431500 311964
rect 431460 311924 431466 311936
rect 431494 311924 431500 311936
rect 431552 311924 431558 311976
rect 323210 311856 323216 311908
rect 323268 311856 323274 311908
rect 341242 311856 341248 311908
rect 341300 311896 341306 311908
rect 341426 311896 341432 311908
rect 341300 311868 341432 311896
rect 341300 311856 341306 311868
rect 341426 311856 341432 311868
rect 341484 311856 341490 311908
rect 389358 311856 389364 311908
rect 389416 311896 389422 311908
rect 389542 311896 389548 311908
rect 389416 311868 389548 311896
rect 389416 311856 389422 311868
rect 389542 311856 389548 311868
rect 389600 311856 389606 311908
rect 284754 311788 284760 311840
rect 284812 311788 284818 311840
rect 299750 311788 299756 311840
rect 299808 311788 299814 311840
rect 302510 311788 302516 311840
rect 302568 311788 302574 311840
rect 245930 311760 245936 311772
rect 245856 311732 245936 311760
rect 245930 311720 245936 311732
rect 245988 311720 245994 311772
rect 239122 311652 239128 311704
rect 239180 311652 239186 311704
rect 239140 311568 239168 311652
rect 239122 311516 239128 311568
rect 239180 311516 239186 311568
rect 267737 311151 267795 311157
rect 267737 311117 267749 311151
rect 267783 311148 267795 311151
rect 267826 311148 267832 311160
rect 267783 311120 267832 311148
rect 267783 311117 267795 311120
rect 267737 311111 267795 311117
rect 267826 311108 267832 311120
rect 267884 311108 267890 311160
rect 266630 309244 266636 309256
rect 266591 309216 266636 309244
rect 266630 309204 266636 309216
rect 266688 309204 266694 309256
rect 230842 309176 230848 309188
rect 230803 309148 230848 309176
rect 230842 309136 230848 309148
rect 230900 309136 230906 309188
rect 236270 309176 236276 309188
rect 236231 309148 236276 309176
rect 236270 309136 236276 309148
rect 236328 309136 236334 309188
rect 327166 309136 327172 309188
rect 327224 309136 327230 309188
rect 372706 309176 372712 309188
rect 372667 309148 372712 309176
rect 372706 309136 372712 309148
rect 372764 309136 372770 309188
rect 265250 309108 265256 309120
rect 265211 309080 265256 309108
rect 265250 309068 265256 309080
rect 265308 309068 265314 309120
rect 327184 309052 327212 309136
rect 337105 309111 337163 309117
rect 337105 309077 337117 309111
rect 337151 309108 337163 309111
rect 337194 309108 337200 309120
rect 337151 309080 337200 309108
rect 337151 309077 337163 309080
rect 337105 309071 337163 309077
rect 337194 309068 337200 309080
rect 337252 309068 337258 309120
rect 341153 309111 341211 309117
rect 341153 309077 341165 309111
rect 341199 309108 341211 309111
rect 341242 309108 341248 309120
rect 341199 309080 341248 309108
rect 341199 309077 341211 309080
rect 341153 309071 341211 309077
rect 341242 309068 341248 309080
rect 341300 309068 341306 309120
rect 367002 309108 367008 309120
rect 366963 309080 367008 309108
rect 367002 309068 367008 309080
rect 367060 309068 367066 309120
rect 327166 309000 327172 309052
rect 327224 309000 327230 309052
rect 310698 307844 310704 307896
rect 310756 307884 310762 307896
rect 310885 307887 310943 307893
rect 310885 307884 310897 307887
rect 310756 307856 310897 307884
rect 310756 307844 310762 307856
rect 310885 307853 310897 307856
rect 310931 307853 310943 307887
rect 310885 307847 310943 307853
rect 251542 307816 251548 307828
rect 251503 307788 251548 307816
rect 251542 307776 251548 307788
rect 251600 307776 251606 307828
rect 270770 307816 270776 307828
rect 270731 307788 270776 307816
rect 270770 307776 270776 307788
rect 270828 307776 270834 307828
rect 272242 307816 272248 307828
rect 272203 307788 272248 307816
rect 272242 307776 272248 307788
rect 272300 307776 272306 307828
rect 330202 307816 330208 307828
rect 330163 307788 330208 307816
rect 330202 307776 330208 307788
rect 330260 307776 330266 307828
rect 393590 307816 393596 307828
rect 393551 307788 393596 307816
rect 393590 307776 393596 307788
rect 393648 307776 393654 307828
rect 460198 307816 460204 307828
rect 460159 307788 460204 307816
rect 460198 307776 460204 307788
rect 460256 307776 460262 307828
rect 288713 307751 288771 307757
rect 288713 307717 288725 307751
rect 288759 307748 288771 307751
rect 288802 307748 288808 307760
rect 288759 307720 288808 307748
rect 288759 307717 288771 307720
rect 288713 307711 288771 307717
rect 288802 307708 288808 307720
rect 288860 307708 288866 307760
rect 310698 307748 310704 307760
rect 310659 307720 310704 307748
rect 310698 307708 310704 307720
rect 310756 307708 310762 307760
rect 337102 307748 337108 307760
rect 337063 307720 337108 307748
rect 337102 307708 337108 307720
rect 337160 307708 337166 307760
rect 286134 306348 286140 306400
rect 286192 306388 286198 306400
rect 286226 306388 286232 306400
rect 286192 306360 286232 306388
rect 286192 306348 286198 306360
rect 286226 306348 286232 306360
rect 286284 306348 286290 306400
rect 288710 306388 288716 306400
rect 288671 306360 288716 306388
rect 288710 306348 288716 306360
rect 288768 306348 288774 306400
rect 317506 306348 317512 306400
rect 317564 306388 317570 306400
rect 317690 306388 317696 306400
rect 317564 306360 317696 306388
rect 317564 306348 317570 306360
rect 317690 306348 317696 306360
rect 317748 306348 317754 306400
rect 463694 306348 463700 306400
rect 463752 306388 463758 306400
rect 463878 306388 463884 306400
rect 463752 306360 463884 306388
rect 463752 306348 463758 306360
rect 463878 306348 463884 306360
rect 463936 306348 463942 306400
rect 580074 306348 580080 306400
rect 580132 306388 580138 306400
rect 580902 306388 580908 306400
rect 580132 306360 580908 306388
rect 580132 306348 580138 306360
rect 580902 306348 580908 306360
rect 580960 306348 580966 306400
rect 266630 305028 266636 305040
rect 266591 305000 266636 305028
rect 266630 304988 266636 305000
rect 266688 304988 266694 305040
rect 291746 304920 291752 304972
rect 291804 304960 291810 304972
rect 291838 304960 291844 304972
rect 291804 304932 291844 304960
rect 291804 304920 291810 304932
rect 291838 304920 291844 304932
rect 291896 304920 291902 304972
rect 294230 304240 294236 304292
rect 294288 304280 294294 304292
rect 294414 304280 294420 304292
rect 294288 304252 294420 304280
rect 294288 304240 294294 304252
rect 294414 304240 294420 304252
rect 294472 304240 294478 304292
rect 295518 304240 295524 304292
rect 295576 304280 295582 304292
rect 295702 304280 295708 304292
rect 295576 304252 295708 304280
rect 295576 304240 295582 304252
rect 295702 304240 295708 304252
rect 295760 304240 295766 304292
rect 323210 304280 323216 304292
rect 323171 304252 323216 304280
rect 323210 304240 323216 304252
rect 323268 304240 323274 304292
rect 291565 303603 291623 303609
rect 291565 303569 291577 303603
rect 291611 303600 291623 303603
rect 291746 303600 291752 303612
rect 291611 303572 291752 303600
rect 291611 303569 291623 303572
rect 291565 303563 291623 303569
rect 291746 303560 291752 303572
rect 291804 303560 291810 303612
rect 259641 302311 259699 302317
rect 259641 302277 259653 302311
rect 259687 302308 259699 302311
rect 259730 302308 259736 302320
rect 259687 302280 259736 302308
rect 259687 302277 259699 302280
rect 259641 302271 259699 302277
rect 259730 302268 259736 302280
rect 259788 302268 259794 302320
rect 357526 302200 357532 302252
rect 357584 302240 357590 302252
rect 357710 302240 357716 302252
rect 357584 302212 357716 302240
rect 357584 302200 357590 302212
rect 357710 302200 357716 302212
rect 357768 302200 357774 302252
rect 389174 302200 389180 302252
rect 389232 302240 389238 302252
rect 389358 302240 389364 302252
rect 389232 302212 389364 302240
rect 389232 302200 389238 302212
rect 389358 302200 389364 302212
rect 389416 302200 389422 302252
rect 431310 302200 431316 302252
rect 431368 302240 431374 302252
rect 431494 302240 431500 302252
rect 431368 302212 431500 302240
rect 431368 302200 431374 302212
rect 431494 302200 431500 302212
rect 431552 302200 431558 302252
rect 296806 301112 296812 301164
rect 296864 301152 296870 301164
rect 296990 301152 296996 301164
rect 296864 301124 296996 301152
rect 296864 301112 296870 301124
rect 296990 301112 296996 301124
rect 297048 301112 297054 301164
rect 265253 300135 265311 300141
rect 265253 300101 265265 300135
rect 265299 300132 265311 300135
rect 265342 300132 265348 300144
rect 265299 300104 265348 300132
rect 265299 300101 265311 300104
rect 265253 300095 265311 300101
rect 265342 300092 265348 300104
rect 265400 300092 265406 300144
rect 262585 299659 262643 299665
rect 262585 299625 262597 299659
rect 262631 299656 262643 299659
rect 262674 299656 262680 299668
rect 262631 299628 262680 299656
rect 262631 299625 262643 299628
rect 262585 299619 262643 299625
rect 262674 299616 262680 299628
rect 262732 299616 262738 299668
rect 331398 299588 331404 299600
rect 331359 299560 331404 299588
rect 331398 299548 331404 299560
rect 331456 299548 331462 299600
rect 266630 299480 266636 299532
rect 266688 299520 266694 299532
rect 266722 299520 266728 299532
rect 266688 299492 266728 299520
rect 266688 299480 266694 299492
rect 266722 299480 266728 299492
rect 266780 299480 266786 299532
rect 299750 299480 299756 299532
rect 299808 299520 299814 299532
rect 299842 299520 299848 299532
rect 299808 299492 299848 299520
rect 299808 299480 299814 299492
rect 299842 299480 299848 299492
rect 299900 299480 299906 299532
rect 302510 299480 302516 299532
rect 302568 299520 302574 299532
rect 302602 299520 302608 299532
rect 302568 299492 302608 299520
rect 302568 299480 302574 299492
rect 302602 299480 302608 299492
rect 302660 299480 302666 299532
rect 306834 299520 306840 299532
rect 306795 299492 306840 299520
rect 306834 299480 306840 299492
rect 306892 299480 306898 299532
rect 323213 299523 323271 299529
rect 323213 299489 323225 299523
rect 323259 299520 323271 299523
rect 323302 299520 323308 299532
rect 323259 299492 323308 299520
rect 323259 299489 323271 299492
rect 323213 299483 323271 299489
rect 323302 299480 323308 299492
rect 323360 299480 323366 299532
rect 341150 299520 341156 299532
rect 341111 299492 341156 299520
rect 341150 299480 341156 299492
rect 341208 299480 341214 299532
rect 367002 299520 367008 299532
rect 366963 299492 367008 299520
rect 367002 299480 367008 299492
rect 367060 299480 367066 299532
rect 235074 299452 235080 299464
rect 235035 299424 235080 299452
rect 235074 299412 235080 299424
rect 235132 299412 235138 299464
rect 236270 299452 236276 299464
rect 236231 299424 236276 299452
rect 236270 299412 236276 299424
rect 236328 299412 236334 299464
rect 270770 299452 270776 299464
rect 270731 299424 270776 299452
rect 270770 299412 270776 299424
rect 270828 299412 270834 299464
rect 272242 299452 272248 299464
rect 272203 299424 272248 299452
rect 272242 299412 272248 299424
rect 272300 299412 272306 299464
rect 273530 299412 273536 299464
rect 273588 299412 273594 299464
rect 281718 299412 281724 299464
rect 281776 299452 281782 299464
rect 281810 299452 281816 299464
rect 281776 299424 281816 299452
rect 281776 299412 281782 299424
rect 281810 299412 281816 299424
rect 281868 299412 281874 299464
rect 284662 299412 284668 299464
rect 284720 299452 284726 299464
rect 284754 299452 284760 299464
rect 284720 299424 284760 299452
rect 284720 299412 284726 299424
rect 284754 299412 284760 299424
rect 284812 299412 284818 299464
rect 324682 299452 324688 299464
rect 324643 299424 324688 299452
rect 324682 299412 324688 299424
rect 324740 299412 324746 299464
rect 325878 299412 325884 299464
rect 325936 299412 325942 299464
rect 372706 299452 372712 299464
rect 372667 299424 372712 299452
rect 372706 299412 372712 299424
rect 372764 299412 372770 299464
rect 469858 299412 469864 299464
rect 469916 299452 469922 299464
rect 580166 299452 580172 299464
rect 469916 299424 580172 299452
rect 469916 299412 469922 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 273548 299328 273576 299412
rect 325896 299384 325924 299412
rect 325970 299384 325976 299396
rect 325896 299356 325976 299384
rect 325970 299344 325976 299356
rect 326028 299344 326034 299396
rect 273530 299276 273536 299328
rect 273588 299276 273594 299328
rect 286042 298188 286048 298240
rect 286100 298228 286106 298240
rect 286134 298228 286140 298240
rect 286100 298200 286140 298228
rect 286100 298188 286106 298200
rect 286134 298188 286140 298200
rect 286192 298188 286198 298240
rect 247034 298120 247040 298172
rect 247092 298160 247098 298172
rect 247310 298160 247316 298172
rect 247092 298132 247316 298160
rect 247092 298120 247098 298132
rect 247310 298120 247316 298132
rect 247368 298120 247374 298172
rect 288894 298120 288900 298172
rect 288952 298120 288958 298172
rect 310701 298163 310759 298169
rect 310701 298129 310713 298163
rect 310747 298160 310759 298163
rect 310882 298160 310888 298172
rect 310747 298132 310888 298160
rect 310747 298129 310759 298132
rect 310701 298123 310759 298129
rect 310882 298120 310888 298132
rect 310940 298120 310946 298172
rect 337105 298163 337163 298169
rect 337105 298129 337117 298163
rect 337151 298160 337163 298163
rect 337286 298160 337292 298172
rect 337151 298132 337292 298160
rect 337151 298129 337163 298132
rect 337105 298123 337163 298129
rect 337286 298120 337292 298132
rect 337344 298120 337350 298172
rect 251361 298095 251419 298101
rect 251361 298061 251373 298095
rect 251407 298092 251419 298095
rect 251542 298092 251548 298104
rect 251407 298064 251548 298092
rect 251407 298061 251419 298064
rect 251361 298055 251419 298061
rect 251542 298052 251548 298064
rect 251600 298052 251606 298104
rect 266722 298092 266728 298104
rect 266683 298064 266728 298092
rect 266722 298052 266728 298064
rect 266780 298052 266786 298104
rect 281718 298052 281724 298104
rect 281776 298092 281782 298104
rect 281810 298092 281816 298104
rect 281776 298064 281816 298092
rect 281776 298052 281782 298064
rect 281810 298052 281816 298064
rect 281868 298052 281874 298104
rect 284662 298052 284668 298104
rect 284720 298092 284726 298104
rect 284754 298092 284760 298104
rect 284720 298064 284760 298092
rect 284720 298052 284726 298064
rect 284754 298052 284760 298064
rect 284812 298052 284818 298104
rect 286042 298052 286048 298104
rect 286100 298092 286106 298104
rect 286134 298092 286140 298104
rect 286100 298064 286140 298092
rect 286100 298052 286106 298064
rect 286134 298052 286140 298064
rect 286192 298052 286198 298104
rect 288912 298036 288940 298120
rect 301038 298092 301044 298104
rect 300999 298064 301044 298092
rect 301038 298052 301044 298064
rect 301096 298052 301102 298104
rect 393590 298092 393596 298104
rect 393551 298064 393596 298092
rect 393590 298052 393596 298064
rect 393648 298052 393654 298104
rect 460014 298092 460020 298104
rect 459975 298064 460020 298092
rect 460014 298052 460020 298064
rect 460072 298052 460078 298104
rect 288894 297984 288900 298036
rect 288952 297984 288958 298036
rect 580074 296760 580080 296812
rect 580132 296800 580138 296812
rect 580994 296800 581000 296812
rect 580132 296772 581000 296800
rect 580132 296760 580138 296772
rect 580994 296760 581000 296772
rect 581052 296760 581058 296812
rect 259638 296732 259644 296744
rect 259599 296704 259644 296732
rect 259638 296692 259644 296704
rect 259696 296692 259702 296744
rect 262582 296732 262588 296744
rect 262543 296704 262588 296732
rect 262582 296692 262588 296704
rect 262640 296692 262646 296744
rect 267734 296692 267740 296744
rect 267792 296732 267798 296744
rect 268010 296732 268016 296744
rect 267792 296704 268016 296732
rect 267792 296692 267798 296704
rect 268010 296692 268016 296704
rect 268068 296692 268074 296744
rect 580166 296624 580172 296676
rect 580224 296664 580230 296676
rect 580994 296664 581000 296676
rect 580224 296636 581000 296664
rect 580224 296624 580230 296636
rect 580994 296624 581000 296636
rect 581052 296624 581058 296676
rect 267734 296556 267740 296608
rect 267792 296596 267798 296608
rect 267829 296599 267887 296605
rect 267829 296596 267841 296599
rect 267792 296568 267841 296596
rect 267792 296556 267798 296568
rect 267829 296565 267841 296568
rect 267875 296565 267887 296599
rect 267829 296559 267887 296565
rect 291562 296528 291568 296540
rect 291523 296500 291568 296528
rect 291562 296488 291568 296500
rect 291620 296488 291626 296540
rect 289998 294584 290004 294636
rect 290056 294624 290062 294636
rect 290182 294624 290188 294636
rect 290056 294596 290188 294624
rect 290056 294584 290062 294596
rect 290182 294584 290188 294596
rect 290240 294584 290246 294636
rect 265342 293904 265348 293956
rect 265400 293944 265406 293956
rect 265526 293944 265532 293956
rect 265400 293916 265532 293944
rect 265400 293904 265406 293916
rect 265526 293904 265532 293916
rect 265584 293904 265590 293956
rect 310882 293060 310888 293072
rect 310843 293032 310888 293060
rect 310882 293020 310888 293032
rect 310940 293020 310946 293072
rect 299842 292612 299848 292664
rect 299900 292612 299906 292664
rect 306834 292612 306840 292664
rect 306892 292612 306898 292664
rect 295518 292544 295524 292596
rect 295576 292544 295582 292596
rect 239122 292476 239128 292528
rect 239180 292476 239186 292528
rect 291381 292519 291439 292525
rect 291381 292485 291393 292519
rect 291427 292516 291439 292519
rect 291562 292516 291568 292528
rect 291427 292488 291568 292516
rect 291427 292485 291439 292488
rect 291381 292479 291439 292485
rect 291562 292476 291568 292488
rect 291620 292476 291626 292528
rect 295536 292516 295564 292544
rect 299860 292528 299888 292612
rect 306852 292528 306880 292612
rect 295610 292516 295616 292528
rect 295536 292488 295616 292516
rect 295610 292476 295616 292488
rect 295668 292476 295674 292528
rect 299842 292476 299848 292528
rect 299900 292476 299906 292528
rect 301038 292516 301044 292528
rect 300999 292488 301044 292516
rect 301038 292476 301044 292488
rect 301096 292476 301102 292528
rect 306834 292476 306840 292528
rect 306892 292476 306898 292528
rect 239140 292392 239168 292476
rect 239122 292340 239128 292392
rect 239180 292340 239186 292392
rect 337102 290368 337108 290420
rect 337160 290408 337166 290420
rect 337286 290408 337292 290420
rect 337160 290380 337292 290408
rect 337160 290368 337166 290380
rect 337286 290368 337292 290380
rect 337344 290368 337350 290420
rect 235074 289864 235080 289876
rect 235035 289836 235080 289864
rect 235074 289824 235080 289836
rect 235132 289824 235138 289876
rect 236270 289864 236276 289876
rect 236231 289836 236276 289864
rect 236270 289824 236276 289836
rect 236328 289824 236334 289876
rect 247034 289824 247040 289876
rect 247092 289864 247098 289876
rect 247218 289864 247224 289876
rect 247092 289836 247224 289864
rect 247092 289824 247098 289836
rect 247218 289824 247224 289836
rect 247276 289824 247282 289876
rect 270770 289864 270776 289876
rect 270731 289836 270776 289864
rect 270770 289824 270776 289836
rect 270828 289824 270834 289876
rect 324682 289864 324688 289876
rect 324643 289836 324688 289864
rect 324682 289824 324688 289836
rect 324740 289824 324746 289876
rect 372706 289864 372712 289876
rect 372667 289836 372712 289864
rect 372706 289824 372712 289836
rect 372764 289824 372770 289876
rect 375834 289824 375840 289876
rect 375892 289864 375898 289876
rect 375926 289864 375932 289876
rect 375892 289836 375932 289864
rect 375892 289824 375898 289836
rect 375926 289824 375932 289836
rect 375984 289824 375990 289876
rect 377122 289824 377128 289876
rect 377180 289864 377186 289876
rect 377214 289864 377220 289876
rect 377180 289836 377220 289864
rect 377180 289824 377186 289836
rect 377214 289824 377220 289836
rect 377272 289824 377278 289876
rect 289998 289756 290004 289808
rect 290056 289796 290062 289808
rect 290182 289796 290188 289808
rect 290056 289768 290188 289796
rect 290056 289756 290062 289768
rect 290182 289756 290188 289768
rect 290240 289756 290246 289808
rect 341153 289799 341211 289805
rect 341153 289765 341165 289799
rect 341199 289796 341211 289799
rect 341242 289796 341248 289808
rect 341199 289768 341248 289796
rect 341199 289765 341211 289768
rect 341153 289759 341211 289765
rect 341242 289756 341248 289768
rect 341300 289756 341306 289808
rect 367002 289796 367008 289808
rect 366963 289768 367008 289796
rect 367002 289756 367008 289768
rect 367060 289756 367066 289808
rect 389361 289799 389419 289805
rect 389361 289765 389373 289799
rect 389407 289796 389419 289799
rect 389450 289796 389456 289808
rect 389407 289768 389456 289796
rect 389407 289765 389419 289768
rect 389361 289759 389419 289765
rect 389450 289756 389456 289768
rect 389508 289756 389514 289808
rect 272242 289320 272248 289332
rect 272203 289292 272248 289320
rect 272242 289280 272248 289292
rect 272300 289280 272306 289332
rect 244458 288396 244464 288448
rect 244516 288436 244522 288448
rect 244550 288436 244556 288448
rect 244516 288408 244556 288436
rect 244516 288396 244522 288408
rect 244550 288396 244556 288408
rect 244608 288396 244614 288448
rect 251358 288436 251364 288448
rect 251319 288408 251364 288436
rect 251358 288396 251364 288408
rect 251416 288396 251422 288448
rect 266725 288439 266783 288445
rect 266725 288405 266737 288439
rect 266771 288436 266783 288439
rect 266814 288436 266820 288448
rect 266771 288408 266820 288436
rect 266771 288405 266783 288408
rect 266725 288399 266783 288405
rect 266814 288396 266820 288408
rect 266872 288396 266878 288448
rect 330110 288396 330116 288448
rect 330168 288436 330174 288448
rect 330202 288436 330208 288448
rect 330168 288408 330208 288436
rect 330168 288396 330174 288408
rect 330202 288396 330208 288408
rect 330260 288396 330266 288448
rect 331398 288396 331404 288448
rect 331456 288436 331462 288448
rect 331490 288436 331496 288448
rect 331456 288408 331496 288436
rect 331456 288396 331462 288408
rect 331490 288396 331496 288408
rect 331548 288396 331554 288448
rect 460017 288439 460075 288445
rect 460017 288405 460029 288439
rect 460063 288436 460075 288439
rect 460106 288436 460112 288448
rect 460063 288408 460112 288436
rect 460063 288405 460075 288408
rect 460017 288399 460075 288405
rect 460106 288396 460112 288408
rect 460164 288396 460170 288448
rect 272242 288328 272248 288380
rect 272300 288368 272306 288380
rect 272334 288368 272340 288380
rect 272300 288340 272340 288368
rect 272300 288328 272306 288340
rect 272334 288328 272340 288340
rect 272392 288328 272398 288380
rect 337102 288368 337108 288380
rect 337063 288340 337108 288368
rect 337102 288328 337108 288340
rect 337160 288328 337166 288380
rect 267734 287036 267740 287088
rect 267792 287076 267798 287088
rect 267829 287079 267887 287085
rect 267829 287076 267841 287079
rect 267792 287048 267841 287076
rect 267792 287036 267798 287048
rect 267829 287045 267841 287048
rect 267875 287045 267887 287079
rect 267829 287039 267887 287045
rect 323302 287036 323308 287088
rect 323360 287076 323366 287088
rect 323486 287076 323492 287088
rect 323360 287048 323492 287076
rect 323360 287036 323366 287048
rect 323486 287036 323492 287048
rect 323544 287036 323550 287088
rect 580166 287036 580172 287088
rect 580224 287076 580230 287088
rect 580902 287076 580908 287088
rect 580224 287048 580908 287076
rect 580224 287036 580230 287048
rect 580902 287036 580908 287048
rect 580960 287036 580966 287088
rect 325970 286968 325976 287020
rect 326028 287008 326034 287020
rect 326062 287008 326068 287020
rect 326028 286980 326068 287008
rect 326028 286968 326034 286980
rect 326062 286968 326068 286980
rect 326120 286968 326126 287020
rect 288897 284291 288955 284297
rect 288897 284257 288909 284291
rect 288943 284288 288955 284291
rect 288986 284288 288992 284300
rect 288943 284260 288992 284288
rect 288943 284257 288955 284260
rect 288897 284251 288955 284257
rect 288986 284248 288992 284260
rect 289044 284248 289050 284300
rect 270770 282996 270776 283008
rect 270696 282968 270776 282996
rect 270696 282872 270724 282968
rect 270770 282956 270776 282968
rect 270828 282956 270834 283008
rect 295610 282996 295616 283008
rect 295536 282968 295616 282996
rect 295536 282872 295564 282968
rect 295610 282956 295616 282968
rect 295668 282956 295674 283008
rect 460106 282956 460112 283008
rect 460164 282956 460170 283008
rect 357526 282888 357532 282940
rect 357584 282928 357590 282940
rect 357710 282928 357716 282940
rect 357584 282900 357716 282928
rect 357584 282888 357590 282900
rect 357710 282888 357716 282900
rect 357768 282888 357774 282940
rect 431310 282888 431316 282940
rect 431368 282928 431374 282940
rect 431494 282928 431500 282940
rect 431368 282900 431500 282928
rect 431368 282888 431374 282900
rect 431494 282888 431500 282900
rect 431552 282888 431558 282940
rect 270678 282820 270684 282872
rect 270736 282820 270742 282872
rect 295518 282820 295524 282872
rect 295576 282820 295582 282872
rect 460124 282804 460152 282956
rect 310882 282792 310888 282804
rect 310843 282764 310888 282792
rect 310882 282752 310888 282764
rect 310940 282752 310946 282804
rect 460106 282752 460112 282804
rect 460164 282752 460170 282804
rect 266722 280168 266728 280220
rect 266780 280208 266786 280220
rect 266814 280208 266820 280220
rect 266780 280180 266820 280208
rect 266780 280168 266786 280180
rect 266814 280168 266820 280180
rect 266872 280168 266878 280220
rect 294230 280168 294236 280220
rect 294288 280208 294294 280220
rect 294322 280208 294328 280220
rect 294288 280180 294328 280208
rect 294288 280168 294294 280180
rect 294322 280168 294328 280180
rect 294380 280168 294386 280220
rect 327166 280208 327172 280220
rect 327127 280180 327172 280208
rect 327166 280168 327172 280180
rect 327224 280168 327230 280220
rect 341150 280208 341156 280220
rect 341111 280180 341156 280208
rect 341150 280168 341156 280180
rect 341208 280168 341214 280220
rect 367002 280208 367008 280220
rect 366963 280180 367008 280208
rect 367002 280168 367008 280180
rect 367060 280168 367066 280220
rect 389358 280208 389364 280220
rect 389319 280180 389364 280208
rect 389358 280168 389364 280180
rect 389416 280168 389422 280220
rect 393590 280208 393596 280220
rect 393551 280180 393596 280208
rect 393590 280168 393596 280180
rect 393648 280168 393654 280220
rect 3326 280100 3332 280152
rect 3384 280140 3390 280152
rect 15838 280140 15844 280152
rect 3384 280112 15844 280140
rect 3384 280100 3390 280112
rect 15838 280100 15844 280112
rect 15896 280100 15902 280152
rect 235074 280140 235080 280152
rect 235035 280112 235080 280140
rect 235074 280100 235080 280112
rect 235132 280100 235138 280152
rect 236270 280140 236276 280152
rect 236231 280112 236276 280140
rect 236270 280100 236276 280112
rect 236328 280100 236334 280152
rect 250070 280100 250076 280152
rect 250128 280140 250134 280152
rect 250162 280140 250168 280152
rect 250128 280112 250168 280140
rect 250128 280100 250134 280112
rect 250162 280100 250168 280112
rect 250220 280100 250226 280152
rect 270678 280140 270684 280152
rect 270639 280112 270684 280140
rect 270678 280100 270684 280112
rect 270736 280100 270742 280152
rect 273530 280140 273536 280152
rect 273491 280112 273536 280140
rect 273530 280100 273536 280112
rect 273588 280100 273594 280152
rect 281718 280100 281724 280152
rect 281776 280140 281782 280152
rect 281810 280140 281816 280152
rect 281776 280112 281816 280140
rect 281776 280100 281782 280112
rect 281810 280100 281816 280112
rect 281868 280100 281874 280152
rect 284754 280100 284760 280152
rect 284812 280140 284818 280152
rect 284846 280140 284852 280152
rect 284812 280112 284852 280140
rect 284812 280100 284818 280112
rect 284846 280100 284852 280112
rect 284904 280100 284910 280152
rect 372706 280140 372712 280152
rect 372667 280112 372712 280140
rect 372706 280100 372712 280112
rect 372764 280100 372770 280152
rect 375834 280140 375840 280152
rect 375795 280112 375840 280140
rect 375834 280100 375840 280112
rect 375892 280100 375898 280152
rect 377122 280140 377128 280152
rect 377083 280112 377128 280140
rect 377122 280100 377128 280112
rect 377180 280100 377186 280152
rect 460106 280140 460112 280152
rect 460067 280112 460112 280140
rect 460106 280100 460112 280112
rect 460164 280100 460170 280152
rect 329926 278876 329932 278928
rect 329984 278916 329990 278928
rect 330202 278916 330208 278928
rect 329984 278888 330208 278916
rect 329984 278876 329990 278888
rect 330202 278876 330208 278888
rect 330260 278876 330266 278928
rect 331490 278848 331496 278860
rect 331416 278820 331496 278848
rect 327166 278780 327172 278792
rect 327127 278752 327172 278780
rect 327166 278740 327172 278752
rect 327224 278740 327230 278792
rect 331416 278724 331444 278820
rect 331490 278808 331496 278820
rect 331548 278808 331554 278860
rect 337105 278783 337163 278789
rect 337105 278749 337117 278783
rect 337151 278780 337163 278783
rect 337194 278780 337200 278792
rect 337151 278752 337200 278780
rect 337151 278749 337163 278752
rect 337105 278743 337163 278749
rect 337194 278740 337200 278752
rect 337252 278740 337258 278792
rect 310882 278712 310888 278724
rect 310843 278684 310888 278712
rect 310882 278672 310888 278684
rect 310940 278672 310946 278724
rect 331398 278672 331404 278724
rect 331456 278672 331462 278724
rect 393590 278712 393596 278724
rect 393551 278684 393596 278712
rect 393590 278672 393596 278684
rect 393648 278672 393654 278724
rect 296806 277380 296812 277432
rect 296864 277420 296870 277432
rect 296898 277420 296904 277432
rect 296864 277392 296904 277420
rect 296864 277380 296870 277392
rect 296898 277380 296904 277392
rect 296956 277380 296962 277432
rect 331398 277352 331404 277364
rect 331359 277324 331404 277352
rect 331398 277312 331404 277324
rect 331456 277312 331462 277364
rect 580166 277312 580172 277364
rect 580224 277352 580230 277364
rect 580902 277352 580908 277364
rect 580224 277324 580908 277352
rect 580224 277312 580230 277324
rect 580902 277312 580908 277324
rect 580960 277312 580966 277364
rect 294230 275952 294236 276004
rect 294288 275992 294294 276004
rect 294322 275992 294328 276004
rect 294288 275964 294328 275992
rect 294288 275952 294294 275964
rect 294322 275952 294328 275964
rect 294380 275952 294386 276004
rect 296993 275995 297051 276001
rect 296993 275961 297005 275995
rect 297039 275992 297051 275995
rect 297082 275992 297088 276004
rect 297039 275964 297088 275992
rect 297039 275961 297051 275964
rect 296993 275955 297051 275961
rect 297082 275952 297088 275964
rect 297140 275952 297146 276004
rect 270678 275312 270684 275324
rect 270639 275284 270684 275312
rect 270678 275272 270684 275284
rect 270736 275272 270742 275324
rect 463786 275312 463792 275324
rect 463747 275284 463792 275312
rect 463786 275272 463792 275284
rect 463844 275272 463850 275324
rect 288894 274700 288900 274712
rect 288855 274672 288900 274700
rect 288894 274660 288900 274672
rect 288952 274660 288958 274712
rect 291378 274700 291384 274712
rect 291339 274672 291384 274700
rect 291378 274660 291384 274672
rect 291436 274660 291442 274712
rect 250070 273912 250076 273964
rect 250128 273952 250134 273964
rect 250254 273952 250260 273964
rect 250128 273924 250260 273952
rect 250128 273912 250134 273924
rect 250254 273912 250260 273924
rect 250312 273912 250318 273964
rect 323302 273340 323308 273352
rect 323263 273312 323308 273340
rect 323302 273300 323308 273312
rect 323360 273300 323366 273352
rect 337194 273340 337200 273352
rect 337120 273312 337200 273340
rect 301038 273232 301044 273284
rect 301096 273232 301102 273284
rect 239122 273164 239128 273216
rect 239180 273164 239186 273216
rect 301056 273204 301084 273232
rect 337120 273216 337148 273312
rect 337194 273300 337200 273312
rect 337252 273300 337258 273352
rect 301130 273204 301136 273216
rect 301056 273176 301136 273204
rect 301130 273164 301136 273176
rect 301188 273164 301194 273216
rect 337102 273164 337108 273216
rect 337160 273164 337166 273216
rect 239140 273080 239168 273164
rect 460106 273136 460112 273148
rect 460067 273108 460112 273136
rect 460106 273096 460112 273108
rect 460164 273096 460170 273148
rect 239122 273028 239128 273080
rect 239180 273028 239186 273080
rect 299842 270620 299848 270632
rect 299768 270592 299848 270620
rect 299768 270564 299796 270592
rect 299842 270580 299848 270592
rect 299900 270580 299906 270632
rect 235074 270552 235080 270564
rect 235035 270524 235080 270552
rect 235074 270512 235080 270524
rect 235132 270512 235138 270564
rect 236270 270552 236276 270564
rect 236231 270524 236276 270552
rect 236270 270512 236276 270524
rect 236328 270512 236334 270564
rect 247034 270512 247040 270564
rect 247092 270552 247098 270564
rect 247218 270552 247224 270564
rect 247092 270524 247224 270552
rect 247092 270512 247098 270524
rect 247218 270512 247224 270524
rect 247276 270512 247282 270564
rect 251174 270512 251180 270564
rect 251232 270552 251238 270564
rect 251450 270552 251456 270564
rect 251232 270524 251456 270552
rect 251232 270512 251238 270524
rect 251450 270512 251456 270524
rect 251508 270512 251514 270564
rect 273530 270552 273536 270564
rect 273491 270524 273536 270552
rect 273530 270512 273536 270524
rect 273588 270512 273594 270564
rect 299750 270512 299756 270564
rect 299808 270512 299814 270564
rect 302510 270512 302516 270564
rect 302568 270552 302574 270564
rect 302694 270552 302700 270564
rect 302568 270524 302700 270552
rect 302568 270512 302574 270524
rect 302694 270512 302700 270524
rect 302752 270512 302758 270564
rect 327166 270512 327172 270564
rect 327224 270552 327230 270564
rect 327258 270552 327264 270564
rect 327224 270524 327264 270552
rect 327224 270512 327230 270524
rect 327258 270512 327264 270524
rect 327316 270512 327322 270564
rect 372706 270552 372712 270564
rect 372667 270524 372712 270552
rect 372706 270512 372712 270524
rect 372764 270512 372770 270564
rect 375834 270552 375840 270564
rect 375795 270524 375840 270552
rect 375834 270512 375840 270524
rect 375892 270512 375898 270564
rect 377122 270552 377128 270564
rect 377083 270524 377128 270552
rect 377122 270512 377128 270524
rect 377180 270512 377186 270564
rect 463789 270555 463847 270561
rect 463789 270521 463801 270555
rect 463835 270552 463847 270555
rect 463878 270552 463884 270564
rect 463835 270524 463884 270552
rect 463835 270521 463847 270524
rect 463789 270515 463847 270521
rect 463878 270512 463884 270524
rect 463936 270512 463942 270564
rect 286042 270444 286048 270496
rect 286100 270484 286106 270496
rect 286134 270484 286140 270496
rect 286100 270456 286140 270484
rect 286100 270444 286106 270456
rect 286134 270444 286140 270456
rect 286192 270444 286198 270496
rect 341153 270487 341211 270493
rect 341153 270453 341165 270487
rect 341199 270484 341211 270487
rect 341242 270484 341248 270496
rect 341199 270456 341248 270484
rect 341199 270453 341211 270456
rect 341153 270447 341211 270453
rect 341242 270444 341248 270456
rect 341300 270444 341306 270496
rect 367002 270484 367008 270496
rect 366963 270456 367008 270484
rect 367002 270444 367008 270456
rect 367060 270444 367066 270496
rect 389361 270487 389419 270493
rect 389361 270453 389373 270487
rect 389407 270484 389419 270487
rect 389450 270484 389456 270496
rect 389407 270456 389456 270484
rect 389407 270453 389419 270456
rect 389361 270447 389419 270453
rect 389450 270444 389456 270456
rect 389508 270444 389514 270496
rect 460017 270487 460075 270493
rect 460017 270453 460029 270487
rect 460063 270484 460075 270487
rect 460106 270484 460112 270496
rect 460063 270456 460112 270484
rect 460063 270453 460075 270456
rect 460017 270447 460075 270453
rect 460106 270444 460112 270456
rect 460164 270444 460170 270496
rect 245930 269084 245936 269136
rect 245988 269124 245994 269136
rect 246114 269124 246120 269136
rect 245988 269096 246120 269124
rect 245988 269084 245994 269096
rect 246114 269084 246120 269096
rect 246172 269084 246178 269136
rect 259638 269084 259644 269136
rect 259696 269124 259702 269136
rect 259730 269124 259736 269136
rect 259696 269096 259736 269124
rect 259696 269084 259702 269096
rect 259730 269084 259736 269096
rect 259788 269084 259794 269136
rect 265250 269084 265256 269136
rect 265308 269084 265314 269136
rect 290090 269084 290096 269136
rect 290148 269124 290154 269136
rect 290182 269124 290188 269136
rect 290148 269096 290188 269124
rect 290148 269084 290154 269096
rect 290182 269084 290188 269096
rect 290240 269084 290246 269136
rect 295518 269084 295524 269136
rect 295576 269124 295582 269136
rect 295794 269124 295800 269136
rect 295576 269096 295800 269124
rect 295576 269084 295582 269096
rect 295794 269084 295800 269096
rect 295852 269084 295858 269136
rect 265158 269016 265164 269068
rect 265216 269056 265222 269068
rect 265268 269056 265296 269084
rect 265216 269028 265296 269056
rect 265216 269016 265222 269028
rect 324498 267792 324504 267844
rect 324556 267832 324562 267844
rect 324682 267832 324688 267844
rect 324556 267804 324688 267832
rect 324556 267792 324562 267804
rect 324682 267792 324688 267804
rect 324740 267792 324746 267844
rect 323302 267764 323308 267776
rect 323263 267736 323308 267764
rect 323302 267724 323308 267736
rect 323360 267724 323366 267776
rect 325970 267724 325976 267776
rect 326028 267764 326034 267776
rect 326062 267764 326068 267776
rect 326028 267736 326068 267764
rect 326028 267724 326034 267736
rect 326062 267724 326068 267736
rect 326120 267724 326126 267776
rect 329926 267724 329932 267776
rect 329984 267764 329990 267776
rect 330110 267764 330116 267776
rect 329984 267736 330116 267764
rect 329984 267724 329990 267736
rect 330110 267724 330116 267736
rect 330168 267724 330174 267776
rect 331398 267764 331404 267776
rect 331359 267736 331404 267764
rect 331398 267724 331404 267736
rect 331456 267724 331462 267776
rect 296990 266404 296996 266416
rect 296951 266376 296996 266404
rect 296990 266364 296996 266376
rect 297048 266364 297054 266416
rect 294322 266296 294328 266348
rect 294380 266336 294386 266348
rect 294414 266336 294420 266348
rect 294380 266308 294420 266336
rect 294380 266296 294386 266308
rect 294414 266296 294420 266308
rect 294472 266296 294478 266348
rect 250162 264296 250168 264308
rect 250123 264268 250168 264296
rect 250162 264256 250168 264268
rect 250220 264256 250226 264308
rect 266722 263616 266728 263628
rect 266683 263588 266728 263616
rect 266722 263576 266728 263588
rect 266780 263576 266786 263628
rect 270678 263576 270684 263628
rect 270736 263576 270742 263628
rect 357526 263576 357532 263628
rect 357584 263616 357590 263628
rect 357710 263616 357716 263628
rect 357584 263588 357716 263616
rect 357584 263576 357590 263588
rect 357710 263576 357716 263588
rect 357768 263576 357774 263628
rect 431310 263576 431316 263628
rect 431368 263616 431374 263628
rect 431494 263616 431500 263628
rect 431368 263588 431500 263616
rect 431368 263576 431374 263588
rect 431494 263576 431500 263588
rect 431552 263576 431558 263628
rect 270696 263492 270724 263576
rect 270678 263440 270684 263492
rect 270736 263440 270742 263492
rect 310882 263480 310888 263492
rect 310843 263452 310888 263480
rect 310882 263440 310888 263452
rect 310940 263440 310946 263492
rect 296806 262896 296812 262948
rect 296864 262936 296870 262948
rect 296990 262936 296996 262948
rect 296864 262908 296996 262936
rect 296864 262896 296870 262908
rect 296990 262896 296996 262908
rect 297048 262896 297054 262948
rect 272334 260964 272340 260976
rect 272168 260936 272340 260964
rect 247126 260856 247132 260908
rect 247184 260896 247190 260908
rect 247221 260899 247279 260905
rect 247221 260896 247233 260899
rect 247184 260868 247233 260896
rect 247184 260856 247190 260868
rect 247221 260865 247233 260868
rect 247267 260865 247279 260899
rect 247221 260859 247279 260865
rect 235074 260828 235080 260840
rect 235035 260800 235080 260828
rect 235074 260788 235080 260800
rect 235132 260788 235138 260840
rect 236270 260828 236276 260840
rect 236231 260800 236276 260828
rect 236270 260788 236276 260800
rect 236328 260788 236334 260840
rect 270678 260828 270684 260840
rect 270639 260800 270684 260828
rect 270678 260788 270684 260800
rect 270736 260788 270742 260840
rect 272168 260772 272196 260936
rect 272334 260924 272340 260936
rect 272392 260924 272398 260976
rect 327258 260964 327264 260976
rect 327184 260936 327264 260964
rect 281810 260896 281816 260908
rect 281771 260868 281816 260896
rect 281810 260856 281816 260868
rect 281868 260856 281874 260908
rect 324590 260896 324596 260908
rect 324551 260868 324596 260896
rect 324590 260856 324596 260868
rect 324648 260856 324654 260908
rect 273530 260828 273536 260840
rect 273491 260800 273536 260828
rect 273530 260788 273536 260800
rect 273588 260788 273594 260840
rect 327184 260772 327212 260936
rect 327258 260924 327264 260936
rect 327316 260924 327322 260976
rect 460014 260964 460020 260976
rect 459975 260936 460020 260964
rect 460014 260924 460020 260936
rect 460072 260924 460078 260976
rect 341150 260896 341156 260908
rect 341111 260868 341156 260896
rect 341150 260856 341156 260868
rect 341208 260856 341214 260908
rect 367002 260896 367008 260908
rect 366963 260868 367008 260896
rect 367002 260856 367008 260868
rect 367060 260856 367066 260908
rect 389358 260896 389364 260908
rect 389319 260868 389364 260896
rect 389358 260856 389364 260868
rect 389416 260856 389422 260908
rect 393590 260896 393596 260908
rect 393551 260868 393596 260896
rect 393590 260856 393596 260868
rect 393648 260856 393654 260908
rect 372706 260828 372712 260840
rect 372667 260800 372712 260828
rect 372706 260788 372712 260800
rect 372764 260788 372770 260840
rect 375834 260828 375840 260840
rect 375795 260800 375840 260828
rect 375834 260788 375840 260800
rect 375892 260788 375898 260840
rect 377122 260828 377128 260840
rect 377083 260800 377128 260828
rect 377122 260788 377128 260800
rect 377180 260788 377186 260840
rect 460014 260788 460020 260840
rect 460072 260828 460078 260840
rect 460198 260828 460204 260840
rect 460072 260800 460204 260828
rect 460072 260788 460078 260800
rect 460198 260788 460204 260800
rect 460256 260788 460262 260840
rect 463697 260831 463755 260837
rect 463697 260797 463709 260831
rect 463743 260828 463755 260831
rect 463786 260828 463792 260840
rect 463743 260800 463792 260828
rect 463743 260797 463755 260800
rect 463697 260791 463755 260797
rect 463786 260788 463792 260800
rect 463844 260788 463850 260840
rect 272150 260720 272156 260772
rect 272208 260720 272214 260772
rect 327166 260720 327172 260772
rect 327224 260720 327230 260772
rect 247218 259604 247224 259616
rect 247179 259576 247224 259604
rect 247218 259564 247224 259576
rect 247276 259564 247282 259616
rect 244366 259428 244372 259480
rect 244424 259468 244430 259480
rect 244458 259468 244464 259480
rect 244424 259440 244464 259468
rect 244424 259428 244430 259440
rect 244458 259428 244464 259440
rect 244516 259428 244522 259480
rect 250162 259468 250168 259480
rect 250123 259440 250168 259468
rect 250162 259428 250168 259440
rect 250220 259428 250226 259480
rect 266722 259468 266728 259480
rect 266683 259440 266728 259468
rect 266722 259428 266728 259440
rect 266780 259428 266786 259480
rect 281810 259468 281816 259480
rect 281771 259440 281816 259468
rect 281810 259428 281816 259440
rect 281868 259428 281874 259480
rect 284754 259428 284760 259480
rect 284812 259468 284818 259480
rect 284846 259468 284852 259480
rect 284812 259440 284852 259468
rect 284812 259428 284818 259440
rect 284846 259428 284852 259440
rect 284904 259428 284910 259480
rect 337102 259428 337108 259480
rect 337160 259468 337166 259480
rect 337286 259468 337292 259480
rect 337160 259440 337292 259468
rect 337160 259428 337166 259440
rect 337286 259428 337292 259440
rect 337344 259428 337350 259480
rect 331398 259400 331404 259412
rect 331359 259372 331404 259400
rect 331398 259360 331404 259372
rect 331456 259360 331462 259412
rect 288805 259131 288863 259137
rect 288805 259097 288817 259131
rect 288851 259128 288863 259131
rect 288894 259128 288900 259140
rect 288851 259100 288900 259128
rect 288851 259097 288863 259100
rect 288805 259091 288863 259097
rect 288894 259088 288900 259100
rect 288952 259088 288958 259140
rect 324590 258108 324596 258120
rect 324551 258080 324596 258108
rect 324590 258068 324596 258080
rect 324648 258068 324654 258120
rect 247218 258040 247224 258052
rect 247179 258012 247224 258040
rect 247218 258000 247224 258012
rect 247276 258000 247282 258052
rect 262306 258000 262312 258052
rect 262364 258040 262370 258052
rect 262582 258040 262588 258052
rect 262364 258012 262588 258040
rect 262364 258000 262370 258012
rect 262582 258000 262588 258012
rect 262640 258000 262646 258052
rect 291470 258000 291476 258052
rect 291528 258040 291534 258052
rect 291562 258040 291568 258052
rect 291528 258012 291568 258040
rect 291528 258000 291534 258012
rect 291562 258000 291568 258012
rect 291620 258000 291626 258052
rect 295518 258000 295524 258052
rect 295576 258040 295582 258052
rect 295702 258040 295708 258052
rect 295576 258012 295708 258040
rect 295576 258000 295582 258012
rect 295702 258000 295708 258012
rect 295760 258000 295766 258052
rect 330110 258000 330116 258052
rect 330168 258040 330174 258052
rect 330294 258040 330300 258052
rect 330168 258012 330300 258040
rect 330168 258000 330174 258012
rect 330294 258000 330300 258012
rect 330352 258000 330358 258052
rect 296809 257975 296867 257981
rect 296809 257941 296821 257975
rect 296855 257972 296867 257975
rect 296990 257972 296996 257984
rect 296855 257944 296996 257972
rect 296855 257941 296867 257944
rect 296809 257935 296867 257941
rect 296990 257932 296996 257944
rect 297048 257932 297054 257984
rect 310882 256068 310888 256080
rect 310843 256040 310888 256068
rect 310882 256028 310888 256040
rect 310940 256028 310946 256080
rect 270678 256000 270684 256012
rect 270639 255972 270684 256000
rect 270678 255960 270684 255972
rect 270736 255960 270742 256012
rect 286045 255935 286103 255941
rect 286045 255901 286057 255935
rect 286091 255932 286103 255935
rect 286134 255932 286140 255944
rect 286091 255904 286140 255932
rect 286091 255901 286103 255904
rect 286045 255895 286103 255901
rect 286134 255892 286140 255904
rect 286192 255892 286198 255944
rect 259641 254643 259699 254649
rect 259641 254609 259653 254643
rect 259687 254640 259699 254643
rect 259730 254640 259736 254652
rect 259687 254612 259736 254640
rect 259687 254609 259699 254612
rect 259641 254603 259699 254609
rect 259730 254600 259736 254612
rect 259788 254600 259794 254652
rect 323302 253920 323308 253972
rect 323360 253960 323366 253972
rect 323397 253963 323455 253969
rect 323397 253960 323409 253963
rect 323360 253932 323409 253960
rect 323360 253920 323366 253932
rect 323397 253929 323409 253932
rect 323443 253929 323455 253963
rect 323397 253923 323455 253929
rect 337102 253920 337108 253972
rect 337160 253920 337166 253972
rect 239122 253852 239128 253904
rect 239180 253852 239186 253904
rect 239140 253768 239168 253852
rect 337120 253824 337148 253920
rect 337286 253824 337292 253836
rect 337120 253796 337292 253824
rect 337286 253784 337292 253796
rect 337344 253784 337350 253836
rect 239122 253716 239128 253768
rect 239180 253716 239186 253768
rect 294233 251855 294291 251861
rect 294233 251821 294245 251855
rect 294279 251852 294291 251855
rect 294414 251852 294420 251864
rect 294279 251824 294420 251852
rect 294279 251821 294291 251824
rect 294233 251815 294291 251821
rect 294414 251812 294420 251824
rect 294472 251812 294478 251864
rect 367002 251404 367008 251456
rect 367060 251404 367066 251456
rect 310698 251268 310704 251320
rect 310756 251308 310762 251320
rect 310885 251311 310943 251317
rect 310885 251308 310897 251311
rect 310756 251280 310897 251308
rect 310756 251268 310762 251280
rect 310885 251277 310897 251280
rect 310931 251277 310943 251311
rect 310885 251271 310943 251277
rect 366818 251268 366824 251320
rect 366876 251308 366882 251320
rect 366876 251280 366956 251308
rect 366876 251268 366882 251280
rect 366928 251252 366956 251280
rect 367020 251252 367048 251404
rect 235074 251240 235080 251252
rect 235035 251212 235080 251240
rect 235074 251200 235080 251212
rect 235132 251200 235138 251252
rect 236270 251240 236276 251252
rect 236231 251212 236276 251240
rect 236270 251200 236276 251212
rect 236328 251200 236334 251252
rect 251174 251200 251180 251252
rect 251232 251240 251238 251252
rect 251450 251240 251456 251252
rect 251232 251212 251456 251240
rect 251232 251200 251238 251212
rect 251450 251200 251456 251212
rect 251508 251200 251514 251252
rect 273530 251240 273536 251252
rect 273491 251212 273536 251240
rect 273530 251200 273536 251212
rect 273588 251200 273594 251252
rect 289998 251200 290004 251252
rect 290056 251240 290062 251252
rect 290090 251240 290096 251252
rect 290056 251212 290096 251240
rect 290056 251200 290062 251212
rect 290090 251200 290096 251212
rect 290148 251200 290154 251252
rect 366910 251200 366916 251252
rect 366968 251200 366974 251252
rect 367002 251200 367008 251252
rect 367060 251200 367066 251252
rect 372706 251240 372712 251252
rect 372667 251212 372712 251240
rect 372706 251200 372712 251212
rect 372764 251200 372770 251252
rect 375834 251240 375840 251252
rect 375795 251212 375840 251240
rect 375834 251200 375840 251212
rect 375892 251200 375898 251252
rect 377122 251240 377128 251252
rect 377083 251212 377128 251240
rect 377122 251200 377128 251212
rect 377180 251200 377186 251252
rect 389174 251200 389180 251252
rect 389232 251240 389238 251252
rect 389358 251240 389364 251252
rect 389232 251212 389364 251240
rect 389232 251200 389238 251212
rect 389358 251200 389364 251212
rect 389416 251200 389422 251252
rect 463694 251200 463700 251252
rect 463752 251240 463758 251252
rect 463752 251212 463797 251240
rect 463752 251200 463758 251212
rect 250162 251172 250168 251184
rect 250123 251144 250168 251172
rect 250162 251132 250168 251144
rect 250220 251132 250226 251184
rect 281810 251172 281816 251184
rect 281771 251144 281816 251172
rect 281810 251132 281816 251144
rect 281868 251132 281874 251184
rect 284662 251132 284668 251184
rect 284720 251172 284726 251184
rect 284754 251172 284760 251184
rect 284720 251144 284760 251172
rect 284720 251132 284726 251144
rect 284754 251132 284760 251144
rect 284812 251132 284818 251184
rect 310698 251172 310704 251184
rect 310659 251144 310704 251172
rect 310698 251132 310704 251144
rect 310756 251132 310762 251184
rect 460017 251175 460075 251181
rect 460017 251141 460029 251175
rect 460063 251172 460075 251175
rect 460106 251172 460112 251184
rect 460063 251144 460112 251172
rect 460063 251141 460075 251144
rect 460017 251135 460075 251141
rect 460106 251132 460112 251144
rect 460164 251132 460170 251184
rect 367002 251104 367008 251116
rect 366963 251076 367008 251104
rect 367002 251064 367008 251076
rect 367060 251064 367066 251116
rect 301041 249883 301099 249889
rect 301041 249849 301053 249883
rect 301087 249880 301099 249883
rect 301130 249880 301136 249892
rect 301087 249852 301136 249880
rect 301087 249849 301099 249852
rect 301041 249843 301099 249849
rect 301130 249840 301136 249852
rect 301188 249840 301194 249892
rect 330018 249840 330024 249892
rect 330076 249840 330082 249892
rect 245838 249772 245844 249824
rect 245896 249812 245902 249824
rect 246022 249812 246028 249824
rect 245896 249784 246028 249812
rect 245896 249772 245902 249784
rect 246022 249772 246028 249784
rect 246080 249772 246086 249824
rect 299750 249772 299756 249824
rect 299808 249812 299814 249824
rect 299934 249812 299940 249824
rect 299808 249784 299940 249812
rect 299808 249772 299814 249784
rect 299934 249772 299940 249784
rect 299992 249772 299998 249824
rect 302510 249772 302516 249824
rect 302568 249812 302574 249824
rect 302602 249812 302608 249824
rect 302568 249784 302608 249812
rect 302568 249772 302574 249784
rect 302602 249772 302608 249784
rect 302660 249772 302666 249824
rect 306742 249772 306748 249824
rect 306800 249812 306806 249824
rect 306926 249812 306932 249824
rect 306800 249784 306932 249812
rect 306800 249772 306806 249784
rect 306926 249772 306932 249784
rect 306984 249772 306990 249824
rect 323394 249812 323400 249824
rect 323355 249784 323400 249812
rect 323394 249772 323400 249784
rect 323452 249772 323458 249824
rect 330036 249756 330064 249840
rect 393590 249772 393596 249824
rect 393648 249812 393654 249824
rect 393774 249812 393780 249824
rect 393648 249784 393780 249812
rect 393648 249772 393654 249784
rect 393774 249772 393780 249784
rect 393832 249772 393838 249824
rect 247218 249744 247224 249756
rect 247179 249716 247224 249744
rect 247218 249704 247224 249716
rect 247276 249704 247282 249756
rect 330018 249704 330024 249756
rect 330076 249704 330082 249756
rect 296806 249472 296812 249484
rect 296767 249444 296812 249472
rect 296806 249432 296812 249444
rect 296864 249432 296870 249484
rect 301038 248452 301044 248464
rect 300999 248424 301044 248452
rect 301038 248412 301044 248424
rect 301096 248412 301102 248464
rect 284662 248384 284668 248396
rect 284623 248356 284668 248384
rect 284662 248344 284668 248356
rect 284720 248344 284726 248396
rect 306742 248384 306748 248396
rect 306703 248356 306748 248384
rect 306742 248344 306748 248356
rect 306800 248344 306806 248396
rect 286042 247092 286048 247104
rect 286003 247064 286048 247092
rect 286042 247052 286048 247064
rect 286100 247052 286106 247104
rect 329926 244944 329932 244996
rect 329984 244984 329990 244996
rect 330202 244984 330208 244996
rect 329984 244956 330208 244984
rect 329984 244944 329990 244956
rect 330202 244944 330208 244956
rect 330260 244944 330266 244996
rect 341242 244372 341248 244384
rect 341168 244344 341248 244372
rect 341168 244248 341196 244344
rect 341242 244332 341248 244344
rect 341300 244332 341306 244384
rect 357526 244264 357532 244316
rect 357584 244304 357590 244316
rect 357710 244304 357716 244316
rect 357584 244276 357716 244304
rect 357584 244264 357590 244276
rect 357710 244264 357716 244276
rect 357768 244264 357774 244316
rect 431310 244264 431316 244316
rect 431368 244304 431374 244316
rect 431494 244304 431500 244316
rect 431368 244276 431500 244304
rect 431368 244264 431374 244276
rect 431494 244264 431500 244276
rect 431552 244264 431558 244316
rect 341150 244196 341156 244248
rect 341208 244196 341214 244248
rect 259638 241584 259644 241596
rect 259599 241556 259644 241584
rect 259638 241544 259644 241556
rect 259696 241544 259702 241596
rect 250162 241516 250168 241528
rect 250123 241488 250168 241516
rect 250162 241476 250168 241488
rect 250220 241476 250226 241528
rect 266630 241476 266636 241528
rect 266688 241516 266694 241528
rect 266722 241516 266728 241528
rect 266688 241488 266728 241516
rect 266688 241476 266694 241488
rect 266722 241476 266728 241488
rect 266780 241476 266786 241528
rect 281810 241516 281816 241528
rect 281771 241488 281816 241516
rect 281810 241476 281816 241488
rect 281868 241476 281874 241528
rect 288802 241516 288808 241528
rect 288763 241488 288808 241516
rect 288802 241476 288808 241488
rect 288860 241476 288866 241528
rect 289998 241476 290004 241528
rect 290056 241516 290062 241528
rect 290182 241516 290188 241528
rect 290056 241488 290188 241516
rect 290056 241476 290062 241488
rect 290182 241476 290188 241488
rect 290240 241476 290246 241528
rect 291470 241476 291476 241528
rect 291528 241516 291534 241528
rect 291654 241516 291660 241528
rect 291528 241488 291660 241516
rect 291528 241476 291534 241488
rect 291654 241476 291660 241488
rect 291712 241476 291718 241528
rect 310701 241519 310759 241525
rect 310701 241485 310713 241519
rect 310747 241516 310759 241519
rect 310882 241516 310888 241528
rect 310747 241488 310888 241516
rect 310747 241485 310759 241488
rect 310701 241479 310759 241485
rect 310882 241476 310888 241488
rect 310940 241476 310946 241528
rect 367002 241516 367008 241528
rect 366963 241488 367008 241516
rect 367002 241476 367008 241488
rect 367060 241476 367066 241528
rect 460014 241516 460020 241528
rect 459975 241488 460020 241516
rect 460014 241476 460020 241488
rect 460072 241476 460078 241528
rect 270678 241408 270684 241460
rect 270736 241448 270742 241460
rect 270862 241448 270868 241460
rect 270736 241420 270868 241448
rect 270736 241408 270742 241420
rect 270862 241408 270868 241420
rect 270920 241408 270926 241460
rect 272150 241408 272156 241460
rect 272208 241448 272214 241460
rect 272334 241448 272340 241460
rect 272208 241420 272340 241448
rect 272208 241408 272214 241420
rect 272334 241408 272340 241420
rect 272392 241408 272398 241460
rect 299474 241408 299480 241460
rect 299532 241448 299538 241460
rect 375834 241448 375840 241460
rect 299532 241420 299577 241448
rect 375795 241420 375840 241448
rect 299532 241408 299538 241420
rect 375834 241408 375840 241420
rect 375892 241408 375898 241460
rect 463786 241448 463792 241460
rect 463747 241420 463792 241448
rect 463786 241408 463792 241420
rect 463844 241408 463850 241460
rect 244366 240116 244372 240168
rect 244424 240156 244430 240168
rect 244550 240156 244556 240168
rect 244424 240128 244556 240156
rect 244424 240116 244430 240128
rect 244550 240116 244556 240128
rect 244608 240116 244614 240168
rect 245930 240116 245936 240168
rect 245988 240156 245994 240168
rect 246114 240156 246120 240168
rect 245988 240128 246120 240156
rect 245988 240116 245994 240128
rect 246114 240116 246120 240128
rect 246172 240116 246178 240168
rect 251174 240116 251180 240168
rect 251232 240156 251238 240168
rect 251358 240156 251364 240168
rect 251232 240128 251364 240156
rect 251232 240116 251238 240128
rect 251358 240116 251364 240128
rect 251416 240116 251422 240168
rect 262490 240116 262496 240168
rect 262548 240156 262554 240168
rect 262582 240156 262588 240168
rect 262548 240128 262588 240156
rect 262548 240116 262554 240128
rect 262582 240116 262588 240128
rect 262640 240116 262646 240168
rect 267734 240116 267740 240168
rect 267792 240156 267798 240168
rect 267826 240156 267832 240168
rect 267792 240128 267832 240156
rect 267792 240116 267798 240128
rect 267826 240116 267832 240128
rect 267884 240116 267890 240168
rect 299750 240116 299756 240168
rect 299808 240156 299814 240168
rect 299934 240156 299940 240168
rect 299808 240128 299940 240156
rect 299808 240116 299814 240128
rect 299934 240116 299940 240128
rect 299992 240116 299998 240168
rect 301038 240116 301044 240168
rect 301096 240156 301102 240168
rect 301130 240156 301136 240168
rect 301096 240128 301136 240156
rect 301096 240116 301102 240128
rect 301130 240116 301136 240128
rect 301188 240116 301194 240168
rect 302510 240116 302516 240168
rect 302568 240156 302574 240168
rect 302694 240156 302700 240168
rect 302568 240128 302700 240156
rect 302568 240116 302574 240128
rect 302694 240116 302700 240128
rect 302752 240116 302758 240168
rect 306745 240091 306803 240097
rect 306745 240057 306757 240091
rect 306791 240088 306803 240091
rect 306834 240088 306840 240100
rect 306791 240060 306840 240088
rect 306791 240057 306803 240060
rect 306745 240051 306803 240057
rect 306834 240048 306840 240060
rect 306892 240048 306898 240100
rect 284665 238799 284723 238805
rect 284665 238765 284677 238799
rect 284711 238796 284723 238799
rect 284754 238796 284760 238808
rect 284711 238768 284760 238796
rect 284711 238765 284723 238768
rect 284665 238759 284723 238765
rect 284754 238756 284760 238768
rect 284812 238756 284818 238808
rect 294233 238799 294291 238805
rect 294233 238765 294245 238799
rect 294279 238796 294291 238799
rect 294414 238796 294420 238808
rect 294279 238768 294420 238796
rect 294279 238765 294291 238768
rect 294233 238759 294291 238765
rect 294414 238756 294420 238768
rect 294472 238756 294478 238808
rect 285950 238688 285956 238740
rect 286008 238688 286014 238740
rect 393314 238688 393320 238740
rect 393372 238728 393378 238740
rect 393498 238728 393504 238740
rect 393372 238700 393504 238728
rect 393372 238688 393378 238700
rect 393498 238688 393504 238700
rect 393556 238688 393562 238740
rect 285968 238592 285996 238688
rect 286134 238592 286140 238604
rect 285968 238564 286140 238592
rect 286134 238552 286140 238564
rect 286192 238552 286198 238604
rect 3326 237328 3332 237380
rect 3384 237368 3390 237380
rect 17218 237368 17224 237380
rect 3384 237340 17224 237368
rect 3384 237328 3390 237340
rect 17218 237328 17224 237340
rect 17276 237328 17282 237380
rect 331398 236688 331404 236700
rect 331359 236660 331404 236688
rect 331398 236648 331404 236660
rect 331456 236648 331462 236700
rect 267734 234676 267740 234728
rect 267792 234676 267798 234728
rect 281810 234676 281816 234728
rect 281868 234676 281874 234728
rect 310882 234716 310888 234728
rect 310808 234688 310888 234716
rect 244458 234648 244464 234660
rect 244384 234620 244464 234648
rect 244384 234592 244412 234620
rect 244458 234608 244464 234620
rect 244516 234608 244522 234660
rect 250070 234608 250076 234660
rect 250128 234648 250134 234660
rect 250165 234651 250223 234657
rect 250165 234648 250177 234651
rect 250128 234620 250177 234648
rect 250128 234608 250134 234620
rect 250165 234617 250177 234620
rect 250211 234617 250223 234651
rect 250165 234611 250223 234617
rect 267752 234592 267780 234676
rect 281828 234592 281856 234676
rect 310808 234592 310836 234688
rect 310882 234676 310888 234688
rect 310940 234676 310946 234728
rect 463789 234651 463847 234657
rect 463789 234617 463801 234651
rect 463835 234648 463847 234651
rect 463970 234648 463976 234660
rect 463835 234620 463976 234648
rect 463835 234617 463847 234620
rect 463789 234611 463847 234617
rect 463970 234608 463976 234620
rect 464028 234608 464034 234660
rect 239122 234540 239128 234592
rect 239180 234540 239186 234592
rect 244366 234540 244372 234592
rect 244424 234540 244430 234592
rect 267734 234540 267740 234592
rect 267792 234540 267798 234592
rect 281810 234540 281816 234592
rect 281868 234540 281874 234592
rect 310790 234540 310796 234592
rect 310848 234540 310854 234592
rect 239140 234456 239168 234540
rect 239122 234404 239128 234456
rect 239180 234404 239186 234456
rect 323394 233860 323400 233912
rect 323452 233900 323458 233912
rect 323578 233900 323584 233912
rect 323452 233872 323584 233900
rect 323452 233860 323458 233872
rect 323578 233860 323584 233872
rect 323636 233860 323642 233912
rect 302694 231928 302700 231940
rect 302620 231900 302700 231928
rect 234890 231820 234896 231872
rect 234948 231860 234954 231872
rect 235074 231860 235080 231872
rect 234948 231832 235080 231860
rect 234948 231820 234954 231832
rect 235074 231820 235080 231832
rect 235132 231820 235138 231872
rect 236270 231820 236276 231872
rect 236328 231860 236334 231872
rect 236454 231860 236460 231872
rect 236328 231832 236460 231860
rect 236328 231820 236334 231832
rect 236454 231820 236460 231832
rect 236512 231820 236518 231872
rect 273530 231820 273536 231872
rect 273588 231860 273594 231872
rect 273714 231860 273720 231872
rect 273588 231832 273720 231860
rect 273588 231820 273594 231832
rect 273714 231820 273720 231832
rect 273772 231820 273778 231872
rect 299474 231820 299480 231872
rect 299532 231860 299538 231872
rect 299532 231832 299577 231860
rect 299532 231820 299538 231832
rect 301130 231820 301136 231872
rect 301188 231820 301194 231872
rect 301148 231792 301176 231820
rect 302620 231804 302648 231900
rect 302694 231888 302700 231900
rect 302752 231888 302758 231940
rect 306926 231928 306932 231940
rect 306852 231900 306932 231928
rect 306852 231804 306880 231900
rect 306926 231888 306932 231900
rect 306984 231888 306990 231940
rect 324682 231820 324688 231872
rect 324740 231860 324746 231872
rect 324774 231860 324780 231872
rect 324740 231832 324780 231860
rect 324740 231820 324746 231832
rect 324774 231820 324780 231832
rect 324832 231820 324838 231872
rect 325970 231820 325976 231872
rect 326028 231860 326034 231872
rect 326062 231860 326068 231872
rect 326028 231832 326068 231860
rect 326028 231820 326034 231832
rect 326062 231820 326068 231832
rect 326120 231820 326126 231872
rect 327258 231820 327264 231872
rect 327316 231860 327322 231872
rect 327350 231860 327356 231872
rect 327316 231832 327356 231860
rect 327316 231820 327322 231832
rect 327350 231820 327356 231832
rect 327408 231820 327414 231872
rect 372522 231820 372528 231872
rect 372580 231860 372586 231872
rect 372706 231860 372712 231872
rect 372580 231832 372712 231860
rect 372580 231820 372586 231832
rect 372706 231820 372712 231832
rect 372764 231820 372770 231872
rect 375834 231860 375840 231872
rect 375795 231832 375840 231860
rect 375834 231820 375840 231832
rect 375892 231820 375898 231872
rect 376938 231820 376944 231872
rect 376996 231860 377002 231872
rect 377122 231860 377128 231872
rect 376996 231832 377128 231860
rect 376996 231820 377002 231832
rect 377122 231820 377128 231832
rect 377180 231820 377186 231872
rect 301222 231792 301228 231804
rect 301148 231764 301228 231792
rect 301222 231752 301228 231764
rect 301280 231752 301286 231804
rect 302602 231752 302608 231804
rect 302660 231752 302666 231804
rect 306834 231752 306840 231804
rect 306892 231752 306898 231804
rect 310790 231792 310796 231804
rect 310751 231764 310796 231792
rect 310790 231752 310796 231764
rect 310848 231752 310854 231804
rect 367002 231792 367008 231804
rect 366963 231764 367008 231792
rect 367002 231752 367008 231764
rect 367060 231752 367066 231804
rect 250162 230500 250168 230512
rect 250123 230472 250168 230500
rect 250162 230460 250168 230472
rect 250220 230460 250226 230512
rect 251082 230460 251088 230512
rect 251140 230500 251146 230512
rect 251358 230500 251364 230512
rect 251140 230472 251364 230500
rect 251140 230460 251146 230472
rect 251358 230460 251364 230472
rect 251416 230460 251422 230512
rect 259546 230460 259552 230512
rect 259604 230500 259610 230512
rect 259638 230500 259644 230512
rect 259604 230472 259644 230500
rect 259604 230460 259610 230472
rect 259638 230460 259644 230472
rect 259696 230460 259702 230512
rect 270678 230460 270684 230512
rect 270736 230500 270742 230512
rect 270770 230500 270776 230512
rect 270736 230472 270776 230500
rect 270736 230460 270742 230472
rect 270770 230460 270776 230472
rect 270828 230460 270834 230512
rect 288710 230460 288716 230512
rect 288768 230500 288774 230512
rect 288802 230500 288808 230512
rect 288768 230472 288808 230500
rect 288768 230460 288774 230472
rect 288802 230460 288808 230472
rect 288860 230460 288866 230512
rect 330202 230460 330208 230512
rect 330260 230500 330266 230512
rect 330386 230500 330392 230512
rect 330260 230472 330392 230500
rect 330260 230460 330266 230472
rect 330386 230460 330392 230472
rect 330444 230460 330450 230512
rect 341242 230460 341248 230512
rect 341300 230500 341306 230512
rect 341426 230500 341432 230512
rect 341300 230472 341432 230500
rect 341300 230460 341306 230472
rect 341426 230460 341432 230472
rect 341484 230460 341490 230512
rect 337286 225332 337292 225344
rect 337247 225304 337292 225332
rect 337286 225292 337292 225304
rect 337344 225292 337350 225344
rect 341242 225060 341248 225072
rect 341168 225032 341248 225060
rect 270678 224952 270684 225004
rect 270736 224952 270742 225004
rect 288710 224952 288716 225004
rect 288768 224952 288774 225004
rect 270696 224868 270724 224952
rect 270678 224816 270684 224868
rect 270736 224816 270742 224868
rect 288728 224856 288756 224952
rect 341168 224936 341196 225032
rect 341242 225020 341248 225032
rect 341300 225020 341306 225072
rect 460106 225060 460112 225072
rect 460032 225032 460112 225060
rect 357526 224952 357532 225004
rect 357584 224992 357590 225004
rect 357710 224992 357716 225004
rect 357584 224964 357716 224992
rect 357584 224952 357590 224964
rect 357710 224952 357716 224964
rect 357768 224952 357774 225004
rect 431310 224952 431316 225004
rect 431368 224992 431374 225004
rect 431494 224992 431500 225004
rect 431368 224964 431500 224992
rect 431368 224952 431374 224964
rect 431494 224952 431500 224964
rect 431552 224952 431558 225004
rect 460032 224936 460060 225032
rect 460106 225020 460112 225032
rect 460164 225020 460170 225072
rect 341150 224884 341156 224936
rect 341208 224884 341214 224936
rect 460014 224884 460020 224936
rect 460072 224884 460078 224936
rect 288802 224856 288808 224868
rect 288728 224828 288808 224856
rect 288802 224816 288808 224828
rect 288860 224816 288866 224868
rect 393314 224204 393320 224256
rect 393372 224244 393378 224256
rect 393498 224244 393504 224256
rect 393372 224216 393504 224244
rect 393372 224204 393378 224216
rect 393498 224204 393504 224216
rect 393556 224204 393562 224256
rect 2774 223048 2780 223100
rect 2832 223088 2838 223100
rect 5166 223088 5172 223100
rect 2832 223060 5172 223088
rect 2832 223048 2838 223060
rect 5166 223048 5172 223060
rect 5224 223048 5230 223100
rect 325970 222272 325976 222284
rect 325896 222244 325976 222272
rect 325896 222216 325924 222244
rect 325970 222232 325976 222244
rect 326028 222232 326034 222284
rect 327258 222272 327264 222284
rect 327184 222244 327264 222272
rect 327184 222216 327212 222244
rect 327258 222232 327264 222244
rect 327316 222232 327322 222284
rect 265158 222164 265164 222216
rect 265216 222204 265222 222216
rect 265342 222204 265348 222216
rect 265216 222176 265348 222204
rect 265216 222164 265222 222176
rect 265342 222164 265348 222176
rect 265400 222164 265406 222216
rect 294322 222164 294328 222216
rect 294380 222204 294386 222216
rect 294414 222204 294420 222216
rect 294380 222176 294420 222204
rect 294380 222164 294386 222176
rect 294414 222164 294420 222176
rect 294472 222164 294478 222216
rect 295518 222164 295524 222216
rect 295576 222204 295582 222216
rect 295610 222204 295616 222216
rect 295576 222176 295616 222204
rect 295576 222164 295582 222176
rect 295610 222164 295616 222176
rect 295668 222164 295674 222216
rect 296806 222164 296812 222216
rect 296864 222204 296870 222216
rect 296898 222204 296904 222216
rect 296864 222176 296904 222204
rect 296864 222164 296870 222176
rect 296898 222164 296904 222176
rect 296956 222164 296962 222216
rect 301038 222164 301044 222216
rect 301096 222204 301102 222216
rect 301222 222204 301228 222216
rect 301096 222176 301228 222204
rect 301096 222164 301102 222176
rect 301222 222164 301228 222176
rect 301280 222164 301286 222216
rect 310793 222207 310851 222213
rect 310793 222173 310805 222207
rect 310839 222204 310851 222207
rect 310882 222204 310888 222216
rect 310839 222176 310888 222204
rect 310839 222173 310851 222176
rect 310793 222167 310851 222173
rect 310882 222164 310888 222176
rect 310940 222164 310946 222216
rect 325878 222164 325884 222216
rect 325936 222164 325942 222216
rect 327166 222164 327172 222216
rect 327224 222164 327230 222216
rect 330110 222164 330116 222216
rect 330168 222204 330174 222216
rect 330202 222204 330208 222216
rect 330168 222176 330208 222204
rect 330168 222164 330174 222176
rect 330202 222164 330208 222176
rect 330260 222164 330266 222216
rect 331398 222204 331404 222216
rect 331359 222176 331404 222204
rect 331398 222164 331404 222176
rect 331456 222164 331462 222216
rect 337286 222204 337292 222216
rect 337247 222176 337292 222204
rect 337286 222164 337292 222176
rect 337344 222164 337350 222216
rect 367002 222204 367008 222216
rect 366963 222176 367008 222204
rect 367002 222164 367008 222176
rect 367060 222164 367066 222216
rect 389266 222164 389272 222216
rect 389324 222204 389330 222216
rect 389542 222204 389548 222216
rect 389324 222176 389548 222204
rect 389324 222164 389330 222176
rect 389542 222164 389548 222176
rect 389600 222164 389606 222216
rect 463786 222164 463792 222216
rect 463844 222204 463850 222216
rect 464062 222204 464068 222216
rect 463844 222176 464068 222204
rect 463844 222164 463850 222176
rect 464062 222164 464068 222176
rect 464120 222164 464126 222216
rect 270678 222136 270684 222148
rect 270639 222108 270684 222136
rect 270678 222096 270684 222108
rect 270736 222096 270742 222148
rect 272150 222096 272156 222148
rect 272208 222136 272214 222148
rect 272242 222136 272248 222148
rect 272208 222108 272248 222136
rect 272208 222096 272214 222108
rect 272242 222096 272248 222108
rect 272300 222096 272306 222148
rect 375834 222136 375840 222148
rect 375795 222108 375840 222136
rect 375834 222096 375840 222108
rect 375892 222096 375898 222148
rect 291838 220980 291844 220992
rect 291672 220952 291844 220980
rect 290366 220912 290372 220924
rect 290200 220884 290372 220912
rect 290200 220856 290228 220884
rect 290366 220872 290372 220884
rect 290424 220872 290430 220924
rect 291672 220856 291700 220952
rect 291838 220940 291844 220952
rect 291896 220940 291902 220992
rect 245838 220804 245844 220856
rect 245896 220844 245902 220856
rect 246022 220844 246028 220856
rect 245896 220816 246028 220844
rect 245896 220804 245902 220816
rect 246022 220804 246028 220816
rect 246080 220804 246086 220856
rect 251542 220804 251548 220856
rect 251600 220844 251606 220856
rect 251634 220844 251640 220856
rect 251600 220816 251640 220844
rect 251600 220804 251606 220816
rect 251634 220804 251640 220816
rect 251692 220804 251698 220856
rect 290182 220804 290188 220856
rect 290240 220804 290246 220856
rect 291654 220804 291660 220856
rect 291712 220804 291718 220856
rect 331398 220844 331404 220856
rect 331359 220816 331404 220844
rect 331398 220804 331404 220816
rect 331456 220804 331462 220856
rect 244366 220776 244372 220788
rect 244327 220748 244372 220776
rect 244366 220736 244372 220748
rect 244424 220736 244430 220788
rect 341150 220776 341156 220788
rect 341111 220748 341156 220776
rect 341150 220736 341156 220748
rect 341208 220736 341214 220788
rect 290182 219416 290188 219428
rect 290143 219388 290188 219416
rect 290182 219376 290188 219388
rect 290240 219376 290246 219428
rect 291654 219416 291660 219428
rect 291615 219388 291660 219416
rect 291654 219376 291660 219388
rect 291712 219376 291718 219428
rect 317506 219376 317512 219428
rect 317564 219416 317570 219428
rect 317690 219416 317696 219428
rect 317564 219388 317696 219416
rect 317564 219376 317570 219388
rect 317690 219376 317696 219388
rect 317748 219376 317754 219428
rect 310882 215404 310888 215416
rect 310808 215376 310888 215404
rect 301038 215296 301044 215348
rect 301096 215296 301102 215348
rect 239122 215228 239128 215280
rect 239180 215228 239186 215280
rect 239140 215144 239168 215228
rect 301056 215200 301084 215296
rect 310808 215280 310836 215376
rect 310882 215364 310888 215376
rect 310940 215364 310946 215416
rect 389542 215404 389548 215416
rect 389468 215376 389548 215404
rect 389468 215280 389496 215376
rect 389542 215364 389548 215376
rect 389600 215364 389606 215416
rect 464062 215404 464068 215416
rect 463988 215376 464068 215404
rect 463988 215280 464016 215376
rect 464062 215364 464068 215376
rect 464120 215364 464126 215416
rect 310790 215228 310796 215280
rect 310848 215228 310854 215280
rect 341150 215268 341156 215280
rect 341111 215240 341156 215268
rect 341150 215228 341156 215240
rect 341208 215228 341214 215280
rect 389450 215228 389456 215280
rect 389508 215228 389514 215280
rect 459830 215228 459836 215280
rect 459888 215268 459894 215280
rect 460014 215268 460020 215280
rect 459888 215240 460020 215268
rect 459888 215228 459894 215240
rect 460014 215228 460020 215240
rect 460072 215228 460078 215280
rect 463970 215228 463976 215280
rect 464028 215228 464034 215280
rect 301130 215200 301136 215212
rect 301056 215172 301136 215200
rect 301130 215160 301136 215172
rect 301188 215160 301194 215212
rect 239122 215092 239128 215144
rect 239180 215092 239186 215144
rect 299750 213664 299756 213716
rect 299808 213704 299814 213716
rect 299934 213704 299940 213716
rect 299808 213676 299940 213704
rect 299808 213664 299814 213676
rect 299934 213664 299940 213676
rect 299992 213664 299998 213716
rect 306742 213664 306748 213716
rect 306800 213704 306806 213716
rect 306926 213704 306932 213716
rect 306800 213676 306932 213704
rect 306800 213664 306806 213676
rect 306926 213664 306932 213676
rect 306984 213664 306990 213716
rect 330202 212576 330208 212628
rect 330260 212576 330266 212628
rect 234890 212508 234896 212560
rect 234948 212548 234954 212560
rect 235074 212548 235080 212560
rect 234948 212520 235080 212548
rect 234948 212508 234954 212520
rect 235074 212508 235080 212520
rect 235132 212508 235138 212560
rect 236270 212508 236276 212560
rect 236328 212548 236334 212560
rect 236454 212548 236460 212560
rect 236328 212520 236460 212548
rect 236328 212508 236334 212520
rect 236454 212508 236460 212520
rect 236512 212508 236518 212560
rect 245838 212508 245844 212560
rect 245896 212548 245902 212560
rect 245930 212548 245936 212560
rect 245896 212520 245936 212548
rect 245896 212508 245902 212520
rect 245930 212508 245936 212520
rect 245988 212508 245994 212560
rect 250070 212508 250076 212560
rect 250128 212548 250134 212560
rect 250254 212548 250260 212560
rect 250128 212520 250260 212548
rect 250128 212508 250134 212520
rect 250254 212508 250260 212520
rect 250312 212508 250318 212560
rect 270681 212551 270739 212557
rect 270681 212517 270693 212551
rect 270727 212548 270739 212551
rect 270770 212548 270776 212560
rect 270727 212520 270776 212548
rect 270727 212517 270739 212520
rect 270681 212511 270739 212517
rect 270770 212508 270776 212520
rect 270828 212508 270834 212560
rect 273530 212508 273536 212560
rect 273588 212548 273594 212560
rect 273714 212548 273720 212560
rect 273588 212520 273720 212548
rect 273588 212508 273594 212520
rect 273714 212508 273720 212520
rect 273772 212508 273778 212560
rect 281718 212508 281724 212560
rect 281776 212548 281782 212560
rect 281902 212548 281908 212560
rect 281776 212520 281908 212548
rect 281776 212508 281782 212520
rect 281902 212508 281908 212520
rect 281960 212508 281966 212560
rect 284662 212508 284668 212560
rect 284720 212548 284726 212560
rect 284846 212548 284852 212560
rect 284720 212520 284852 212548
rect 284720 212508 284726 212520
rect 284846 212508 284852 212520
rect 284904 212508 284910 212560
rect 324682 212508 324688 212560
rect 324740 212548 324746 212560
rect 324774 212548 324780 212560
rect 324740 212520 324780 212548
rect 324740 212508 324746 212520
rect 324774 212508 324780 212520
rect 324832 212508 324838 212560
rect 325878 212508 325884 212560
rect 325936 212548 325942 212560
rect 325970 212548 325976 212560
rect 325936 212520 325976 212548
rect 325936 212508 325942 212520
rect 325970 212508 325976 212520
rect 326028 212508 326034 212560
rect 327166 212508 327172 212560
rect 327224 212548 327230 212560
rect 327258 212548 327264 212560
rect 327224 212520 327264 212548
rect 327224 212508 327230 212520
rect 327258 212508 327264 212520
rect 327316 212508 327322 212560
rect 330220 212492 330248 212576
rect 372522 212508 372528 212560
rect 372580 212548 372586 212560
rect 372706 212548 372712 212560
rect 372580 212520 372712 212548
rect 372580 212508 372586 212520
rect 372706 212508 372712 212520
rect 372764 212508 372770 212560
rect 375834 212548 375840 212560
rect 375795 212520 375840 212548
rect 375834 212508 375840 212520
rect 375892 212508 375898 212560
rect 376938 212508 376944 212560
rect 376996 212548 377002 212560
rect 377122 212548 377128 212560
rect 376996 212520 377128 212548
rect 376996 212508 377002 212520
rect 377122 212508 377128 212520
rect 377180 212508 377186 212560
rect 244369 212483 244427 212489
rect 244369 212449 244381 212483
rect 244415 212480 244427 212483
rect 244458 212480 244464 212492
rect 244415 212452 244464 212480
rect 244415 212449 244427 212452
rect 244369 212443 244427 212449
rect 244458 212440 244464 212452
rect 244516 212440 244522 212492
rect 286042 212480 286048 212492
rect 286003 212452 286048 212480
rect 286042 212440 286048 212452
rect 286100 212440 286106 212492
rect 310790 212480 310796 212492
rect 310751 212452 310796 212480
rect 310790 212440 310796 212452
rect 310848 212440 310854 212492
rect 330202 212440 330208 212492
rect 330260 212440 330266 212492
rect 367002 212480 367008 212492
rect 366963 212452 367008 212480
rect 367002 212440 367008 212452
rect 367060 212440 367066 212492
rect 262490 212100 262496 212152
rect 262548 212140 262554 212152
rect 262674 212140 262680 212152
rect 262548 212112 262680 212140
rect 262548 212100 262554 212112
rect 262674 212100 262680 212112
rect 262732 212100 262738 212152
rect 246942 211080 246948 211132
rect 247000 211120 247006 211132
rect 247218 211120 247224 211132
rect 247000 211092 247224 211120
rect 247000 211080 247006 211092
rect 247218 211080 247224 211092
rect 247276 211080 247282 211132
rect 249978 211080 249984 211132
rect 250036 211120 250042 211132
rect 250070 211120 250076 211132
rect 250036 211092 250076 211120
rect 250036 211080 250042 211092
rect 250070 211080 250076 211092
rect 250128 211080 250134 211132
rect 290182 211120 290188 211132
rect 290143 211092 290188 211120
rect 290182 211080 290188 211092
rect 290240 211080 290246 211132
rect 330113 211123 330171 211129
rect 330113 211089 330125 211123
rect 330159 211120 330171 211123
rect 330294 211120 330300 211132
rect 330159 211092 330300 211120
rect 330159 211089 330171 211092
rect 330113 211083 330171 211089
rect 330294 211080 330300 211092
rect 330352 211080 330358 211132
rect 317506 209788 317512 209840
rect 317564 209828 317570 209840
rect 317690 209828 317696 209840
rect 317564 209800 317696 209828
rect 317564 209788 317570 209800
rect 317690 209788 317696 209800
rect 317748 209788 317754 209840
rect 460106 205748 460112 205760
rect 460032 205720 460112 205748
rect 281718 205640 281724 205692
rect 281776 205640 281782 205692
rect 284662 205640 284668 205692
rect 284720 205640 284726 205692
rect 288710 205640 288716 205692
rect 288768 205640 288774 205692
rect 357526 205640 357532 205692
rect 357584 205680 357590 205692
rect 357710 205680 357716 205692
rect 357584 205652 357716 205680
rect 357584 205640 357590 205652
rect 357710 205640 357716 205652
rect 357768 205640 357774 205692
rect 431310 205640 431316 205692
rect 431368 205680 431374 205692
rect 431494 205680 431500 205692
rect 431368 205652 431500 205680
rect 431368 205640 431374 205652
rect 431494 205640 431500 205652
rect 431552 205640 431558 205692
rect 281736 205544 281764 205640
rect 281810 205544 281816 205556
rect 281736 205516 281816 205544
rect 281810 205504 281816 205516
rect 281868 205504 281874 205556
rect 284680 205544 284708 205640
rect 288728 205612 288756 205640
rect 460032 205624 460060 205720
rect 460106 205708 460112 205720
rect 460164 205708 460170 205760
rect 288802 205612 288808 205624
rect 288728 205584 288808 205612
rect 288802 205572 288808 205584
rect 288860 205572 288866 205624
rect 460014 205572 460020 205624
rect 460072 205572 460078 205624
rect 284754 205544 284760 205556
rect 284680 205516 284760 205544
rect 284754 205504 284760 205516
rect 284812 205504 284818 205556
rect 393498 204932 393504 204944
rect 393459 204904 393504 204932
rect 393498 204892 393504 204904
rect 393556 204892 393562 204944
rect 291654 204320 291660 204332
rect 291615 204292 291660 204320
rect 291654 204280 291660 204292
rect 291712 204280 291718 204332
rect 331398 202988 331404 203040
rect 331456 202988 331462 203040
rect 325970 202960 325976 202972
rect 325896 202932 325976 202960
rect 325896 202904 325924 202932
rect 325970 202920 325976 202932
rect 326028 202920 326034 202972
rect 327258 202960 327264 202972
rect 327184 202932 327264 202960
rect 327184 202904 327212 202932
rect 327258 202920 327264 202932
rect 327316 202920 327322 202972
rect 331416 202904 331444 202988
rect 244366 202852 244372 202904
rect 244424 202892 244430 202904
rect 244550 202892 244556 202904
rect 244424 202864 244556 202892
rect 244424 202852 244430 202864
rect 244550 202852 244556 202864
rect 244608 202852 244614 202904
rect 245838 202852 245844 202904
rect 245896 202892 245902 202904
rect 245930 202892 245936 202904
rect 245896 202864 245936 202892
rect 245896 202852 245902 202864
rect 245930 202852 245936 202864
rect 245988 202852 245994 202904
rect 262490 202852 262496 202904
rect 262548 202892 262554 202904
rect 262582 202892 262588 202904
rect 262548 202864 262588 202892
rect 262548 202852 262554 202864
rect 262582 202852 262588 202864
rect 262640 202852 262646 202904
rect 270494 202852 270500 202904
rect 270552 202892 270558 202904
rect 270678 202892 270684 202904
rect 270552 202864 270684 202892
rect 270552 202852 270558 202864
rect 270678 202852 270684 202864
rect 270736 202852 270742 202904
rect 286045 202895 286103 202901
rect 286045 202861 286057 202895
rect 286091 202892 286103 202895
rect 286134 202892 286140 202904
rect 286091 202864 286140 202892
rect 286091 202861 286103 202864
rect 286045 202855 286103 202861
rect 286134 202852 286140 202864
rect 286192 202852 286198 202904
rect 294230 202852 294236 202904
rect 294288 202892 294294 202904
rect 294322 202892 294328 202904
rect 294288 202864 294328 202892
rect 294288 202852 294294 202864
rect 294322 202852 294328 202864
rect 294380 202852 294386 202904
rect 295518 202852 295524 202904
rect 295576 202892 295582 202904
rect 295610 202892 295616 202904
rect 295576 202864 295616 202892
rect 295576 202852 295582 202864
rect 295610 202852 295616 202864
rect 295668 202852 295674 202904
rect 296806 202852 296812 202904
rect 296864 202892 296870 202904
rect 296898 202892 296904 202904
rect 296864 202864 296904 202892
rect 296864 202852 296870 202864
rect 296898 202852 296904 202864
rect 296956 202852 296962 202904
rect 299750 202852 299756 202904
rect 299808 202892 299814 202904
rect 299842 202892 299848 202904
rect 299808 202864 299848 202892
rect 299808 202852 299814 202864
rect 299842 202852 299848 202864
rect 299900 202852 299906 202904
rect 301038 202852 301044 202904
rect 301096 202892 301102 202904
rect 301130 202892 301136 202904
rect 301096 202864 301136 202892
rect 301096 202852 301102 202864
rect 301130 202852 301136 202864
rect 301188 202852 301194 202904
rect 302510 202852 302516 202904
rect 302568 202892 302574 202904
rect 302602 202892 302608 202904
rect 302568 202864 302608 202892
rect 302568 202852 302574 202864
rect 302602 202852 302608 202864
rect 302660 202852 302666 202904
rect 306742 202852 306748 202904
rect 306800 202892 306806 202904
rect 306834 202892 306840 202904
rect 306800 202864 306840 202892
rect 306800 202852 306806 202864
rect 306834 202852 306840 202864
rect 306892 202852 306898 202904
rect 310793 202895 310851 202901
rect 310793 202861 310805 202895
rect 310839 202892 310851 202895
rect 310882 202892 310888 202904
rect 310839 202864 310888 202892
rect 310839 202861 310851 202864
rect 310793 202855 310851 202861
rect 310882 202852 310888 202864
rect 310940 202852 310946 202904
rect 325878 202852 325884 202904
rect 325936 202852 325942 202904
rect 327166 202852 327172 202904
rect 327224 202852 327230 202904
rect 331398 202852 331404 202904
rect 331456 202852 331462 202904
rect 337194 202852 337200 202904
rect 337252 202892 337258 202904
rect 337286 202892 337292 202904
rect 337252 202864 337292 202892
rect 337252 202852 337258 202864
rect 337286 202852 337292 202864
rect 337344 202852 337350 202904
rect 341150 202852 341156 202904
rect 341208 202892 341214 202904
rect 341242 202892 341248 202904
rect 341208 202864 341248 202892
rect 341208 202852 341214 202864
rect 341242 202852 341248 202864
rect 341300 202852 341306 202904
rect 367002 202892 367008 202904
rect 366963 202864 367008 202892
rect 367002 202852 367008 202864
rect 367060 202852 367066 202904
rect 389266 202852 389272 202904
rect 389324 202892 389330 202904
rect 389542 202892 389548 202904
rect 389324 202864 389548 202892
rect 389324 202852 389330 202864
rect 389542 202852 389548 202864
rect 389600 202852 389606 202904
rect 463786 202852 463792 202904
rect 463844 202892 463850 202904
rect 464062 202892 464068 202904
rect 463844 202864 464068 202892
rect 463844 202852 463850 202864
rect 464062 202852 464068 202864
rect 464120 202852 464126 202904
rect 330110 202824 330116 202836
rect 330071 202796 330116 202824
rect 330110 202784 330116 202796
rect 330168 202784 330174 202836
rect 375834 202824 375840 202836
rect 375795 202796 375840 202824
rect 375834 202784 375840 202796
rect 375892 202784 375898 202836
rect 250070 201424 250076 201476
rect 250128 201464 250134 201476
rect 250162 201464 250168 201476
rect 250128 201436 250168 201464
rect 250128 201424 250134 201436
rect 250162 201424 250168 201436
rect 250220 201424 250226 201476
rect 306834 201424 306840 201476
rect 306892 201464 306898 201476
rect 306926 201464 306932 201476
rect 306892 201436 306932 201464
rect 306892 201424 306898 201436
rect 306926 201424 306932 201436
rect 306984 201424 306990 201476
rect 324590 201464 324596 201476
rect 324551 201436 324596 201464
rect 324590 201424 324596 201436
rect 324648 201424 324654 201476
rect 327166 201464 327172 201476
rect 327127 201436 327172 201464
rect 327166 201424 327172 201436
rect 327224 201424 327230 201476
rect 330110 201424 330116 201476
rect 330168 201464 330174 201476
rect 330294 201464 330300 201476
rect 330168 201436 330300 201464
rect 330168 201424 330174 201436
rect 330294 201424 330300 201436
rect 330352 201424 330358 201476
rect 250070 200064 250076 200116
rect 250128 200104 250134 200116
rect 250254 200104 250260 200116
rect 250128 200076 250260 200104
rect 250128 200064 250134 200076
rect 250254 200064 250260 200076
rect 250312 200064 250318 200116
rect 290001 200107 290059 200113
rect 290001 200073 290013 200107
rect 290047 200104 290059 200107
rect 290182 200104 290188 200116
rect 290047 200076 290188 200104
rect 290047 200073 290059 200076
rect 290001 200067 290059 200073
rect 290182 200064 290188 200076
rect 290240 200064 290246 200116
rect 317506 200064 317512 200116
rect 317564 200104 317570 200116
rect 317690 200104 317696 200116
rect 317564 200076 317696 200104
rect 317564 200064 317570 200076
rect 317690 200064 317696 200076
rect 317748 200064 317754 200116
rect 330294 200064 330300 200116
rect 330352 200104 330358 200116
rect 330478 200104 330484 200116
rect 330352 200076 330484 200104
rect 330352 200064 330358 200076
rect 330478 200064 330484 200076
rect 330536 200064 330542 200116
rect 331398 200104 331404 200116
rect 331359 200076 331404 200104
rect 331398 200064 331404 200076
rect 331456 200064 331462 200116
rect 266722 198092 266728 198144
rect 266780 198092 266786 198144
rect 266740 198008 266768 198092
rect 266722 197956 266728 198008
rect 266780 197956 266786 198008
rect 299842 196092 299848 196104
rect 299768 196064 299848 196092
rect 232222 195984 232228 196036
rect 232280 195984 232286 196036
rect 232240 195956 232268 195984
rect 299768 195968 299796 196064
rect 299842 196052 299848 196064
rect 299900 196052 299906 196104
rect 302602 196092 302608 196104
rect 302528 196064 302608 196092
rect 301038 195984 301044 196036
rect 301096 195984 301102 196036
rect 232314 195956 232320 195968
rect 232240 195928 232320 195956
rect 232314 195916 232320 195928
rect 232372 195916 232378 195968
rect 235074 195916 235080 195968
rect 235132 195916 235138 195968
rect 299750 195916 299756 195968
rect 299808 195916 299814 195968
rect 235092 195832 235120 195916
rect 301056 195888 301084 195984
rect 302528 195968 302556 196064
rect 302602 196052 302608 196064
rect 302660 196052 302666 196104
rect 310882 196092 310888 196104
rect 310808 196064 310888 196092
rect 310808 195968 310836 196064
rect 310882 196052 310888 196064
rect 310940 196052 310946 196104
rect 337194 196092 337200 196104
rect 337120 196064 337200 196092
rect 337120 195968 337148 196064
rect 337194 196052 337200 196064
rect 337252 196052 337258 196104
rect 389542 196092 389548 196104
rect 389468 196064 389548 196092
rect 389468 195968 389496 196064
rect 389542 196052 389548 196064
rect 389600 196052 389606 196104
rect 464062 196092 464068 196104
rect 463988 196064 464068 196092
rect 460014 195984 460020 196036
rect 460072 195984 460078 196036
rect 302510 195916 302516 195968
rect 302568 195916 302574 195968
rect 310790 195916 310796 195968
rect 310848 195916 310854 195968
rect 337102 195916 337108 195968
rect 337160 195916 337166 195968
rect 389450 195916 389456 195968
rect 389508 195916 389514 195968
rect 301130 195888 301136 195900
rect 301056 195860 301136 195888
rect 301130 195848 301136 195860
rect 301188 195848 301194 195900
rect 460032 195888 460060 195984
rect 463988 195968 464016 196064
rect 464062 196052 464068 196064
rect 464120 196052 464126 196104
rect 463970 195916 463976 195968
rect 464028 195916 464034 195968
rect 460106 195888 460112 195900
rect 460032 195860 460112 195888
rect 460106 195848 460112 195860
rect 460164 195848 460170 195900
rect 235074 195780 235080 195832
rect 235132 195780 235138 195832
rect 230842 193196 230848 193248
rect 230900 193236 230906 193248
rect 231026 193236 231032 193248
rect 230900 193208 231032 193236
rect 230900 193196 230906 193208
rect 231026 193196 231032 193208
rect 231084 193196 231090 193248
rect 236270 193196 236276 193248
rect 236328 193236 236334 193248
rect 236454 193236 236460 193248
rect 236328 193208 236460 193236
rect 236328 193196 236334 193208
rect 236454 193196 236460 193208
rect 236512 193196 236518 193248
rect 244366 193196 244372 193248
rect 244424 193236 244430 193248
rect 244458 193236 244464 193248
rect 244424 193208 244464 193236
rect 244424 193196 244430 193208
rect 244458 193196 244464 193208
rect 244516 193196 244522 193248
rect 247126 193196 247132 193248
rect 247184 193236 247190 193248
rect 247218 193236 247224 193248
rect 247184 193208 247224 193236
rect 247184 193196 247190 193208
rect 247218 193196 247224 193208
rect 247276 193196 247282 193248
rect 259730 193196 259736 193248
rect 259788 193236 259794 193248
rect 259914 193236 259920 193248
rect 259788 193208 259920 193236
rect 259788 193196 259794 193208
rect 259914 193196 259920 193208
rect 259972 193196 259978 193248
rect 265250 193196 265256 193248
rect 265308 193236 265314 193248
rect 265342 193236 265348 193248
rect 265308 193208 265348 193236
rect 265308 193196 265314 193208
rect 265342 193196 265348 193208
rect 265400 193196 265406 193248
rect 267826 193196 267832 193248
rect 267884 193236 267890 193248
rect 267918 193236 267924 193248
rect 267884 193208 267924 193236
rect 267884 193196 267890 193208
rect 267918 193196 267924 193208
rect 267976 193196 267982 193248
rect 270494 193196 270500 193248
rect 270552 193236 270558 193248
rect 270770 193236 270776 193248
rect 270552 193208 270776 193236
rect 270552 193196 270558 193208
rect 270770 193196 270776 193208
rect 270828 193196 270834 193248
rect 273530 193196 273536 193248
rect 273588 193236 273594 193248
rect 273714 193236 273720 193248
rect 273588 193208 273720 193236
rect 273588 193196 273594 193208
rect 273714 193196 273720 193208
rect 273772 193196 273778 193248
rect 281718 193196 281724 193248
rect 281776 193236 281782 193248
rect 281902 193236 281908 193248
rect 281776 193208 281908 193236
rect 281776 193196 281782 193208
rect 281902 193196 281908 193208
rect 281960 193196 281966 193248
rect 284662 193196 284668 193248
rect 284720 193236 284726 193248
rect 284846 193236 284852 193248
rect 284720 193208 284852 193236
rect 284720 193196 284726 193208
rect 284846 193196 284852 193208
rect 284904 193196 284910 193248
rect 288710 193196 288716 193248
rect 288768 193236 288774 193248
rect 288894 193236 288900 193248
rect 288768 193208 288900 193236
rect 288768 193196 288774 193208
rect 288894 193196 288900 193208
rect 288952 193196 288958 193248
rect 341242 193196 341248 193248
rect 341300 193236 341306 193248
rect 341426 193236 341432 193248
rect 341300 193208 341432 193236
rect 341300 193196 341306 193208
rect 341426 193196 341432 193208
rect 341484 193196 341490 193248
rect 372522 193196 372528 193248
rect 372580 193236 372586 193248
rect 372706 193236 372712 193248
rect 372580 193208 372712 193236
rect 372580 193196 372586 193208
rect 372706 193196 372712 193208
rect 372764 193196 372770 193248
rect 375834 193236 375840 193248
rect 375795 193208 375840 193236
rect 375834 193196 375840 193208
rect 375892 193196 375898 193248
rect 376938 193196 376944 193248
rect 376996 193236 377002 193248
rect 377122 193236 377128 193248
rect 376996 193208 377128 193236
rect 376996 193196 377002 193208
rect 377122 193196 377128 193208
rect 377180 193196 377186 193248
rect 324593 193171 324651 193177
rect 324593 193137 324605 193171
rect 324639 193168 324651 193171
rect 324682 193168 324688 193180
rect 324639 193140 324688 193168
rect 324639 193137 324651 193140
rect 324593 193131 324651 193137
rect 324682 193128 324688 193140
rect 324740 193128 324746 193180
rect 327169 193171 327227 193177
rect 327169 193137 327181 193171
rect 327215 193168 327227 193171
rect 327258 193168 327264 193180
rect 327215 193140 327264 193168
rect 327215 193137 327227 193140
rect 327169 193131 327227 193137
rect 327258 193128 327264 193140
rect 327316 193128 327322 193180
rect 367002 193168 367008 193180
rect 366963 193140 367008 193168
rect 367002 193128 367008 193140
rect 367060 193128 367066 193180
rect 393498 193100 393504 193112
rect 393459 193072 393504 193100
rect 393498 193060 393504 193072
rect 393556 193060 393562 193112
rect 245838 191876 245844 191888
rect 245799 191848 245844 191876
rect 245838 191836 245844 191848
rect 245896 191836 245902 191888
rect 285950 191768 285956 191820
rect 286008 191808 286014 191820
rect 286042 191808 286048 191820
rect 286008 191780 286048 191808
rect 286008 191768 286014 191780
rect 286042 191768 286048 191780
rect 286100 191768 286106 191820
rect 331401 191811 331459 191817
rect 331401 191777 331413 191811
rect 331447 191808 331459 191811
rect 331582 191808 331588 191820
rect 331447 191780 331588 191808
rect 331447 191777 331459 191780
rect 331401 191771 331459 191777
rect 331582 191768 331588 191780
rect 331640 191768 331646 191820
rect 337102 191808 337108 191820
rect 337063 191780 337108 191808
rect 337102 191768 337108 191780
rect 337160 191768 337166 191820
rect 393498 191808 393504 191820
rect 393459 191780 393504 191808
rect 393498 191768 393504 191780
rect 393556 191768 393562 191820
rect 289998 190516 290004 190528
rect 289959 190488 290004 190516
rect 289998 190476 290004 190488
rect 290056 190476 290062 190528
rect 317506 190476 317512 190528
rect 317564 190516 317570 190528
rect 317690 190516 317696 190528
rect 317564 190488 317696 190516
rect 317564 190476 317570 190488
rect 317690 190476 317696 190488
rect 317748 190476 317754 190528
rect 267734 190408 267740 190460
rect 267792 190448 267798 190460
rect 267826 190448 267832 190460
rect 267792 190420 267832 190448
rect 267792 190408 267798 190420
rect 267826 190408 267832 190420
rect 267884 190408 267890 190460
rect 331398 190408 331404 190460
rect 331456 190448 331462 190460
rect 331674 190448 331680 190460
rect 331456 190420 331680 190448
rect 331456 190408 331462 190420
rect 331674 190408 331680 190420
rect 331732 190408 331738 190460
rect 245378 189048 245384 189100
rect 245436 189088 245442 189100
rect 245841 189091 245899 189097
rect 245841 189088 245853 189091
rect 245436 189060 245853 189088
rect 245436 189048 245442 189060
rect 245841 189057 245853 189060
rect 245887 189057 245899 189091
rect 245841 189051 245899 189057
rect 289998 188300 290004 188352
rect 290056 188300 290062 188352
rect 290016 188216 290044 188300
rect 289998 188164 290004 188216
rect 290056 188164 290062 188216
rect 339770 186940 339776 186992
rect 339828 186980 339834 186992
rect 339954 186980 339960 186992
rect 339828 186952 339960 186980
rect 339828 186940 339834 186952
rect 339954 186940 339960 186952
rect 340012 186940 340018 186992
rect 296898 186436 296904 186448
rect 296824 186408 296904 186436
rect 251358 186328 251364 186380
rect 251416 186328 251422 186380
rect 266630 186328 266636 186380
rect 266688 186328 266694 186380
rect 295610 186368 295616 186380
rect 295536 186340 295616 186368
rect 251376 186244 251404 186328
rect 251358 186192 251364 186244
rect 251416 186192 251422 186244
rect 266648 186232 266676 186328
rect 295536 186312 295564 186340
rect 295610 186328 295616 186340
rect 295668 186328 295674 186380
rect 296824 186312 296852 186408
rect 296898 186396 296904 186408
rect 296956 186396 296962 186448
rect 357526 186328 357532 186380
rect 357584 186368 357590 186380
rect 357710 186368 357716 186380
rect 357584 186340 357716 186368
rect 357584 186328 357590 186340
rect 357710 186328 357716 186340
rect 357768 186328 357774 186380
rect 431310 186328 431316 186380
rect 431368 186368 431374 186380
rect 431494 186368 431500 186380
rect 431368 186340 431500 186368
rect 431368 186328 431374 186340
rect 431494 186328 431500 186340
rect 431552 186328 431558 186380
rect 460014 186328 460020 186380
rect 460072 186368 460078 186380
rect 460072 186340 460152 186368
rect 460072 186328 460078 186340
rect 460124 186312 460152 186340
rect 295518 186260 295524 186312
rect 295576 186260 295582 186312
rect 296806 186260 296812 186312
rect 296864 186260 296870 186312
rect 337102 186300 337108 186312
rect 337063 186272 337108 186300
rect 337102 186260 337108 186272
rect 337160 186260 337166 186312
rect 460106 186260 460112 186312
rect 460164 186260 460170 186312
rect 266722 186232 266728 186244
rect 266648 186204 266728 186232
rect 266722 186192 266728 186204
rect 266780 186192 266786 186244
rect 264974 183540 264980 183592
rect 265032 183580 265038 183592
rect 265158 183580 265164 183592
rect 265032 183552 265164 183580
rect 265032 183540 265038 183552
rect 265158 183540 265164 183552
rect 265216 183540 265222 183592
rect 270494 183540 270500 183592
rect 270552 183580 270558 183592
rect 270678 183580 270684 183592
rect 270552 183552 270684 183580
rect 270552 183540 270558 183552
rect 270678 183540 270684 183552
rect 270736 183540 270742 183592
rect 291562 183540 291568 183592
rect 291620 183580 291626 183592
rect 291654 183580 291660 183592
rect 291620 183552 291660 183580
rect 291620 183540 291626 183552
rect 291654 183540 291660 183552
rect 291712 183540 291718 183592
rect 299750 183540 299756 183592
rect 299808 183580 299814 183592
rect 299842 183580 299848 183592
rect 299808 183552 299848 183580
rect 299808 183540 299814 183552
rect 299842 183540 299848 183552
rect 299900 183540 299906 183592
rect 301038 183540 301044 183592
rect 301096 183580 301102 183592
rect 301130 183580 301136 183592
rect 301096 183552 301136 183580
rect 301096 183540 301102 183552
rect 301130 183540 301136 183552
rect 301188 183540 301194 183592
rect 302510 183540 302516 183592
rect 302568 183580 302574 183592
rect 302602 183580 302608 183592
rect 302568 183552 302608 183580
rect 302568 183540 302574 183552
rect 302602 183540 302608 183552
rect 302660 183540 302666 183592
rect 306834 183540 306840 183592
rect 306892 183580 306898 183592
rect 306926 183580 306932 183592
rect 306892 183552 306932 183580
rect 306892 183540 306898 183552
rect 306926 183540 306932 183552
rect 306984 183540 306990 183592
rect 310882 183540 310888 183592
rect 310940 183580 310946 183592
rect 311066 183580 311072 183592
rect 310940 183552 311072 183580
rect 310940 183540 310946 183552
rect 311066 183540 311072 183552
rect 311124 183540 311130 183592
rect 324590 183540 324596 183592
rect 324648 183580 324654 183592
rect 324774 183580 324780 183592
rect 324648 183552 324780 183580
rect 324648 183540 324654 183552
rect 324774 183540 324780 183552
rect 324832 183540 324838 183592
rect 327166 183540 327172 183592
rect 327224 183580 327230 183592
rect 327350 183580 327356 183592
rect 327224 183552 327356 183580
rect 327224 183540 327230 183552
rect 327350 183540 327356 183552
rect 327408 183540 327414 183592
rect 367002 183580 367008 183592
rect 366963 183552 367008 183580
rect 367002 183540 367008 183552
rect 367060 183540 367066 183592
rect 389266 183540 389272 183592
rect 389324 183580 389330 183592
rect 389542 183580 389548 183592
rect 389324 183552 389548 183580
rect 389324 183540 389330 183552
rect 389542 183540 389548 183552
rect 389600 183540 389606 183592
rect 463786 183540 463792 183592
rect 463844 183580 463850 183592
rect 464062 183580 464068 183592
rect 463844 183552 464068 183580
rect 463844 183540 463850 183552
rect 464062 183540 464068 183552
rect 464120 183540 464126 183592
rect 251358 183472 251364 183524
rect 251416 183512 251422 183524
rect 251542 183512 251548 183524
rect 251416 183484 251548 183512
rect 251416 183472 251422 183484
rect 251542 183472 251548 183484
rect 251600 183472 251606 183524
rect 393498 183512 393504 183524
rect 393459 183484 393504 183512
rect 393498 183472 393504 183484
rect 393556 183472 393562 183524
rect 460106 183512 460112 183524
rect 460067 183484 460112 183512
rect 460106 183472 460112 183484
rect 460164 183472 460170 183524
rect 272058 182112 272064 182164
rect 272116 182152 272122 182164
rect 272334 182152 272340 182164
rect 272116 182124 272340 182152
rect 272116 182112 272122 182124
rect 272334 182112 272340 182124
rect 272392 182112 272398 182164
rect 273533 182155 273591 182161
rect 273533 182121 273545 182155
rect 273579 182152 273591 182155
rect 273714 182152 273720 182164
rect 273579 182124 273720 182152
rect 273579 182121 273591 182124
rect 273533 182115 273591 182121
rect 273714 182112 273720 182124
rect 273772 182112 273778 182164
rect 289998 182152 290004 182164
rect 289959 182124 290004 182152
rect 289998 182112 290004 182124
rect 290056 182112 290062 182164
rect 291654 182152 291660 182164
rect 291615 182124 291660 182152
rect 291654 182112 291660 182124
rect 291712 182112 291718 182164
rect 341150 182112 341156 182164
rect 341208 182152 341214 182164
rect 341242 182152 341248 182164
rect 341208 182124 341248 182152
rect 341208 182112 341214 182124
rect 341242 182112 341248 182124
rect 341300 182112 341306 182164
rect 393314 182112 393320 182164
rect 393372 182152 393378 182164
rect 393498 182152 393504 182164
rect 393372 182124 393504 182152
rect 393372 182112 393378 182124
rect 393498 182112 393504 182124
rect 393556 182112 393562 182164
rect 329926 182044 329932 182096
rect 329984 182084 329990 182096
rect 330110 182084 330116 182096
rect 329984 182056 330116 182084
rect 329984 182044 329990 182056
rect 330110 182044 330116 182056
rect 330168 182044 330174 182096
rect 245746 180928 245752 180940
rect 245707 180900 245752 180928
rect 245746 180888 245752 180900
rect 245804 180888 245810 180940
rect 245654 180820 245660 180872
rect 245712 180820 245718 180872
rect 245672 180736 245700 180820
rect 267826 180752 267832 180804
rect 267884 180792 267890 180804
rect 267918 180792 267924 180804
rect 267884 180764 267924 180792
rect 267884 180752 267890 180764
rect 267918 180752 267924 180764
rect 267976 180752 267982 180804
rect 301038 180792 301044 180804
rect 300999 180764 301044 180792
rect 301038 180752 301044 180764
rect 301096 180752 301102 180804
rect 306834 180792 306840 180804
rect 306795 180764 306840 180792
rect 306834 180752 306840 180764
rect 306892 180752 306898 180804
rect 317506 180752 317512 180804
rect 317564 180792 317570 180804
rect 317690 180792 317696 180804
rect 317564 180764 317696 180792
rect 317564 180752 317570 180764
rect 317690 180752 317696 180764
rect 317748 180752 317754 180804
rect 245654 180684 245660 180736
rect 245712 180684 245718 180736
rect 245378 180616 245384 180668
rect 245436 180656 245442 180668
rect 245838 180656 245844 180668
rect 245436 180628 245844 180656
rect 245436 180616 245442 180628
rect 245838 180616 245844 180628
rect 245896 180616 245902 180668
rect 245746 179432 245752 179444
rect 245707 179404 245752 179432
rect 245746 179392 245752 179404
rect 245804 179392 245810 179444
rect 267826 179364 267832 179376
rect 267787 179336 267832 179364
rect 267826 179324 267832 179336
rect 267884 179324 267890 179376
rect 266722 178780 266728 178832
rect 266780 178780 266786 178832
rect 266740 178696 266768 178780
rect 294230 178712 294236 178764
rect 294288 178752 294294 178764
rect 294414 178752 294420 178764
rect 294288 178724 294420 178752
rect 294288 178712 294294 178724
rect 294414 178712 294420 178724
rect 294472 178712 294478 178764
rect 295518 178712 295524 178764
rect 295576 178752 295582 178764
rect 295702 178752 295708 178764
rect 295576 178724 295708 178752
rect 295576 178712 295582 178724
rect 295702 178712 295708 178724
rect 295760 178712 295766 178764
rect 296806 178712 296812 178764
rect 296864 178752 296870 178764
rect 296990 178752 296996 178764
rect 296864 178724 296996 178752
rect 296864 178712 296870 178724
rect 296990 178712 296996 178724
rect 297048 178712 297054 178764
rect 266722 178644 266728 178696
rect 266780 178644 266786 178696
rect 247126 176740 247132 176792
rect 247184 176740 247190 176792
rect 250254 176780 250260 176792
rect 250088 176752 250260 176780
rect 232222 176672 232228 176724
rect 232280 176672 232286 176724
rect 247144 176712 247172 176740
rect 250088 176724 250116 176752
rect 250254 176740 250260 176752
rect 250312 176740 250318 176792
rect 299842 176780 299848 176792
rect 299803 176752 299848 176780
rect 299842 176740 299848 176752
rect 299900 176740 299906 176792
rect 302602 176740 302608 176792
rect 302660 176740 302666 176792
rect 310882 176780 310888 176792
rect 310808 176752 310888 176780
rect 247218 176712 247224 176724
rect 247144 176684 247224 176712
rect 247218 176672 247224 176684
rect 247276 176672 247282 176724
rect 250070 176672 250076 176724
rect 250128 176672 250134 176724
rect 232240 176644 232268 176672
rect 302620 176656 302648 176740
rect 310808 176656 310836 176752
rect 310882 176740 310888 176752
rect 310940 176740 310946 176792
rect 389542 176780 389548 176792
rect 389468 176752 389548 176780
rect 389468 176656 389496 176752
rect 389542 176740 389548 176752
rect 389600 176740 389606 176792
rect 232314 176644 232320 176656
rect 232240 176616 232320 176644
rect 232314 176604 232320 176616
rect 232372 176604 232378 176656
rect 235074 176604 235080 176656
rect 235132 176604 235138 176656
rect 302602 176604 302608 176656
rect 302660 176604 302666 176656
rect 310790 176604 310796 176656
rect 310848 176604 310854 176656
rect 389450 176604 389456 176656
rect 389508 176604 389514 176656
rect 235092 176520 235120 176604
rect 235074 176468 235080 176520
rect 235132 176468 235138 176520
rect 239122 176468 239128 176520
rect 239180 176468 239186 176520
rect 460106 176508 460112 176520
rect 460067 176480 460112 176508
rect 460106 176468 460112 176480
rect 460164 176468 460170 176520
rect 239140 176384 239168 176468
rect 372706 176400 372712 176452
rect 372764 176440 372770 176452
rect 372798 176440 372804 176452
rect 372764 176412 372804 176440
rect 372764 176400 372770 176412
rect 372798 176400 372804 176412
rect 372856 176400 372862 176452
rect 375834 176400 375840 176452
rect 375892 176440 375898 176452
rect 375926 176440 375932 176452
rect 375892 176412 375932 176440
rect 375892 176400 375898 176412
rect 375926 176400 375932 176412
rect 375984 176400 375990 176452
rect 239122 176332 239128 176384
rect 239180 176332 239186 176384
rect 366818 174020 366824 174072
rect 366876 174060 366882 174072
rect 367002 174060 367008 174072
rect 366876 174032 367008 174060
rect 366876 174020 366882 174032
rect 367002 174020 367008 174032
rect 367060 174020 367066 174072
rect 230842 173884 230848 173936
rect 230900 173924 230906 173936
rect 231026 173924 231032 173936
rect 230900 173896 231032 173924
rect 230900 173884 230906 173896
rect 231026 173884 231032 173896
rect 231084 173884 231090 173936
rect 236270 173884 236276 173936
rect 236328 173924 236334 173936
rect 236454 173924 236460 173936
rect 236328 173896 236460 173924
rect 236328 173884 236334 173896
rect 236454 173884 236460 173896
rect 236512 173884 236518 173936
rect 259730 173884 259736 173936
rect 259788 173924 259794 173936
rect 259914 173924 259920 173936
rect 259788 173896 259920 173924
rect 259788 173884 259794 173896
rect 259914 173884 259920 173896
rect 259972 173884 259978 173936
rect 265250 173884 265256 173936
rect 265308 173924 265314 173936
rect 265342 173924 265348 173936
rect 265308 173896 265348 173924
rect 265308 173884 265314 173896
rect 265342 173884 265348 173896
rect 265400 173884 265406 173936
rect 270494 173884 270500 173936
rect 270552 173924 270558 173936
rect 270770 173924 270776 173936
rect 270552 173896 270776 173924
rect 270552 173884 270558 173896
rect 270770 173884 270776 173896
rect 270828 173884 270834 173936
rect 281718 173884 281724 173936
rect 281776 173924 281782 173936
rect 281902 173924 281908 173936
rect 281776 173896 281908 173924
rect 281776 173884 281782 173896
rect 281902 173884 281908 173896
rect 281960 173884 281966 173936
rect 284662 173884 284668 173936
rect 284720 173924 284726 173936
rect 284846 173924 284852 173936
rect 284720 173896 284852 173924
rect 284720 173884 284726 173896
rect 284846 173884 284852 173896
rect 284904 173884 284910 173936
rect 288710 173884 288716 173936
rect 288768 173924 288774 173936
rect 288894 173924 288900 173936
rect 288768 173896 288900 173924
rect 288768 173884 288774 173896
rect 288894 173884 288900 173896
rect 288952 173884 288958 173936
rect 323302 173884 323308 173936
rect 323360 173924 323366 173936
rect 323486 173924 323492 173936
rect 323360 173896 323492 173924
rect 323360 173884 323366 173896
rect 323486 173884 323492 173896
rect 323544 173884 323550 173936
rect 324590 173884 324596 173936
rect 324648 173924 324654 173936
rect 324682 173924 324688 173936
rect 324648 173896 324688 173924
rect 324648 173884 324654 173896
rect 324682 173884 324688 173896
rect 324740 173884 324746 173936
rect 325878 173884 325884 173936
rect 325936 173924 325942 173936
rect 325970 173924 325976 173936
rect 325936 173896 325976 173924
rect 325936 173884 325942 173896
rect 325970 173884 325976 173896
rect 326028 173884 326034 173936
rect 327166 173884 327172 173936
rect 327224 173924 327230 173936
rect 327258 173924 327264 173936
rect 327224 173896 327264 173924
rect 327224 173884 327230 173896
rect 327258 173884 327264 173896
rect 327316 173884 327322 173936
rect 357434 173884 357440 173936
rect 357492 173924 357498 173936
rect 357710 173924 357716 173936
rect 357492 173896 357716 173924
rect 357492 173884 357498 173896
rect 357710 173884 357716 173896
rect 357768 173884 357774 173936
rect 376938 173884 376944 173936
rect 376996 173924 377002 173936
rect 377030 173924 377036 173936
rect 376996 173896 377036 173924
rect 376996 173884 377002 173896
rect 377030 173884 377036 173896
rect 377088 173884 377094 173936
rect 463878 173884 463884 173936
rect 463936 173924 463942 173936
rect 464062 173924 464068 173936
rect 463936 173896 464068 173924
rect 463936 173884 463942 173896
rect 464062 173884 464068 173896
rect 464120 173884 464126 173936
rect 291654 173720 291660 173732
rect 291615 173692 291660 173720
rect 291654 173680 291660 173692
rect 291712 173680 291718 173732
rect 251174 172524 251180 172576
rect 251232 172564 251238 172576
rect 251542 172564 251548 172576
rect 251232 172536 251548 172564
rect 251232 172524 251238 172536
rect 251542 172524 251548 172536
rect 251600 172524 251606 172576
rect 273530 172564 273536 172576
rect 273491 172536 273536 172564
rect 273530 172524 273536 172536
rect 273588 172524 273594 172576
rect 289998 172564 290004 172576
rect 289959 172536 290004 172564
rect 289998 172524 290004 172536
rect 290056 172524 290062 172576
rect 331582 172524 331588 172576
rect 331640 172524 331646 172576
rect 337102 172524 337108 172576
rect 337160 172524 337166 172576
rect 329926 172456 329932 172508
rect 329984 172496 329990 172508
rect 330202 172496 330208 172508
rect 329984 172468 330208 172496
rect 329984 172456 329990 172468
rect 330202 172456 330208 172468
rect 330260 172456 330266 172508
rect 331600 172440 331628 172524
rect 337120 172440 337148 172524
rect 331582 172388 331588 172440
rect 331640 172388 331646 172440
rect 337102 172388 337108 172440
rect 337160 172388 337166 172440
rect 299750 171096 299756 171148
rect 299808 171136 299814 171148
rect 299845 171139 299903 171145
rect 299845 171136 299857 171139
rect 299808 171108 299857 171136
rect 299808 171096 299814 171108
rect 299845 171105 299857 171108
rect 299891 171105 299903 171139
rect 301038 171136 301044 171148
rect 300999 171108 301044 171136
rect 299845 171099 299903 171105
rect 301038 171096 301044 171108
rect 301096 171096 301102 171148
rect 306834 171136 306840 171148
rect 306795 171108 306840 171136
rect 306834 171096 306840 171108
rect 306892 171096 306898 171148
rect 244366 171028 244372 171080
rect 244424 171028 244430 171080
rect 247129 171071 247187 171077
rect 247129 171037 247141 171071
rect 247175 171068 247187 171071
rect 247218 171068 247224 171080
rect 247175 171040 247224 171068
rect 247175 171037 247187 171040
rect 247129 171031 247187 171037
rect 247218 171028 247224 171040
rect 247276 171028 247282 171080
rect 266630 171068 266636 171080
rect 266591 171040 266636 171068
rect 266630 171028 266636 171040
rect 266688 171028 266694 171080
rect 331582 171068 331588 171080
rect 331543 171040 331588 171068
rect 331582 171028 331588 171040
rect 331640 171028 331646 171080
rect 337102 171068 337108 171080
rect 337063 171040 337108 171068
rect 337102 171028 337108 171040
rect 337160 171028 337166 171080
rect 244384 171000 244412 171028
rect 244550 171000 244556 171012
rect 244384 170972 244556 171000
rect 244550 170960 244556 170972
rect 244608 170960 244614 171012
rect 267826 169776 267832 169788
rect 267787 169748 267832 169776
rect 267826 169736 267832 169748
rect 267884 169736 267890 169788
rect 278866 167056 278872 167068
rect 278792 167028 278872 167056
rect 278792 166932 278820 167028
rect 278866 167016 278872 167028
rect 278924 167016 278930 167068
rect 310790 167016 310796 167068
rect 310848 167016 310854 167068
rect 357526 167016 357532 167068
rect 357584 167056 357590 167068
rect 357710 167056 357716 167068
rect 357584 167028 357716 167056
rect 357584 167016 357590 167028
rect 357710 167016 357716 167028
rect 357768 167016 357774 167068
rect 431310 167016 431316 167068
rect 431368 167056 431374 167068
rect 431494 167056 431500 167068
rect 431368 167028 431500 167056
rect 431368 167016 431374 167028
rect 431494 167016 431500 167028
rect 431552 167016 431558 167068
rect 278774 166880 278780 166932
rect 278832 166880 278838 166932
rect 310808 166920 310836 167016
rect 310882 166920 310888 166932
rect 310808 166892 310888 166920
rect 310882 166880 310888 166892
rect 310940 166880 310946 166932
rect 341058 164908 341064 164960
rect 341116 164948 341122 164960
rect 341242 164948 341248 164960
rect 341116 164920 341248 164948
rect 341116 164908 341122 164920
rect 341242 164908 341248 164920
rect 341300 164908 341306 164960
rect 251266 164296 251272 164348
rect 251324 164296 251330 164348
rect 251174 164228 251180 164280
rect 251232 164228 251238 164280
rect 235074 164200 235080 164212
rect 235035 164172 235080 164200
rect 235074 164160 235080 164172
rect 235132 164160 235138 164212
rect 236270 164160 236276 164212
rect 236328 164200 236334 164212
rect 236454 164200 236460 164212
rect 236328 164172 236460 164200
rect 236328 164160 236334 164172
rect 236454 164160 236460 164172
rect 236512 164160 236518 164212
rect 251192 164132 251220 164228
rect 251284 164212 251312 164296
rect 285950 164228 285956 164280
rect 286008 164228 286014 164280
rect 251266 164160 251272 164212
rect 251324 164160 251330 164212
rect 270678 164160 270684 164212
rect 270736 164160 270742 164212
rect 251358 164132 251364 164144
rect 251192 164104 251364 164132
rect 251358 164092 251364 164104
rect 251416 164092 251422 164144
rect 270696 164132 270724 164160
rect 270770 164132 270776 164144
rect 270696 164104 270776 164132
rect 270770 164092 270776 164104
rect 270828 164092 270834 164144
rect 285968 164132 285996 164228
rect 340874 164160 340880 164212
rect 340932 164200 340938 164212
rect 341058 164200 341064 164212
rect 340932 164172 341064 164200
rect 340932 164160 340938 164172
rect 341058 164160 341064 164172
rect 341116 164160 341122 164212
rect 367002 164200 367008 164212
rect 366963 164172 367008 164200
rect 367002 164160 367008 164172
rect 367060 164160 367066 164212
rect 372522 164160 372528 164212
rect 372580 164200 372586 164212
rect 372798 164200 372804 164212
rect 372580 164172 372804 164200
rect 372580 164160 372586 164172
rect 372798 164160 372804 164172
rect 372856 164160 372862 164212
rect 375837 164203 375895 164209
rect 375837 164169 375849 164203
rect 375883 164200 375895 164203
rect 375926 164200 375932 164212
rect 375883 164172 375932 164200
rect 375883 164169 375895 164172
rect 375837 164163 375895 164169
rect 375926 164160 375932 164172
rect 375984 164160 375990 164212
rect 286134 164132 286140 164144
rect 285968 164104 286140 164132
rect 286134 164092 286140 164104
rect 286192 164092 286198 164144
rect 230658 162800 230664 162852
rect 230716 162840 230722 162852
rect 230750 162840 230756 162852
rect 230716 162812 230756 162840
rect 230716 162800 230722 162812
rect 230750 162800 230756 162812
rect 230808 162800 230814 162852
rect 250162 162800 250168 162852
rect 250220 162840 250226 162852
rect 250254 162840 250260 162852
rect 250220 162812 250260 162840
rect 250220 162800 250226 162812
rect 250254 162800 250260 162812
rect 250312 162800 250318 162852
rect 251358 162800 251364 162852
rect 251416 162840 251422 162852
rect 251634 162840 251640 162852
rect 251416 162812 251640 162840
rect 251416 162800 251422 162812
rect 251634 162800 251640 162812
rect 251692 162800 251698 162852
rect 393593 162843 393651 162849
rect 393593 162809 393605 162843
rect 393639 162840 393651 162843
rect 393682 162840 393688 162852
rect 393639 162812 393688 162840
rect 393639 162809 393651 162812
rect 393593 162803 393651 162809
rect 393682 162800 393688 162812
rect 393740 162800 393746 162852
rect 330110 162732 330116 162784
rect 330168 162772 330174 162784
rect 330205 162775 330263 162781
rect 330205 162772 330217 162775
rect 330168 162744 330217 162772
rect 330168 162732 330174 162744
rect 330205 162741 330217 162744
rect 330251 162741 330263 162775
rect 330205 162735 330263 162741
rect 247126 161480 247132 161492
rect 247087 161452 247132 161480
rect 247126 161440 247132 161452
rect 247184 161440 247190 161492
rect 265158 161440 265164 161492
rect 265216 161480 265222 161492
rect 265250 161480 265256 161492
rect 265216 161452 265256 161480
rect 265216 161440 265222 161452
rect 265250 161440 265256 161452
rect 265308 161440 265314 161492
rect 266633 161483 266691 161489
rect 266633 161449 266645 161483
rect 266679 161480 266691 161483
rect 266814 161480 266820 161492
rect 266679 161452 266820 161480
rect 266679 161449 266691 161452
rect 266633 161443 266691 161449
rect 266814 161440 266820 161452
rect 266872 161440 266878 161492
rect 294322 161440 294328 161492
rect 294380 161480 294386 161492
rect 294414 161480 294420 161492
rect 294380 161452 294420 161480
rect 294380 161440 294386 161452
rect 294414 161440 294420 161452
rect 294472 161440 294478 161492
rect 295610 161440 295616 161492
rect 295668 161480 295674 161492
rect 295702 161480 295708 161492
rect 295668 161452 295708 161480
rect 295668 161440 295674 161452
rect 295702 161440 295708 161452
rect 295760 161440 295766 161492
rect 296898 161440 296904 161492
rect 296956 161480 296962 161492
rect 296990 161480 296996 161492
rect 296956 161452 296996 161480
rect 296956 161440 296962 161452
rect 296990 161440 296996 161452
rect 297048 161440 297054 161492
rect 331585 161483 331643 161489
rect 331585 161449 331597 161483
rect 331631 161480 331643 161483
rect 331674 161480 331680 161492
rect 331631 161452 331680 161480
rect 331631 161449 331643 161452
rect 331585 161443 331643 161449
rect 331674 161440 331680 161452
rect 331732 161440 331738 161492
rect 337105 161483 337163 161489
rect 337105 161449 337117 161483
rect 337151 161480 337163 161483
rect 337286 161480 337292 161492
rect 337151 161452 337292 161480
rect 337151 161449 337163 161452
rect 337105 161443 337163 161449
rect 337286 161440 337292 161452
rect 337344 161440 337350 161492
rect 285953 161415 286011 161421
rect 285953 161381 285965 161415
rect 285999 161412 286011 161415
rect 286134 161412 286140 161424
rect 285999 161384 286140 161412
rect 285999 161381 286011 161384
rect 285953 161375 286011 161381
rect 286134 161372 286140 161384
rect 286192 161372 286198 161424
rect 265158 160012 265164 160064
rect 265216 160052 265222 160064
rect 265345 160055 265403 160061
rect 265345 160052 265357 160055
rect 265216 160024 265357 160052
rect 265216 160012 265222 160024
rect 265345 160021 265357 160024
rect 265391 160021 265403 160055
rect 265345 160015 265403 160021
rect 272150 160012 272156 160064
rect 272208 160052 272214 160064
rect 272337 160055 272395 160061
rect 272337 160052 272349 160055
rect 272208 160024 272349 160052
rect 272208 160012 272214 160024
rect 272337 160021 272349 160024
rect 272383 160021 272395 160055
rect 272337 160015 272395 160021
rect 378226 157700 378232 157752
rect 378284 157740 378290 157752
rect 386322 157740 386328 157752
rect 378284 157712 386328 157740
rect 378284 157700 378290 157712
rect 386322 157700 386328 157712
rect 386380 157700 386386 157752
rect 306374 157496 306380 157548
rect 306432 157536 306438 157548
rect 315942 157536 315948 157548
rect 306432 157508 315948 157536
rect 306432 157496 306438 157508
rect 315942 157496 315948 157508
rect 316000 157496 316006 157548
rect 336734 157496 336740 157548
rect 336792 157536 336798 157548
rect 346302 157536 346308 157548
rect 336792 157508 346308 157536
rect 336792 157496 336798 157508
rect 346302 157496 346308 157508
rect 346360 157496 346366 157548
rect 417878 157496 417884 157548
rect 417936 157536 417942 157548
rect 418154 157536 418160 157548
rect 417936 157508 418160 157536
rect 417936 157496 417942 157508
rect 418154 157496 418160 157508
rect 418212 157496 418218 157548
rect 437198 157496 437204 157548
rect 437256 157536 437262 157548
rect 437474 157536 437480 157548
rect 437256 157508 437480 157536
rect 437256 157496 437262 157508
rect 437474 157496 437480 157508
rect 437532 157496 437538 157548
rect 267734 157428 267740 157480
rect 267792 157428 267798 157480
rect 460198 157468 460204 157480
rect 460032 157440 460204 157468
rect 267752 157344 267780 157428
rect 357618 157360 357624 157412
rect 357676 157360 357682 157412
rect 267734 157292 267740 157344
rect 267792 157292 267798 157344
rect 325970 157224 325976 157276
rect 326028 157224 326034 157276
rect 357636 157264 357664 157360
rect 460032 157344 460060 157440
rect 460198 157428 460204 157440
rect 460256 157428 460262 157480
rect 460014 157292 460020 157344
rect 460072 157292 460078 157344
rect 357710 157264 357716 157276
rect 357636 157236 357716 157264
rect 357710 157224 357716 157236
rect 357768 157224 357774 157276
rect 325988 157140 326016 157224
rect 325970 157088 325976 157140
rect 326028 157088 326034 157140
rect 299750 156612 299756 156664
rect 299808 156652 299814 156664
rect 299934 156652 299940 156664
rect 299808 156624 299940 156652
rect 299808 156612 299814 156624
rect 299934 156612 299940 156624
rect 299992 156612 299998 156664
rect 245838 156544 245844 156596
rect 245896 156584 245902 156596
rect 246022 156584 246028 156596
rect 245896 156556 246028 156584
rect 245896 156544 245902 156556
rect 246022 156544 246028 156556
rect 246080 156544 246086 156596
rect 367002 154680 367008 154692
rect 366963 154652 367008 154680
rect 367002 154640 367008 154652
rect 367060 154640 367066 154692
rect 235074 154612 235080 154624
rect 235035 154584 235080 154612
rect 235074 154572 235080 154584
rect 235132 154572 235138 154624
rect 375834 154612 375840 154624
rect 375795 154584 375840 154612
rect 375834 154572 375840 154584
rect 375892 154572 375898 154624
rect 232317 154547 232375 154553
rect 232317 154513 232329 154547
rect 232363 154544 232375 154547
rect 232406 154544 232412 154556
rect 232363 154516 232412 154544
rect 232363 154513 232375 154516
rect 232317 154507 232375 154513
rect 232406 154504 232412 154516
rect 232464 154504 232470 154556
rect 259730 154544 259736 154556
rect 259691 154516 259736 154544
rect 259730 154504 259736 154516
rect 259788 154504 259794 154556
rect 366726 154504 366732 154556
rect 366784 154544 366790 154556
rect 367002 154544 367008 154556
rect 366784 154516 367008 154544
rect 366784 154504 366790 154516
rect 367002 154504 367008 154516
rect 367060 154504 367066 154556
rect 247126 153252 247132 153264
rect 247052 153224 247132 153252
rect 247052 153196 247080 153224
rect 247126 153212 247132 153224
rect 247184 153212 247190 153264
rect 337286 153252 337292 153264
rect 337212 153224 337292 153252
rect 337212 153196 337240 153224
rect 337286 153212 337292 153224
rect 337344 153212 337350 153264
rect 393590 153252 393596 153264
rect 393551 153224 393596 153252
rect 393590 153212 393596 153224
rect 393648 153212 393654 153264
rect 247034 153144 247040 153196
rect 247092 153144 247098 153196
rect 270770 153144 270776 153196
rect 270828 153184 270834 153196
rect 270862 153184 270868 153196
rect 270828 153156 270868 153184
rect 270828 153144 270834 153156
rect 270862 153144 270868 153156
rect 270920 153144 270926 153196
rect 273530 153184 273536 153196
rect 273491 153156 273536 153184
rect 273530 153144 273536 153156
rect 273588 153144 273594 153196
rect 289998 153144 290004 153196
rect 290056 153184 290062 153196
rect 290090 153184 290096 153196
rect 290056 153156 290096 153184
rect 290056 153144 290062 153156
rect 290090 153144 290096 153156
rect 290148 153144 290154 153196
rect 291470 153144 291476 153196
rect 291528 153184 291534 153196
rect 291562 153184 291568 153196
rect 291528 153156 291568 153184
rect 291528 153144 291534 153156
rect 291562 153144 291568 153156
rect 291620 153144 291626 153196
rect 294230 153144 294236 153196
rect 294288 153184 294294 153196
rect 294322 153184 294328 153196
rect 294288 153156 294328 153184
rect 294288 153144 294294 153156
rect 294322 153144 294328 153156
rect 294380 153144 294386 153196
rect 310790 153184 310796 153196
rect 310751 153156 310796 153184
rect 310790 153144 310796 153156
rect 310848 153144 310854 153196
rect 337194 153144 337200 153196
rect 337252 153144 337258 153196
rect 266814 151784 266820 151836
rect 266872 151784 266878 151836
rect 285950 151824 285956 151836
rect 285911 151796 285956 151824
rect 285950 151784 285956 151796
rect 286008 151784 286014 151836
rect 3326 151716 3332 151768
rect 3384 151756 3390 151768
rect 24118 151756 24124 151768
rect 3384 151728 24124 151756
rect 3384 151716 3390 151728
rect 24118 151716 24124 151728
rect 24176 151716 24182 151768
rect 266832 151700 266860 151784
rect 266814 151648 266820 151700
rect 266872 151648 266878 151700
rect 245746 150424 245752 150476
rect 245804 150464 245810 150476
rect 246114 150464 246120 150476
rect 245804 150436 246120 150464
rect 245804 150424 245810 150436
rect 246114 150424 246120 150436
rect 246172 150424 246178 150476
rect 265342 150464 265348 150476
rect 265303 150436 265348 150464
rect 265342 150424 265348 150436
rect 265400 150424 265406 150476
rect 296622 150356 296628 150408
rect 296680 150396 296686 150408
rect 296898 150396 296904 150408
rect 296680 150368 296904 150396
rect 296680 150356 296686 150368
rect 296898 150356 296904 150368
rect 296956 150356 296962 150408
rect 393590 148492 393596 148504
rect 393551 148464 393596 148492
rect 393590 148452 393596 148464
rect 393648 148452 393654 148504
rect 281718 148356 281724 148368
rect 281679 148328 281724 148356
rect 281718 148316 281724 148328
rect 281776 148316 281782 148368
rect 272334 148288 272340 148300
rect 272295 148260 272340 148288
rect 272334 148248 272340 148260
rect 272392 148248 272398 148300
rect 235074 147704 235080 147756
rect 235132 147704 235138 147756
rect 463697 147747 463755 147753
rect 463697 147713 463709 147747
rect 463743 147744 463755 147747
rect 463786 147744 463792 147756
rect 463743 147716 463792 147744
rect 463743 147713 463755 147716
rect 463697 147707 463755 147713
rect 463786 147704 463792 147716
rect 463844 147704 463850 147756
rect 235092 147620 235120 147704
rect 357526 147636 357532 147688
rect 357584 147676 357590 147688
rect 357710 147676 357716 147688
rect 357584 147648 357716 147676
rect 357584 147636 357590 147648
rect 357710 147636 357716 147648
rect 357768 147636 357774 147688
rect 235074 147568 235080 147620
rect 235132 147568 235138 147620
rect 259730 147608 259736 147620
rect 259691 147580 259736 147608
rect 259730 147568 259736 147580
rect 259788 147568 259794 147620
rect 310790 147608 310796 147620
rect 310751 147580 310796 147608
rect 310790 147568 310796 147580
rect 310848 147568 310854 147620
rect 331398 146044 331404 146056
rect 331359 146016 331404 146044
rect 331398 146004 331404 146016
rect 331456 146004 331462 146056
rect 232314 145024 232320 145036
rect 232275 144996 232320 145024
rect 232314 144984 232320 144996
rect 232372 144984 232378 145036
rect 330202 144956 330208 144968
rect 330163 144928 330208 144956
rect 330202 144916 330208 144928
rect 330260 144916 330266 144968
rect 463694 144916 463700 144968
rect 463752 144956 463758 144968
rect 463752 144928 463797 144956
rect 463752 144916 463758 144928
rect 267734 144848 267740 144900
rect 267792 144888 267798 144900
rect 267918 144888 267924 144900
rect 267792 144860 267924 144888
rect 267792 144848 267798 144860
rect 267918 144848 267924 144860
rect 267976 144848 267982 144900
rect 273530 144888 273536 144900
rect 273491 144860 273536 144888
rect 273530 144848 273536 144860
rect 273588 144848 273594 144900
rect 284662 144848 284668 144900
rect 284720 144888 284726 144900
rect 284754 144888 284760 144900
rect 284720 144860 284760 144888
rect 284720 144848 284726 144860
rect 284754 144848 284760 144860
rect 284812 144848 284818 144900
rect 323394 144848 323400 144900
rect 323452 144888 323458 144900
rect 323486 144888 323492 144900
rect 323452 144860 323492 144888
rect 323452 144848 323458 144860
rect 323486 144848 323492 144860
rect 323544 144848 323550 144900
rect 324590 144848 324596 144900
rect 324648 144888 324654 144900
rect 324774 144888 324780 144900
rect 324648 144860 324780 144888
rect 324648 144848 324654 144860
rect 324774 144848 324780 144860
rect 324832 144848 324838 144900
rect 325878 144848 325884 144900
rect 325936 144888 325942 144900
rect 326062 144888 326068 144900
rect 325936 144860 326068 144888
rect 325936 144848 325942 144860
rect 326062 144848 326068 144860
rect 326120 144848 326126 144900
rect 357618 144888 357624 144900
rect 357579 144860 357624 144888
rect 357618 144848 357624 144860
rect 357676 144848 357682 144900
rect 367002 144888 367008 144900
rect 366963 144860 367008 144888
rect 367002 144848 367008 144860
rect 367060 144848 367066 144900
rect 459922 144848 459928 144900
rect 459980 144888 459986 144900
rect 460198 144888 460204 144900
rect 459980 144860 460204 144888
rect 459980 144848 459986 144860
rect 460198 144848 460204 144860
rect 460256 144848 460262 144900
rect 251358 143624 251364 143676
rect 251416 143664 251422 143676
rect 251542 143664 251548 143676
rect 251416 143636 251548 143664
rect 251416 143624 251422 143636
rect 251542 143624 251548 143636
rect 251600 143624 251606 143676
rect 281718 143596 281724 143608
rect 281679 143568 281724 143596
rect 281718 143556 281724 143568
rect 281776 143556 281782 143608
rect 230842 143528 230848 143540
rect 230803 143500 230848 143528
rect 230842 143488 230848 143500
rect 230900 143488 230906 143540
rect 232314 143528 232320 143540
rect 232275 143500 232320 143528
rect 232314 143488 232320 143500
rect 232372 143488 232378 143540
rect 245838 143528 245844 143540
rect 245799 143500 245844 143528
rect 245838 143488 245844 143500
rect 245896 143488 245902 143540
rect 250162 143528 250168 143540
rect 250123 143500 250168 143528
rect 250162 143488 250168 143500
rect 250220 143488 250226 143540
rect 329926 143488 329932 143540
rect 329984 143528 329990 143540
rect 330202 143528 330208 143540
rect 329984 143500 330208 143528
rect 329984 143488 329990 143500
rect 330202 143488 330208 143500
rect 330260 143488 330266 143540
rect 393593 142171 393651 142177
rect 393593 142137 393605 142171
rect 393639 142168 393651 142171
rect 393682 142168 393688 142180
rect 393639 142140 393688 142168
rect 393639 142137 393651 142140
rect 393593 142131 393651 142137
rect 393682 142128 393688 142140
rect 393740 142128 393746 142180
rect 251358 142100 251364 142112
rect 251319 142072 251364 142100
rect 251358 142060 251364 142072
rect 251416 142060 251422 142112
rect 296806 140700 296812 140752
rect 296864 140740 296870 140752
rect 296990 140740 296996 140752
rect 296864 140712 296996 140740
rect 296864 140700 296870 140712
rect 296990 140700 296996 140712
rect 297048 140700 297054 140752
rect 324774 139924 324780 139936
rect 324735 139896 324780 139924
rect 324774 139884 324780 139896
rect 324832 139884 324838 139936
rect 296901 139383 296959 139389
rect 296901 139349 296913 139383
rect 296947 139380 296959 139383
rect 296990 139380 296996 139392
rect 296947 139352 296996 139380
rect 296947 139349 296959 139352
rect 296901 139343 296959 139349
rect 296990 139340 296996 139352
rect 297048 139340 297054 139392
rect 341242 138660 341248 138712
rect 341300 138700 341306 138712
rect 341337 138703 341395 138709
rect 341337 138700 341349 138703
rect 341300 138672 341349 138700
rect 341300 138660 341306 138672
rect 341337 138669 341349 138672
rect 341383 138669 341395 138703
rect 341337 138663 341395 138669
rect 302510 138524 302516 138576
rect 302568 138564 302574 138576
rect 302694 138564 302700 138576
rect 302568 138536 302700 138564
rect 302568 138524 302574 138536
rect 302694 138524 302700 138536
rect 302752 138524 302758 138576
rect 244366 138048 244372 138100
rect 244424 138048 244430 138100
rect 310882 138088 310888 138100
rect 310808 138060 310888 138088
rect 235074 137980 235080 138032
rect 235132 137980 235138 138032
rect 235092 137896 235120 137980
rect 244384 137964 244412 138048
rect 259638 137980 259644 138032
rect 259696 138020 259702 138032
rect 259822 138020 259828 138032
rect 259696 137992 259828 138020
rect 259696 137980 259702 137992
rect 259822 137980 259828 137992
rect 259880 137980 259886 138032
rect 310808 137964 310836 138060
rect 310882 138048 310888 138060
rect 310940 138048 310946 138100
rect 463694 137980 463700 138032
rect 463752 137980 463758 138032
rect 244366 137912 244372 137964
rect 244424 137912 244430 137964
rect 245838 137952 245844 137964
rect 245799 137924 245844 137952
rect 245838 137912 245844 137924
rect 245896 137912 245902 137964
rect 250162 137952 250168 137964
rect 250123 137924 250168 137952
rect 250162 137912 250168 137924
rect 250220 137912 250226 137964
rect 310790 137912 310796 137964
rect 310848 137912 310854 137964
rect 357618 137952 357624 137964
rect 357579 137924 357624 137952
rect 357618 137912 357624 137924
rect 357676 137912 357682 137964
rect 463712 137952 463740 137980
rect 463878 137952 463884 137964
rect 463712 137924 463884 137952
rect 463878 137912 463884 137924
rect 463936 137912 463942 137964
rect 235074 137844 235080 137896
rect 235132 137844 235138 137896
rect 285766 137708 285772 137760
rect 285824 137748 285830 137760
rect 286134 137748 286140 137760
rect 285824 137720 286140 137748
rect 285824 137708 285830 137720
rect 286134 137708 286140 137720
rect 286192 137708 286198 137760
rect 326062 137748 326068 137760
rect 326023 137720 326068 137748
rect 326062 137708 326068 137720
rect 326120 137708 326126 137760
rect 299750 137368 299756 137420
rect 299808 137408 299814 137420
rect 299934 137408 299940 137420
rect 299808 137380 299940 137408
rect 299808 137368 299814 137380
rect 299934 137368 299940 137380
rect 299992 137368 299998 137420
rect 2774 136484 2780 136536
rect 2832 136524 2838 136536
rect 5074 136524 5080 136536
rect 2832 136496 5080 136524
rect 2832 136484 2838 136496
rect 5074 136484 5080 136496
rect 5132 136484 5138 136536
rect 367002 135368 367008 135380
rect 366963 135340 367008 135368
rect 367002 135328 367008 135340
rect 367060 135328 367066 135380
rect 273530 135260 273536 135312
rect 273588 135300 273594 135312
rect 273622 135300 273628 135312
rect 273588 135272 273628 135300
rect 273588 135260 273594 135272
rect 273622 135260 273628 135272
rect 273680 135260 273686 135312
rect 337102 135192 337108 135244
rect 337160 135232 337166 135244
rect 337194 135232 337200 135244
rect 337160 135204 337200 135232
rect 337160 135192 337166 135204
rect 337194 135192 337200 135204
rect 337252 135192 337258 135244
rect 339770 135232 339776 135244
rect 339731 135204 339776 135232
rect 339770 135192 339776 135204
rect 339828 135192 339834 135244
rect 357526 135192 357532 135244
rect 357584 135232 357590 135244
rect 357710 135232 357716 135244
rect 357584 135204 357716 135232
rect 357584 135192 357590 135204
rect 357710 135192 357716 135204
rect 357768 135192 357774 135244
rect 367002 135232 367008 135244
rect 366963 135204 367008 135232
rect 367002 135192 367008 135204
rect 367060 135192 367066 135244
rect 378226 134172 378232 134224
rect 378284 134212 378290 134224
rect 386322 134212 386328 134224
rect 378284 134184 386328 134212
rect 378284 134172 378290 134184
rect 386322 134172 386328 134184
rect 386380 134172 386386 134224
rect 456518 134104 456524 134156
rect 456576 134144 456582 134156
rect 457438 134144 457444 134156
rect 456576 134116 457444 134144
rect 456576 134104 456582 134116
rect 457438 134104 457444 134116
rect 457496 134104 457502 134156
rect 309042 134036 309048 134088
rect 309100 134076 309106 134088
rect 315942 134076 315948 134088
rect 309100 134048 315948 134076
rect 309100 134036 309106 134048
rect 315942 134036 315948 134048
rect 316000 134036 316006 134088
rect 437198 134036 437204 134088
rect 437256 134076 437262 134088
rect 437566 134076 437572 134088
rect 437256 134048 437572 134076
rect 437256 134036 437262 134048
rect 437566 134036 437572 134048
rect 437624 134036 437630 134088
rect 475562 134036 475568 134088
rect 475620 134076 475626 134088
rect 482922 134076 482928 134088
rect 475620 134048 482928 134076
rect 475620 134036 475626 134048
rect 482922 134036 482928 134048
rect 482980 134036 482986 134088
rect 417878 133968 417884 134020
rect 417936 134008 417942 134020
rect 418154 134008 418160 134020
rect 417936 133980 418160 134008
rect 417936 133968 417942 133980
rect 418154 133968 418160 133980
rect 418212 133968 418218 134020
rect 230842 133940 230848 133952
rect 230803 133912 230848 133940
rect 230842 133900 230848 133912
rect 230900 133900 230906 133952
rect 232314 133940 232320 133952
rect 232275 133912 232320 133940
rect 232314 133900 232320 133912
rect 232372 133900 232378 133952
rect 324774 133940 324780 133952
rect 324735 133912 324780 133940
rect 324774 133900 324780 133912
rect 324832 133900 324838 133952
rect 326062 133940 326068 133952
rect 326023 133912 326068 133940
rect 326062 133900 326068 133912
rect 326120 133900 326126 133952
rect 331398 133940 331404 133952
rect 331359 133912 331404 133940
rect 331398 133900 331404 133912
rect 331456 133900 331462 133952
rect 270770 133832 270776 133884
rect 270828 133872 270834 133884
rect 271046 133872 271052 133884
rect 270828 133844 271052 133872
rect 270828 133832 270834 133844
rect 271046 133832 271052 133844
rect 271104 133832 271110 133884
rect 299750 133872 299756 133884
rect 299711 133844 299756 133872
rect 299750 133832 299756 133844
rect 299808 133832 299814 133884
rect 301038 133872 301044 133884
rect 300999 133844 301044 133872
rect 301038 133832 301044 133844
rect 301096 133832 301102 133884
rect 357526 133872 357532 133884
rect 357487 133844 357532 133872
rect 357526 133832 357532 133844
rect 357584 133832 357590 133884
rect 251361 132515 251419 132521
rect 251361 132481 251373 132515
rect 251407 132512 251419 132515
rect 251450 132512 251456 132524
rect 251407 132484 251456 132512
rect 251407 132481 251419 132484
rect 251361 132475 251419 132481
rect 251450 132472 251456 132484
rect 251508 132472 251514 132524
rect 289906 132472 289912 132524
rect 289964 132512 289970 132524
rect 290090 132512 290096 132524
rect 289964 132484 290096 132512
rect 289964 132472 289970 132484
rect 290090 132472 290096 132484
rect 290148 132472 290154 132524
rect 295518 132472 295524 132524
rect 295576 132512 295582 132524
rect 295610 132512 295616 132524
rect 295576 132484 295616 132512
rect 295576 132472 295582 132484
rect 295610 132472 295616 132484
rect 295668 132472 295674 132524
rect 259641 132447 259699 132453
rect 259641 132413 259653 132447
rect 259687 132444 259699 132447
rect 259730 132444 259736 132456
rect 259687 132416 259736 132444
rect 259687 132413 259699 132416
rect 259641 132407 259699 132413
rect 259730 132404 259736 132416
rect 259788 132404 259794 132456
rect 262585 132447 262643 132453
rect 262585 132413 262597 132447
rect 262631 132444 262643 132447
rect 262674 132444 262680 132456
rect 262631 132416 262680 132444
rect 262631 132413 262643 132416
rect 262585 132407 262643 132413
rect 262674 132404 262680 132416
rect 262732 132404 262738 132456
rect 245746 131112 245752 131164
rect 245804 131152 245810 131164
rect 245930 131152 245936 131164
rect 245804 131124 245936 131152
rect 245804 131112 245810 131124
rect 245930 131112 245936 131124
rect 245988 131112 245994 131164
rect 393590 131044 393596 131096
rect 393648 131084 393654 131096
rect 393774 131084 393780 131096
rect 393648 131056 393780 131084
rect 393648 131044 393654 131056
rect 393774 131044 393780 131056
rect 393832 131044 393838 131096
rect 375834 130364 375840 130416
rect 375892 130404 375898 130416
rect 376110 130404 376116 130416
rect 375892 130376 376116 130404
rect 375892 130364 375898 130376
rect 376110 130364 376116 130376
rect 376168 130364 376174 130416
rect 463878 130364 463884 130416
rect 463936 130404 463942 130416
rect 464062 130404 464068 130416
rect 463936 130376 464068 130404
rect 463936 130364 463942 130376
rect 464062 130364 464068 130376
rect 464120 130364 464126 130416
rect 291381 129931 291439 129937
rect 291381 129897 291393 129931
rect 291427 129928 291439 129931
rect 291562 129928 291568 129940
rect 291427 129900 291568 129928
rect 291427 129897 291439 129900
rect 291381 129891 291439 129897
rect 291562 129888 291568 129900
rect 291620 129888 291626 129940
rect 291381 129659 291439 129665
rect 291381 129625 291393 129659
rect 291427 129656 291439 129659
rect 291470 129656 291476 129668
rect 291427 129628 291476 129656
rect 291427 129625 291439 129628
rect 291381 129619 291439 129625
rect 291470 129616 291476 129628
rect 291528 129616 291534 129668
rect 306742 128324 306748 128376
rect 306800 128324 306806 128376
rect 306760 128296 306788 128324
rect 306834 128296 306840 128308
rect 306760 128268 306840 128296
rect 306834 128256 306840 128268
rect 306892 128256 306898 128308
rect 341334 128296 341340 128308
rect 341295 128268 341340 128296
rect 341334 128256 341340 128268
rect 341392 128256 341398 128308
rect 310790 125780 310796 125792
rect 310751 125752 310796 125780
rect 310790 125740 310796 125752
rect 310848 125740 310854 125792
rect 367002 125644 367008 125656
rect 366963 125616 367008 125644
rect 367002 125604 367008 125616
rect 367060 125604 367066 125656
rect 377122 125604 377128 125656
rect 377180 125644 377186 125656
rect 377214 125644 377220 125656
rect 377180 125616 377220 125644
rect 377180 125604 377186 125616
rect 377214 125604 377220 125616
rect 377272 125604 377278 125656
rect 235074 125576 235080 125588
rect 235035 125548 235080 125576
rect 235074 125536 235080 125548
rect 235132 125536 235138 125588
rect 236270 125536 236276 125588
rect 236328 125576 236334 125588
rect 236454 125576 236460 125588
rect 236328 125548 236460 125576
rect 236328 125536 236334 125548
rect 236454 125536 236460 125548
rect 236512 125536 236518 125588
rect 330110 125536 330116 125588
rect 330168 125576 330174 125588
rect 330294 125576 330300 125588
rect 330168 125548 330300 125576
rect 330168 125536 330174 125548
rect 330294 125536 330300 125548
rect 330352 125536 330358 125588
rect 331398 125536 331404 125588
rect 331456 125576 331462 125588
rect 331582 125576 331588 125588
rect 331456 125548 331588 125576
rect 331456 125536 331462 125548
rect 331582 125536 331588 125548
rect 331640 125536 331646 125588
rect 337102 125536 337108 125588
rect 337160 125576 337166 125588
rect 337286 125576 337292 125588
rect 337160 125548 337292 125576
rect 337160 125536 337166 125548
rect 337286 125536 337292 125548
rect 337344 125536 337350 125588
rect 375745 125579 375803 125585
rect 375745 125545 375757 125579
rect 375791 125576 375803 125579
rect 375834 125576 375840 125588
rect 375791 125548 375840 125576
rect 375791 125545 375803 125548
rect 375745 125539 375803 125545
rect 375834 125536 375840 125548
rect 375892 125536 375898 125588
rect 339678 124244 339684 124296
rect 339736 124284 339742 124296
rect 339773 124287 339831 124293
rect 339773 124284 339785 124287
rect 339736 124256 339785 124284
rect 339736 124244 339742 124256
rect 339773 124253 339785 124256
rect 339819 124253 339831 124287
rect 339773 124247 339831 124253
rect 289906 124176 289912 124228
rect 289964 124216 289970 124228
rect 289998 124216 290004 124228
rect 289964 124188 290004 124216
rect 289964 124176 289970 124188
rect 289998 124176 290004 124188
rect 290056 124176 290062 124228
rect 299753 124219 299811 124225
rect 299753 124185 299765 124219
rect 299799 124216 299811 124219
rect 299842 124216 299848 124228
rect 299799 124188 299848 124216
rect 299799 124185 299811 124188
rect 299753 124179 299811 124185
rect 299842 124176 299848 124188
rect 299900 124176 299906 124228
rect 301041 124219 301099 124225
rect 301041 124185 301053 124219
rect 301087 124216 301099 124219
rect 301130 124216 301136 124228
rect 301087 124188 301136 124216
rect 301087 124185 301099 124188
rect 301041 124179 301099 124185
rect 301130 124176 301136 124188
rect 301188 124176 301194 124228
rect 357529 124219 357587 124225
rect 357529 124185 357541 124219
rect 357575 124216 357587 124219
rect 357618 124216 357624 124228
rect 357575 124188 357624 124216
rect 357575 124185 357587 124188
rect 357529 124179 357587 124185
rect 357618 124176 357624 124188
rect 357676 124176 357682 124228
rect 232314 124148 232320 124160
rect 232275 124120 232320 124148
rect 232314 124108 232320 124120
rect 232372 124108 232378 124160
rect 247310 124148 247316 124160
rect 247271 124120 247316 124148
rect 247310 124108 247316 124120
rect 247368 124108 247374 124160
rect 377033 124151 377091 124157
rect 377033 124117 377045 124151
rect 377079 124148 377091 124151
rect 377122 124148 377128 124160
rect 377079 124120 377128 124148
rect 377079 124117 377091 124120
rect 377033 124111 377091 124117
rect 377122 124108 377128 124120
rect 377180 124108 377186 124160
rect 456518 123088 456524 123140
rect 456576 123128 456582 123140
rect 457438 123128 457444 123140
rect 456576 123100 457444 123128
rect 456576 123088 456582 123100
rect 457438 123088 457444 123100
rect 457496 123088 457502 123140
rect 306006 123020 306012 123072
rect 306064 123060 306070 123072
rect 314562 123060 314568 123072
rect 306064 123032 314568 123060
rect 306064 123020 306070 123032
rect 314562 123020 314568 123032
rect 314620 123020 314626 123072
rect 369670 123020 369676 123072
rect 369728 123060 369734 123072
rect 376662 123060 376668 123072
rect 369728 123032 376668 123060
rect 369728 123020 369734 123032
rect 376662 123020 376668 123032
rect 376720 123020 376726 123072
rect 417878 122952 417884 123004
rect 417936 122992 417942 123004
rect 419350 122992 419356 123004
rect 417936 122964 419356 122992
rect 417936 122952 417942 122964
rect 419350 122952 419356 122964
rect 419408 122952 419414 123004
rect 437198 122952 437204 123004
rect 437256 122992 437262 123004
rect 437474 122992 437480 123004
rect 437256 122964 437480 122992
rect 437256 122952 437262 122964
rect 437474 122952 437480 122964
rect 437532 122952 437538 123004
rect 259638 122856 259644 122868
rect 259599 122828 259644 122856
rect 259638 122816 259644 122828
rect 259696 122816 259702 122868
rect 262582 122856 262588 122868
rect 262543 122828 262588 122856
rect 262582 122816 262588 122828
rect 262640 122816 262646 122868
rect 251358 122788 251364 122800
rect 251319 122760 251364 122788
rect 251358 122748 251364 122760
rect 251416 122748 251422 122800
rect 270773 122791 270831 122797
rect 270773 122757 270785 122791
rect 270819 122788 270831 122791
rect 270862 122788 270868 122800
rect 270819 122760 270868 122788
rect 270819 122757 270831 122760
rect 270773 122751 270831 122757
rect 270862 122748 270868 122760
rect 270920 122748 270926 122800
rect 285950 122748 285956 122800
rect 286008 122788 286014 122800
rect 286042 122788 286048 122800
rect 286008 122760 286048 122788
rect 286008 122748 286014 122760
rect 286042 122748 286048 122760
rect 286100 122748 286106 122800
rect 288710 122748 288716 122800
rect 288768 122788 288774 122800
rect 288802 122788 288808 122800
rect 288768 122760 288808 122788
rect 288768 122748 288774 122760
rect 288802 122748 288808 122760
rect 288860 122748 288866 122800
rect 294414 122788 294420 122800
rect 294375 122760 294420 122788
rect 294414 122748 294420 122760
rect 294472 122748 294478 122800
rect 295702 122788 295708 122800
rect 295663 122760 295708 122788
rect 295702 122748 295708 122760
rect 295760 122748 295766 122800
rect 303890 122788 303896 122800
rect 303851 122760 303896 122788
rect 303890 122748 303896 122760
rect 303948 122748 303954 122800
rect 324590 122788 324596 122800
rect 324551 122760 324596 122788
rect 324590 122748 324596 122760
rect 324648 122748 324654 122800
rect 325878 122788 325884 122800
rect 325839 122760 325884 122788
rect 325878 122748 325884 122760
rect 325936 122748 325942 122800
rect 339770 122788 339776 122800
rect 339731 122760 339776 122788
rect 339770 122748 339776 122760
rect 339828 122748 339834 122800
rect 372798 122788 372804 122800
rect 372759 122760 372804 122788
rect 372798 122748 372804 122760
rect 372856 122748 372862 122800
rect 296901 122723 296959 122729
rect 296901 122689 296913 122723
rect 296947 122720 296959 122723
rect 296990 122720 296996 122732
rect 296947 122692 296996 122720
rect 296947 122689 296959 122692
rect 296901 122683 296959 122689
rect 296990 122680 296996 122692
rect 297048 122680 297054 122732
rect 2774 122272 2780 122324
rect 2832 122312 2838 122324
rect 4982 122312 4988 122324
rect 2832 122284 4988 122312
rect 2832 122272 2838 122284
rect 4982 122272 4988 122284
rect 5040 122272 5046 122324
rect 310790 121496 310796 121508
rect 310751 121468 310796 121496
rect 310790 121456 310796 121468
rect 310848 121456 310854 121508
rect 389358 121428 389364 121440
rect 389319 121400 389364 121428
rect 389358 121388 389364 121400
rect 389416 121388 389422 121440
rect 291470 120068 291476 120080
rect 291431 120040 291476 120068
rect 291470 120028 291476 120040
rect 291528 120028 291534 120080
rect 393590 120068 393596 120080
rect 393551 120040 393596 120068
rect 393590 120028 393596 120040
rect 393648 120028 393654 120080
rect 278866 118736 278872 118788
rect 278924 118736 278930 118788
rect 278884 118652 278912 118736
rect 341242 118668 341248 118720
rect 341300 118708 341306 118720
rect 341426 118708 341432 118720
rect 341300 118680 341432 118708
rect 341300 118668 341306 118680
rect 341426 118668 341432 118680
rect 341484 118668 341490 118720
rect 278866 118600 278872 118652
rect 278924 118600 278930 118652
rect 339770 118028 339776 118040
rect 339731 118000 339776 118028
rect 339770 117988 339776 118000
rect 339828 117988 339834 118040
rect 295705 116603 295763 116609
rect 295705 116569 295717 116603
rect 295751 116600 295763 116603
rect 295794 116600 295800 116612
rect 295751 116572 295800 116600
rect 295751 116569 295763 116572
rect 295705 116563 295763 116569
rect 295794 116560 295800 116572
rect 295852 116560 295858 116612
rect 235074 115988 235080 116000
rect 235035 115960 235080 115988
rect 235074 115948 235080 115960
rect 235132 115948 235138 116000
rect 245930 115988 245936 116000
rect 245891 115960 245936 115988
rect 245930 115948 245936 115960
rect 245988 115948 245994 116000
rect 375742 115988 375748 116000
rect 375703 115960 375748 115988
rect 375742 115948 375748 115960
rect 375800 115948 375806 116000
rect 341153 115923 341211 115929
rect 341153 115889 341165 115923
rect 341199 115920 341211 115923
rect 341242 115920 341248 115932
rect 341199 115892 341248 115920
rect 341199 115889 341211 115892
rect 341153 115883 341211 115889
rect 341242 115880 341248 115892
rect 341300 115880 341306 115932
rect 366726 115880 366732 115932
rect 366784 115920 366790 115932
rect 367002 115920 367008 115932
rect 366784 115892 367008 115920
rect 366784 115880 366790 115892
rect 367002 115880 367008 115892
rect 367060 115880 367066 115932
rect 232314 114560 232320 114572
rect 232275 114532 232320 114560
rect 232314 114520 232320 114532
rect 232372 114520 232378 114572
rect 244274 114520 244280 114572
rect 244332 114560 244338 114572
rect 244458 114560 244464 114572
rect 244332 114532 244464 114560
rect 244332 114520 244338 114532
rect 244458 114520 244464 114532
rect 244516 114520 244522 114572
rect 245930 114560 245936 114572
rect 245891 114532 245936 114560
rect 245930 114520 245936 114532
rect 245988 114520 245994 114572
rect 247126 114520 247132 114572
rect 247184 114560 247190 114572
rect 247313 114563 247371 114569
rect 247313 114560 247325 114563
rect 247184 114532 247325 114560
rect 247184 114520 247190 114532
rect 247313 114529 247325 114532
rect 247359 114529 247371 114563
rect 247313 114523 247371 114529
rect 265158 114520 265164 114572
rect 265216 114560 265222 114572
rect 265250 114560 265256 114572
rect 265216 114532 265256 114560
rect 265216 114520 265222 114532
rect 265250 114520 265256 114532
rect 265308 114520 265314 114572
rect 377030 114560 377036 114572
rect 376991 114532 377036 114560
rect 377030 114520 377036 114532
rect 377088 114520 377094 114572
rect 272242 114452 272248 114504
rect 272300 114492 272306 114504
rect 272334 114492 272340 114504
rect 272300 114464 272340 114492
rect 272300 114452 272306 114464
rect 272334 114452 272340 114464
rect 272392 114452 272398 114504
rect 337013 114495 337071 114501
rect 337013 114461 337025 114495
rect 337059 114492 337071 114495
rect 337194 114492 337200 114504
rect 337059 114464 337200 114492
rect 337059 114461 337071 114464
rect 337013 114455 337071 114461
rect 337194 114452 337200 114464
rect 337252 114452 337258 114504
rect 463881 114495 463939 114501
rect 463881 114461 463893 114495
rect 463927 114492 463939 114495
rect 463970 114492 463976 114504
rect 463927 114464 463976 114492
rect 463927 114461 463939 114464
rect 463881 114455 463939 114461
rect 463970 114452 463976 114464
rect 464028 114452 464034 114504
rect 325881 114427 325939 114433
rect 325881 114393 325893 114427
rect 325927 114424 325939 114427
rect 326062 114424 326068 114436
rect 325927 114396 326068 114424
rect 325927 114393 325939 114396
rect 325881 114387 325939 114393
rect 326062 114384 326068 114396
rect 326120 114384 326126 114436
rect 301130 113268 301136 113280
rect 301056 113240 301136 113268
rect 301056 113212 301084 113240
rect 301130 113228 301136 113240
rect 301188 113228 301194 113280
rect 251361 113203 251419 113209
rect 251361 113169 251373 113203
rect 251407 113200 251419 113203
rect 251450 113200 251456 113212
rect 251407 113172 251456 113200
rect 251407 113169 251419 113172
rect 251361 113163 251419 113169
rect 251450 113160 251456 113172
rect 251508 113160 251514 113212
rect 259730 113160 259736 113212
rect 259788 113200 259794 113212
rect 259914 113200 259920 113212
rect 259788 113172 259920 113200
rect 259788 113160 259794 113172
rect 259914 113160 259920 113172
rect 259972 113160 259978 113212
rect 270770 113200 270776 113212
rect 270731 113172 270776 113200
rect 270770 113160 270776 113172
rect 270828 113160 270834 113212
rect 294414 113200 294420 113212
rect 294375 113172 294420 113200
rect 294414 113160 294420 113172
rect 294472 113160 294478 113212
rect 301038 113160 301044 113212
rect 301096 113160 301102 113212
rect 303890 113200 303896 113212
rect 303851 113172 303896 113200
rect 303890 113160 303896 113172
rect 303948 113160 303954 113212
rect 324590 113200 324596 113212
rect 324551 113172 324596 113200
rect 324590 113160 324596 113172
rect 324648 113160 324654 113212
rect 372798 113200 372804 113212
rect 372759 113172 372804 113200
rect 372798 113160 372804 113172
rect 372856 113160 372862 113212
rect 244274 113092 244280 113144
rect 244332 113132 244338 113144
rect 244369 113135 244427 113141
rect 244369 113132 244381 113135
rect 244332 113104 244381 113132
rect 244332 113092 244338 113104
rect 244369 113101 244381 113104
rect 244415 113101 244427 113135
rect 285950 113132 285956 113144
rect 285911 113104 285956 113132
rect 244369 113095 244427 113101
rect 285950 113092 285956 113104
rect 286008 113092 286014 113144
rect 296990 112820 296996 112872
rect 297048 112820 297054 112872
rect 297008 112736 297036 112820
rect 296990 112684 296996 112736
rect 297048 112684 297054 112736
rect 310790 111800 310796 111852
rect 310848 111840 310854 111852
rect 310974 111840 310980 111852
rect 310848 111812 310980 111840
rect 310848 111800 310854 111812
rect 310974 111800 310980 111812
rect 311032 111800 311038 111852
rect 290001 111775 290059 111781
rect 290001 111741 290013 111775
rect 290047 111772 290059 111775
rect 290090 111772 290096 111784
rect 290047 111744 290096 111772
rect 290047 111741 290059 111744
rect 290001 111735 290059 111741
rect 290090 111732 290096 111744
rect 290148 111732 290154 111784
rect 295702 111772 295708 111784
rect 295663 111744 295708 111772
rect 295702 111732 295708 111744
rect 295760 111732 295766 111784
rect 306282 110780 306288 110832
rect 306340 110820 306346 110832
rect 315942 110820 315948 110832
rect 306340 110792 315948 110820
rect 306340 110780 306346 110792
rect 315942 110780 315948 110792
rect 316000 110780 316006 110832
rect 248414 110712 248420 110764
rect 248472 110752 248478 110764
rect 254118 110752 254124 110764
rect 248472 110724 254124 110752
rect 248472 110712 248478 110724
rect 254118 110712 254124 110724
rect 254176 110712 254182 110764
rect 456518 110712 456524 110764
rect 456576 110752 456582 110764
rect 457438 110752 457444 110764
rect 456576 110724 457444 110752
rect 456576 110712 456582 110724
rect 457438 110712 457444 110724
rect 457496 110712 457502 110764
rect 259362 110576 259368 110628
rect 259420 110616 259426 110628
rect 267642 110616 267648 110628
rect 259420 110588 267648 110616
rect 259420 110576 259426 110588
rect 267642 110576 267648 110588
rect 267700 110576 267706 110628
rect 417878 110576 417884 110628
rect 417936 110616 417942 110628
rect 418154 110616 418160 110628
rect 417936 110588 418160 110616
rect 417936 110576 417942 110588
rect 418154 110576 418160 110588
rect 418212 110576 418218 110628
rect 437198 110576 437204 110628
rect 437256 110616 437262 110628
rect 437474 110616 437480 110628
rect 437256 110588 437480 110616
rect 437256 110576 437262 110588
rect 437474 110576 437480 110588
rect 437532 110576 437538 110628
rect 291470 110480 291476 110492
rect 291431 110452 291476 110480
rect 291470 110440 291476 110452
rect 291528 110440 291534 110492
rect 393590 110480 393596 110492
rect 393551 110452 393596 110480
rect 393590 110440 393596 110452
rect 393648 110440 393654 110492
rect 262493 109735 262551 109741
rect 262493 109701 262505 109735
rect 262539 109732 262551 109735
rect 262582 109732 262588 109744
rect 262539 109704 262588 109732
rect 262539 109701 262551 109704
rect 262493 109695 262551 109701
rect 262582 109692 262588 109704
rect 262640 109692 262646 109744
rect 357621 109735 357679 109741
rect 357621 109701 357633 109735
rect 357667 109732 357679 109735
rect 357710 109732 357716 109744
rect 357667 109704 357716 109732
rect 357667 109701 357679 109704
rect 357621 109695 357679 109701
rect 357710 109692 357716 109704
rect 357768 109692 357774 109744
rect 265158 109012 265164 109064
rect 265216 109012 265222 109064
rect 375742 109012 375748 109064
rect 375800 109012 375806 109064
rect 377030 109012 377036 109064
rect 377088 109012 377094 109064
rect 265176 108984 265204 109012
rect 265250 108984 265256 108996
rect 265176 108956 265256 108984
rect 265250 108944 265256 108956
rect 265308 108944 265314 108996
rect 375760 108984 375788 109012
rect 375834 108984 375840 108996
rect 375760 108956 375840 108984
rect 375834 108944 375840 108956
rect 375892 108944 375898 108996
rect 377048 108984 377076 109012
rect 377122 108984 377128 108996
rect 377048 108956 377128 108984
rect 377122 108944 377128 108956
rect 377180 108944 377186 108996
rect 323394 108032 323400 108044
rect 323355 108004 323400 108032
rect 323394 107992 323400 108004
rect 323452 107992 323458 108044
rect 247126 106292 247132 106344
rect 247184 106292 247190 106344
rect 341150 106332 341156 106344
rect 341111 106304 341156 106332
rect 341150 106292 341156 106304
rect 341208 106292 341214 106344
rect 235074 106264 235080 106276
rect 235035 106236 235080 106264
rect 235074 106224 235080 106236
rect 235132 106224 235138 106276
rect 236270 106224 236276 106276
rect 236328 106264 236334 106276
rect 236454 106264 236460 106276
rect 236328 106236 236460 106264
rect 236328 106224 236334 106236
rect 236454 106224 236460 106236
rect 236512 106224 236518 106276
rect 245930 106264 245936 106276
rect 245891 106236 245936 106264
rect 245930 106224 245936 106236
rect 245988 106224 245994 106276
rect 247144 106208 247172 106292
rect 284754 106224 284760 106276
rect 284812 106264 284818 106276
rect 284846 106264 284852 106276
rect 284812 106236 284852 106264
rect 284812 106224 284818 106236
rect 284846 106224 284852 106236
rect 284904 106224 284910 106276
rect 367002 106264 367008 106276
rect 366963 106236 367008 106264
rect 367002 106224 367008 106236
rect 367060 106224 367066 106276
rect 459922 106224 459928 106276
rect 459980 106264 459986 106276
rect 460106 106264 460112 106276
rect 459980 106236 460112 106264
rect 459980 106224 459986 106236
rect 460106 106224 460112 106236
rect 460164 106224 460170 106276
rect 247126 106156 247132 106208
rect 247184 106156 247190 106208
rect 262490 104904 262496 104916
rect 262451 104876 262496 104904
rect 262490 104864 262496 104876
rect 262548 104864 262554 104916
rect 267734 104864 267740 104916
rect 267792 104904 267798 104916
rect 267826 104904 267832 104916
rect 267792 104876 267832 104904
rect 267792 104864 267798 104876
rect 267826 104864 267832 104876
rect 267884 104864 267890 104916
rect 270678 104864 270684 104916
rect 270736 104904 270742 104916
rect 270770 104904 270776 104916
rect 270736 104876 270776 104904
rect 270736 104864 270742 104876
rect 270770 104864 270776 104876
rect 270828 104864 270834 104916
rect 299658 104864 299664 104916
rect 299716 104904 299722 104916
rect 299750 104904 299756 104916
rect 299716 104876 299756 104904
rect 299716 104864 299722 104876
rect 299750 104864 299756 104876
rect 299808 104864 299814 104916
rect 325970 104864 325976 104916
rect 326028 104904 326034 104916
rect 326062 104904 326068 104916
rect 326028 104876 326068 104904
rect 326028 104864 326034 104876
rect 326062 104864 326068 104876
rect 326120 104864 326126 104916
rect 337010 104904 337016 104916
rect 336971 104876 337016 104904
rect 337010 104864 337016 104876
rect 337068 104864 337074 104916
rect 393590 104864 393596 104916
rect 393648 104864 393654 104916
rect 463878 104904 463884 104916
rect 463839 104876 463884 104904
rect 463878 104864 463884 104876
rect 463936 104864 463942 104916
rect 232314 104836 232320 104848
rect 232275 104808 232320 104836
rect 232314 104796 232320 104808
rect 232372 104796 232378 104848
rect 324590 104836 324596 104848
rect 324551 104808 324596 104836
rect 324590 104796 324596 104808
rect 324648 104796 324654 104848
rect 337010 104728 337016 104780
rect 337068 104768 337074 104780
rect 337197 104771 337255 104777
rect 337197 104768 337209 104771
rect 337068 104740 337209 104768
rect 337068 104728 337074 104740
rect 337197 104737 337209 104740
rect 337243 104737 337255 104771
rect 393608 104768 393636 104864
rect 393682 104768 393688 104780
rect 393608 104740 393688 104768
rect 337197 104731 337255 104737
rect 393682 104728 393688 104740
rect 393740 104728 393746 104780
rect 289998 104224 290004 104236
rect 289959 104196 290004 104224
rect 289998 104184 290004 104196
rect 290056 104184 290062 104236
rect 244366 103544 244372 103556
rect 244327 103516 244372 103544
rect 244366 103504 244372 103516
rect 244424 103504 244430 103556
rect 285953 103547 286011 103553
rect 285953 103513 285965 103547
rect 285999 103544 286011 103547
rect 286042 103544 286048 103556
rect 285999 103516 286048 103544
rect 285999 103513 286011 103516
rect 285953 103507 286011 103513
rect 286042 103504 286048 103516
rect 286100 103504 286106 103556
rect 291470 103504 291476 103556
rect 291528 103504 291534 103556
rect 294414 103504 294420 103556
rect 294472 103504 294478 103556
rect 296898 103504 296904 103556
rect 296956 103544 296962 103556
rect 296990 103544 296996 103556
rect 296956 103516 296996 103544
rect 296956 103504 296962 103516
rect 296990 103504 296996 103516
rect 297048 103504 297054 103556
rect 389358 103544 389364 103556
rect 389319 103516 389364 103544
rect 389358 103504 389364 103516
rect 389416 103504 389422 103556
rect 247126 103476 247132 103488
rect 247087 103448 247132 103476
rect 247126 103436 247132 103448
rect 247184 103436 247190 103488
rect 291488 103476 291516 103504
rect 291654 103476 291660 103488
rect 291488 103448 291660 103476
rect 291654 103436 291660 103448
rect 291712 103436 291718 103488
rect 294432 103476 294460 103504
rect 294598 103476 294604 103488
rect 294432 103448 294604 103476
rect 294598 103436 294604 103448
rect 294656 103436 294662 103488
rect 327166 103476 327172 103488
rect 327127 103448 327172 103476
rect 327166 103436 327172 103448
rect 327224 103436 327230 103488
rect 331398 103476 331404 103488
rect 331359 103448 331404 103476
rect 331398 103436 331404 103448
rect 331456 103436 331462 103488
rect 372798 103436 372804 103488
rect 372856 103436 372862 103488
rect 244366 103368 244372 103420
rect 244424 103408 244430 103420
rect 244550 103408 244556 103420
rect 244424 103380 244556 103408
rect 244424 103368 244430 103380
rect 244550 103368 244556 103380
rect 244608 103368 244614 103420
rect 317690 103408 317696 103420
rect 317651 103380 317696 103408
rect 317690 103368 317696 103380
rect 317748 103368 317754 103420
rect 330110 103408 330116 103420
rect 330071 103380 330116 103408
rect 330110 103368 330116 103380
rect 330168 103368 330174 103420
rect 372709 103411 372767 103417
rect 372709 103377 372721 103411
rect 372755 103408 372767 103411
rect 372816 103408 372844 103436
rect 372755 103380 372844 103408
rect 372755 103377 372767 103380
rect 372709 103371 372767 103377
rect 310974 102252 310980 102264
rect 310900 102224 310980 102252
rect 310900 102196 310928 102224
rect 310974 102212 310980 102224
rect 311032 102212 311038 102264
rect 295705 102187 295763 102193
rect 295705 102153 295717 102187
rect 295751 102184 295763 102187
rect 295886 102184 295892 102196
rect 295751 102156 295892 102184
rect 295751 102153 295763 102156
rect 295705 102147 295763 102153
rect 295886 102144 295892 102156
rect 295944 102144 295950 102196
rect 310882 102144 310888 102196
rect 310940 102144 310946 102196
rect 393593 100691 393651 100697
rect 393593 100657 393605 100691
rect 393639 100688 393651 100691
rect 393682 100688 393688 100700
rect 393639 100660 393688 100688
rect 393639 100657 393651 100660
rect 393593 100651 393651 100657
rect 393682 100648 393688 100660
rect 393740 100648 393746 100700
rect 267826 99464 267832 99476
rect 267752 99436 267832 99464
rect 267752 99340 267780 99436
rect 267826 99424 267832 99436
rect 267884 99424 267890 99476
rect 377122 99424 377128 99476
rect 377180 99424 377186 99476
rect 341150 99356 341156 99408
rect 341208 99356 341214 99408
rect 267734 99288 267740 99340
rect 267792 99288 267798 99340
rect 341168 99328 341196 99356
rect 377140 99340 377168 99424
rect 341242 99328 341248 99340
rect 341168 99300 341248 99328
rect 341242 99288 341248 99300
rect 341300 99288 341306 99340
rect 357618 99328 357624 99340
rect 357579 99300 357624 99328
rect 357618 99288 357624 99300
rect 357676 99288 357682 99340
rect 377122 99288 377128 99340
rect 377180 99288 377186 99340
rect 310793 98719 310851 98725
rect 310793 98685 310805 98719
rect 310839 98716 310851 98719
rect 310882 98716 310888 98728
rect 310839 98688 310888 98716
rect 310839 98685 310851 98688
rect 310793 98679 310851 98685
rect 310882 98676 310888 98688
rect 310940 98676 310946 98728
rect 330113 98719 330171 98725
rect 330113 98685 330125 98719
rect 330159 98716 330171 98719
rect 330202 98716 330208 98728
rect 330159 98688 330208 98716
rect 330159 98685 330171 98688
rect 330113 98679 330171 98685
rect 330202 98676 330208 98688
rect 330260 98676 330266 98728
rect 389269 98719 389327 98725
rect 389269 98685 389281 98719
rect 389315 98716 389327 98719
rect 389358 98716 389364 98728
rect 389315 98688 389364 98716
rect 389315 98685 389327 98688
rect 389269 98679 389327 98685
rect 389358 98676 389364 98688
rect 389416 98676 389422 98728
rect 289998 97968 290004 97980
rect 289959 97940 290004 97968
rect 289998 97928 290004 97940
rect 290056 97928 290062 97980
rect 367002 96744 367008 96756
rect 366963 96716 367008 96744
rect 367002 96704 367008 96716
rect 367060 96704 367066 96756
rect 235074 96676 235080 96688
rect 235035 96648 235080 96676
rect 235074 96636 235080 96648
rect 235132 96636 235138 96688
rect 245930 96676 245936 96688
rect 245891 96648 245936 96676
rect 245930 96636 245936 96648
rect 245988 96636 245994 96688
rect 284846 96676 284852 96688
rect 284772 96648 284852 96676
rect 284772 96620 284800 96648
rect 284846 96636 284852 96648
rect 284904 96636 284910 96688
rect 284754 96568 284760 96620
rect 284812 96568 284818 96620
rect 327166 96608 327172 96620
rect 327127 96580 327172 96608
rect 327166 96568 327172 96580
rect 327224 96568 327230 96620
rect 265250 95316 265256 95328
rect 265211 95288 265256 95316
rect 265250 95276 265256 95288
rect 265308 95276 265314 95328
rect 272334 95276 272340 95328
rect 272392 95276 272398 95328
rect 299750 95276 299756 95328
rect 299808 95316 299814 95328
rect 299808 95288 299888 95316
rect 299808 95276 299814 95288
rect 232314 95248 232320 95260
rect 232275 95220 232320 95248
rect 232314 95208 232320 95220
rect 232372 95208 232378 95260
rect 262490 95208 262496 95260
rect 262548 95248 262554 95260
rect 262582 95248 262588 95260
rect 262548 95220 262588 95248
rect 262548 95208 262554 95220
rect 262582 95208 262588 95220
rect 262640 95208 262646 95260
rect 270678 95208 270684 95260
rect 270736 95248 270742 95260
rect 270770 95248 270776 95260
rect 270736 95220 270776 95248
rect 270736 95208 270742 95220
rect 270770 95208 270776 95220
rect 270828 95208 270834 95260
rect 272242 95208 272248 95260
rect 272300 95248 272306 95260
rect 272352 95248 272380 95276
rect 299860 95260 299888 95288
rect 272300 95220 272380 95248
rect 272300 95208 272306 95220
rect 299842 95208 299848 95260
rect 299900 95208 299906 95260
rect 317693 95251 317751 95257
rect 317693 95217 317705 95251
rect 317739 95248 317751 95251
rect 317782 95248 317788 95260
rect 317739 95220 317788 95248
rect 317739 95217 317751 95220
rect 317693 95211 317751 95217
rect 317782 95208 317788 95220
rect 317840 95208 317846 95260
rect 323394 95248 323400 95260
rect 323355 95220 323400 95248
rect 323394 95208 323400 95220
rect 323452 95208 323458 95260
rect 324590 95248 324596 95260
rect 324551 95220 324596 95248
rect 324590 95208 324596 95220
rect 324648 95208 324654 95260
rect 337194 95248 337200 95260
rect 337155 95220 337200 95248
rect 337194 95208 337200 95220
rect 337252 95208 337258 95260
rect 463694 95208 463700 95260
rect 463752 95248 463758 95260
rect 463878 95248 463884 95260
rect 463752 95220 463884 95248
rect 463752 95208 463758 95220
rect 463878 95208 463884 95220
rect 463936 95208 463942 95260
rect 259638 95140 259644 95192
rect 259696 95180 259702 95192
rect 259733 95183 259791 95189
rect 259733 95180 259745 95183
rect 259696 95152 259745 95180
rect 259696 95140 259702 95152
rect 259733 95149 259745 95152
rect 259779 95149 259791 95183
rect 259733 95143 259791 95149
rect 296898 95140 296904 95192
rect 296956 95180 296962 95192
rect 296990 95180 296996 95192
rect 296956 95152 296996 95180
rect 296956 95140 296962 95152
rect 296990 95140 296996 95152
rect 297048 95140 297054 95192
rect 463694 94160 463700 94172
rect 463655 94132 463700 94160
rect 463694 94120 463700 94132
rect 463752 94120 463758 94172
rect 247129 93891 247187 93897
rect 247129 93857 247141 93891
rect 247175 93888 247187 93891
rect 247218 93888 247224 93900
rect 247175 93860 247224 93888
rect 247175 93857 247187 93860
rect 247129 93851 247187 93857
rect 247218 93848 247224 93860
rect 247276 93848 247282 93900
rect 331398 93888 331404 93900
rect 331359 93860 331404 93888
rect 331398 93848 331404 93860
rect 331456 93848 331462 93900
rect 262582 93820 262588 93832
rect 262543 93792 262588 93820
rect 262582 93780 262588 93792
rect 262640 93780 262646 93832
rect 289998 93820 290004 93832
rect 289959 93792 290004 93820
rect 289998 93780 290004 93792
rect 290056 93780 290062 93832
rect 329929 93823 329987 93829
rect 329929 93789 329941 93823
rect 329975 93820 329987 93823
rect 330110 93820 330116 93832
rect 329975 93792 330116 93820
rect 329975 93789 329987 93792
rect 329929 93783 329987 93789
rect 330110 93780 330116 93792
rect 330168 93780 330174 93832
rect 245746 92488 245752 92540
rect 245804 92528 245810 92540
rect 245838 92528 245844 92540
rect 245804 92500 245844 92528
rect 245804 92488 245810 92500
rect 245838 92488 245844 92500
rect 245896 92488 245902 92540
rect 265250 92528 265256 92540
rect 265211 92500 265256 92528
rect 265250 92488 265256 92500
rect 265308 92488 265314 92540
rect 270681 90423 270739 90429
rect 270681 90389 270693 90423
rect 270727 90420 270739 90423
rect 270770 90420 270776 90432
rect 270727 90392 270776 90420
rect 270727 90389 270739 90392
rect 270681 90383 270739 90389
rect 270770 90380 270776 90392
rect 270828 90380 270834 90432
rect 272153 90423 272211 90429
rect 272153 90389 272165 90423
rect 272199 90420 272211 90423
rect 272242 90420 272248 90432
rect 272199 90392 272248 90420
rect 272199 90389 272211 90392
rect 272153 90383 272211 90389
rect 272242 90380 272248 90392
rect 272300 90380 272306 90432
rect 317782 89700 317788 89752
rect 317840 89700 317846 89752
rect 357526 89700 357532 89752
rect 357584 89740 357590 89752
rect 357710 89740 357716 89752
rect 357584 89712 357716 89740
rect 357584 89700 357590 89712
rect 357710 89700 357716 89712
rect 357768 89700 357774 89752
rect 431310 89700 431316 89752
rect 431368 89740 431374 89752
rect 431494 89740 431500 89752
rect 431368 89712 431500 89740
rect 431368 89700 431374 89712
rect 431494 89700 431500 89712
rect 431552 89700 431558 89752
rect 310790 89672 310796 89684
rect 310751 89644 310796 89672
rect 310790 89632 310796 89644
rect 310848 89632 310854 89684
rect 317800 89604 317828 89700
rect 389266 89672 389272 89684
rect 389227 89644 389272 89672
rect 389266 89632 389272 89644
rect 389324 89632 389330 89684
rect 317874 89604 317880 89616
rect 317800 89576 317880 89604
rect 317874 89564 317880 89576
rect 317932 89564 317938 89616
rect 281718 88952 281724 89004
rect 281776 88992 281782 89004
rect 281813 88995 281871 89001
rect 281813 88992 281825 88995
rect 281776 88964 281825 88992
rect 281776 88952 281782 88964
rect 281813 88961 281825 88964
rect 281859 88961 281871 88995
rect 281813 88955 281871 88961
rect 366910 87224 366916 87236
rect 366871 87196 366916 87224
rect 366910 87184 366916 87196
rect 366968 87184 366974 87236
rect 417878 87116 417884 87168
rect 417936 87156 417942 87168
rect 418614 87156 418620 87168
rect 417936 87128 418620 87156
rect 417936 87116 417942 87128
rect 418614 87116 418620 87128
rect 418672 87116 418678 87168
rect 454034 87116 454040 87168
rect 454092 87156 454098 87168
rect 463418 87156 463424 87168
rect 454092 87128 463424 87156
rect 454092 87116 454098 87128
rect 463418 87116 463424 87128
rect 463476 87116 463482 87168
rect 463694 87116 463700 87168
rect 463752 87156 463758 87168
rect 467926 87156 467932 87168
rect 463752 87128 467932 87156
rect 463752 87116 463758 87128
rect 467926 87116 467932 87128
rect 467984 87116 467990 87168
rect 494606 87116 494612 87168
rect 494664 87156 494670 87168
rect 502242 87156 502248 87168
rect 494664 87128 502248 87156
rect 494664 87116 494670 87128
rect 502242 87116 502248 87128
rect 502300 87116 502306 87168
rect 336734 87048 336740 87100
rect 336792 87088 336798 87100
rect 346302 87088 346308 87100
rect 336792 87060 346308 87088
rect 336792 87048 336798 87060
rect 346302 87048 346308 87060
rect 346360 87048 346366 87100
rect 366910 87088 366916 87100
rect 366871 87060 366916 87088
rect 366910 87048 366916 87060
rect 366968 87048 366974 87100
rect 379054 87048 379060 87100
rect 379112 87088 379118 87100
rect 386230 87088 386236 87100
rect 379112 87060 386236 87088
rect 379112 87048 379118 87060
rect 386230 87048 386236 87060
rect 386288 87048 386294 87100
rect 396074 87048 396080 87100
rect 396132 87088 396138 87100
rect 405550 87088 405556 87100
rect 396132 87060 405556 87088
rect 396132 87048 396138 87060
rect 405550 87048 405556 87060
rect 405608 87048 405614 87100
rect 437198 87048 437204 87100
rect 437256 87088 437262 87100
rect 437474 87088 437480 87100
rect 437256 87060 437480 87088
rect 437256 87048 437262 87060
rect 437474 87048 437480 87060
rect 437532 87048 437538 87100
rect 235074 86952 235080 86964
rect 235035 86924 235080 86952
rect 235074 86912 235080 86924
rect 235132 86912 235138 86964
rect 236270 86952 236276 86964
rect 236231 86924 236276 86952
rect 236270 86912 236276 86924
rect 236328 86912 236334 86964
rect 284570 86912 284576 86964
rect 284628 86952 284634 86964
rect 284754 86952 284760 86964
rect 284628 86924 284760 86952
rect 284628 86912 284634 86924
rect 284754 86912 284760 86924
rect 284812 86912 284818 86964
rect 323302 86912 323308 86964
rect 323360 86952 323366 86964
rect 323394 86952 323400 86964
rect 323360 86924 323400 86952
rect 323360 86912 323366 86924
rect 323394 86912 323400 86924
rect 323452 86912 323458 86964
rect 324590 86912 324596 86964
rect 324648 86912 324654 86964
rect 327166 86912 327172 86964
rect 327224 86912 327230 86964
rect 341061 86955 341119 86961
rect 341061 86921 341073 86955
rect 341107 86952 341119 86955
rect 341150 86952 341156 86964
rect 341107 86924 341156 86952
rect 341107 86921 341119 86924
rect 341061 86915 341119 86921
rect 341150 86912 341156 86924
rect 341208 86912 341214 86964
rect 357618 86952 357624 86964
rect 357579 86924 357624 86952
rect 357618 86912 357624 86924
rect 357676 86912 357682 86964
rect 375834 86952 375840 86964
rect 375795 86924 375840 86952
rect 375834 86912 375840 86924
rect 375892 86912 375898 86964
rect 377122 86952 377128 86964
rect 377083 86924 377128 86952
rect 377122 86912 377128 86924
rect 377180 86912 377186 86964
rect 431310 86952 431316 86964
rect 431271 86924 431316 86952
rect 431310 86912 431316 86924
rect 431368 86912 431374 86964
rect 324608 86884 324636 86912
rect 324682 86884 324688 86896
rect 324608 86856 324688 86884
rect 324682 86844 324688 86856
rect 324740 86844 324746 86896
rect 327184 86884 327212 86912
rect 327258 86884 327264 86896
rect 327184 86856 327264 86884
rect 327258 86844 327264 86856
rect 327316 86844 327322 86896
rect 393590 86884 393596 86896
rect 393551 86856 393596 86884
rect 393590 86844 393596 86856
rect 393648 86844 393654 86896
rect 267734 85552 267740 85604
rect 267792 85552 267798 85604
rect 291562 85552 291568 85604
rect 291620 85592 291626 85604
rect 291654 85592 291660 85604
rect 291620 85564 291660 85592
rect 291620 85552 291626 85564
rect 291654 85552 291660 85564
rect 291712 85552 291718 85604
rect 294414 85552 294420 85604
rect 294472 85592 294478 85604
rect 294598 85592 294604 85604
rect 294472 85564 294604 85592
rect 294472 85552 294478 85564
rect 294598 85552 294604 85564
rect 294656 85552 294662 85604
rect 306834 85552 306840 85604
rect 306892 85592 306898 85604
rect 306926 85592 306932 85604
rect 306892 85564 306932 85592
rect 306892 85552 306898 85564
rect 306926 85552 306932 85564
rect 306984 85552 306990 85604
rect 331398 85552 331404 85604
rect 331456 85592 331462 85604
rect 331674 85592 331680 85604
rect 331456 85564 331680 85592
rect 331456 85552 331462 85564
rect 331674 85552 331680 85564
rect 331732 85552 331738 85604
rect 463697 85595 463755 85601
rect 463697 85561 463709 85595
rect 463743 85592 463755 85595
rect 463878 85592 463884 85604
rect 463743 85564 463884 85592
rect 463743 85561 463755 85564
rect 463697 85555 463755 85561
rect 463878 85552 463884 85564
rect 463936 85552 463942 85604
rect 232314 85524 232320 85536
rect 232275 85496 232320 85524
rect 232314 85484 232320 85496
rect 232372 85484 232378 85536
rect 267752 85456 267780 85552
rect 310790 85524 310796 85536
rect 310751 85496 310796 85524
rect 310790 85484 310796 85496
rect 310848 85484 310854 85536
rect 367002 85524 367008 85536
rect 366963 85496 367008 85524
rect 367002 85484 367008 85496
rect 367060 85484 367066 85536
rect 267826 85456 267832 85468
rect 267752 85428 267832 85456
rect 267826 85416 267832 85428
rect 267884 85416 267890 85468
rect 286045 84983 286103 84989
rect 286045 84949 286057 84983
rect 286091 84980 286103 84983
rect 286134 84980 286140 84992
rect 286091 84952 286140 84980
rect 286091 84949 286103 84952
rect 286045 84943 286103 84949
rect 286134 84940 286140 84952
rect 286192 84940 286198 84992
rect 262585 84303 262643 84309
rect 262585 84269 262597 84303
rect 262631 84300 262643 84303
rect 262631 84272 262720 84300
rect 262631 84269 262643 84272
rect 262585 84263 262643 84269
rect 262692 84244 262720 84272
rect 262674 84192 262680 84244
rect 262732 84192 262738 84244
rect 290090 84192 290096 84244
rect 290148 84192 290154 84244
rect 329926 84232 329932 84244
rect 329887 84204 329932 84232
rect 329926 84192 329932 84204
rect 329984 84192 329990 84244
rect 290108 84096 290136 84192
rect 290182 84096 290188 84108
rect 290108 84068 290188 84096
rect 290182 84056 290188 84068
rect 290240 84056 290246 84108
rect 295702 82832 295708 82884
rect 295760 82872 295766 82884
rect 295886 82872 295892 82884
rect 295760 82844 295892 82872
rect 295760 82832 295766 82844
rect 295886 82832 295892 82844
rect 295944 82832 295950 82884
rect 267826 82804 267832 82816
rect 267787 82776 267832 82804
rect 267826 82764 267832 82776
rect 267884 82764 267890 82816
rect 278866 80112 278872 80164
rect 278924 80112 278930 80164
rect 339770 80112 339776 80164
rect 339828 80112 339834 80164
rect 247129 80087 247187 80093
rect 247129 80053 247141 80087
rect 247175 80084 247187 80087
rect 247218 80084 247224 80096
rect 247175 80056 247224 80084
rect 247175 80053 247187 80056
rect 247129 80047 247187 80053
rect 247218 80044 247224 80056
rect 247276 80044 247282 80096
rect 278884 80028 278912 80112
rect 339788 80028 339816 80112
rect 389358 80044 389364 80096
rect 389416 80044 389422 80096
rect 273530 80016 273536 80028
rect 273491 79988 273536 80016
rect 273530 79976 273536 79988
rect 273588 79976 273594 80028
rect 278866 79976 278872 80028
rect 278924 79976 278930 80028
rect 339770 79976 339776 80028
rect 339828 79976 339834 80028
rect 389376 79948 389404 80044
rect 389450 79948 389456 79960
rect 389376 79920 389456 79948
rect 389450 79908 389456 79920
rect 389508 79908 389514 79960
rect 2774 79772 2780 79824
rect 2832 79812 2838 79824
rect 4890 79812 4896 79824
rect 2832 79784 4896 79812
rect 2832 79772 2838 79784
rect 4890 79772 4896 79784
rect 4948 79772 4954 79824
rect 296990 77364 296996 77376
rect 296824 77336 296996 77364
rect 235074 77296 235080 77308
rect 235035 77268 235080 77296
rect 235074 77256 235080 77268
rect 235132 77256 235138 77308
rect 236270 77296 236276 77308
rect 236231 77268 236276 77296
rect 236270 77256 236276 77268
rect 236328 77256 236334 77308
rect 259730 77296 259736 77308
rect 259691 77268 259736 77296
rect 259730 77256 259736 77268
rect 259788 77256 259794 77308
rect 266630 77256 266636 77308
rect 266688 77296 266694 77308
rect 266722 77296 266728 77308
rect 266688 77268 266728 77296
rect 266688 77256 266694 77268
rect 266722 77256 266728 77268
rect 266780 77256 266786 77308
rect 270681 77299 270739 77305
rect 270681 77265 270693 77299
rect 270727 77296 270739 77299
rect 270770 77296 270776 77308
rect 270727 77268 270776 77296
rect 270727 77265 270739 77268
rect 270681 77259 270739 77265
rect 270770 77256 270776 77268
rect 270828 77256 270834 77308
rect 272153 77299 272211 77305
rect 272153 77265 272165 77299
rect 272199 77296 272211 77299
rect 272242 77296 272248 77308
rect 272199 77268 272248 77296
rect 272199 77265 272211 77268
rect 272153 77259 272211 77265
rect 272242 77256 272248 77268
rect 272300 77256 272306 77308
rect 296824 77240 296852 77336
rect 296990 77324 296996 77336
rect 297048 77324 297054 77376
rect 299842 77324 299848 77376
rect 299900 77324 299906 77376
rect 330018 77324 330024 77376
rect 330076 77324 330082 77376
rect 299860 77240 299888 77324
rect 302510 77256 302516 77308
rect 302568 77296 302574 77308
rect 302602 77296 302608 77308
rect 302568 77268 302608 77296
rect 302568 77256 302574 77268
rect 302602 77256 302608 77268
rect 302660 77256 302666 77308
rect 306742 77256 306748 77308
rect 306800 77296 306806 77308
rect 306834 77296 306840 77308
rect 306800 77268 306840 77296
rect 306800 77256 306806 77268
rect 306834 77256 306840 77268
rect 306892 77256 306898 77308
rect 330036 77240 330064 77324
rect 341058 77296 341064 77308
rect 341019 77268 341064 77296
rect 341058 77256 341064 77268
rect 341116 77256 341122 77308
rect 357621 77299 357679 77305
rect 357621 77265 357633 77299
rect 357667 77296 357679 77299
rect 357710 77296 357716 77308
rect 357667 77268 357716 77296
rect 357667 77265 357679 77268
rect 357621 77259 357679 77265
rect 357710 77256 357716 77268
rect 357768 77256 357774 77308
rect 372706 77296 372712 77308
rect 372667 77268 372712 77296
rect 372706 77256 372712 77268
rect 372764 77256 372770 77308
rect 375834 77296 375840 77308
rect 375795 77268 375840 77296
rect 375834 77256 375840 77268
rect 375892 77256 375898 77308
rect 377122 77296 377128 77308
rect 377083 77268 377128 77296
rect 377122 77256 377128 77268
rect 377180 77256 377186 77308
rect 431310 77296 431316 77308
rect 431271 77268 431316 77296
rect 431310 77256 431316 77268
rect 431368 77256 431374 77308
rect 251361 77231 251419 77237
rect 251361 77197 251373 77231
rect 251407 77228 251419 77231
rect 251450 77228 251456 77240
rect 251407 77200 251456 77228
rect 251407 77197 251419 77200
rect 251361 77191 251419 77197
rect 251450 77188 251456 77200
rect 251508 77188 251514 77240
rect 296806 77188 296812 77240
rect 296864 77188 296870 77240
rect 299842 77188 299848 77240
rect 299900 77188 299906 77240
rect 330018 77188 330024 77240
rect 330076 77188 330082 77240
rect 341058 77160 341064 77172
rect 341019 77132 341064 77160
rect 341058 77120 341064 77132
rect 341116 77120 341122 77172
rect 431310 77160 431316 77172
rect 431271 77132 431316 77160
rect 431310 77120 431316 77132
rect 431368 77120 431374 77172
rect 378226 76236 378232 76288
rect 378284 76276 378290 76288
rect 386322 76276 386328 76288
rect 378284 76248 386328 76276
rect 378284 76236 378290 76248
rect 386322 76236 386328 76248
rect 386380 76236 386386 76288
rect 434714 76100 434720 76152
rect 434772 76140 434778 76152
rect 437474 76140 437480 76152
rect 434772 76112 437480 76140
rect 434772 76100 434778 76112
rect 437474 76100 437480 76112
rect 437532 76100 437538 76152
rect 463694 76100 463700 76152
rect 463752 76140 463758 76152
rect 467926 76140 467932 76152
rect 463752 76112 467932 76140
rect 463752 76100 463758 76112
rect 467926 76100 467932 76112
rect 467984 76100 467990 76152
rect 417878 76032 417884 76084
rect 417936 76072 417942 76084
rect 419350 76072 419356 76084
rect 417936 76044 419356 76072
rect 417936 76032 417942 76044
rect 419350 76032 419356 76044
rect 419408 76032 419414 76084
rect 270494 75964 270500 76016
rect 270552 76004 270558 76016
rect 275370 76004 275376 76016
rect 270552 75976 275376 76004
rect 270552 75964 270558 75976
rect 275370 75964 275376 75976
rect 275428 75964 275434 76016
rect 232314 75936 232320 75948
rect 232275 75908 232320 75936
rect 232314 75896 232320 75908
rect 232372 75896 232378 75948
rect 273530 75936 273536 75948
rect 273491 75908 273536 75936
rect 273530 75896 273536 75908
rect 273588 75896 273594 75948
rect 281810 75936 281816 75948
rect 281771 75908 281816 75936
rect 281810 75896 281816 75908
rect 281868 75896 281874 75948
rect 286045 75939 286103 75945
rect 286045 75905 286057 75939
rect 286091 75936 286103 75939
rect 286134 75936 286140 75948
rect 286091 75908 286140 75936
rect 286091 75905 286103 75908
rect 286045 75899 286103 75905
rect 286134 75896 286140 75908
rect 286192 75896 286198 75948
rect 310790 75936 310796 75948
rect 310751 75908 310796 75936
rect 310790 75896 310796 75908
rect 310848 75896 310854 75948
rect 317690 75896 317696 75948
rect 317748 75936 317754 75948
rect 317966 75936 317972 75948
rect 317748 75908 317972 75936
rect 317748 75896 317754 75908
rect 317966 75896 317972 75908
rect 318024 75896 318030 75948
rect 331398 75896 331404 75948
rect 331456 75936 331462 75948
rect 331674 75936 331680 75948
rect 331456 75908 331680 75936
rect 331456 75896 331462 75908
rect 331674 75896 331680 75908
rect 331732 75896 331738 75948
rect 367002 75936 367008 75948
rect 366963 75908 367008 75936
rect 367002 75896 367008 75908
rect 367060 75896 367066 75948
rect 389361 75871 389419 75877
rect 389361 75837 389373 75871
rect 389407 75868 389419 75871
rect 389450 75868 389456 75880
rect 389407 75840 389456 75868
rect 389407 75837 389419 75840
rect 389361 75831 389419 75837
rect 389450 75828 389456 75840
rect 389508 75828 389514 75880
rect 303890 74672 303896 74724
rect 303948 74672 303954 74724
rect 303908 74588 303936 74672
rect 291378 74536 291384 74588
rect 291436 74576 291442 74588
rect 291562 74576 291568 74588
rect 291436 74548 291568 74576
rect 291436 74536 291442 74548
rect 291562 74536 291568 74548
rect 291620 74536 291626 74588
rect 303890 74536 303896 74588
rect 303948 74536 303954 74588
rect 294233 74511 294291 74517
rect 294233 74477 294245 74511
rect 294279 74508 294291 74511
rect 294414 74508 294420 74520
rect 294279 74480 294420 74508
rect 294279 74477 294291 74480
rect 294233 74471 294291 74477
rect 294414 74468 294420 74480
rect 294472 74468 294478 74520
rect 393682 74508 393688 74520
rect 393643 74480 393688 74508
rect 393682 74468 393688 74480
rect 393740 74468 393746 74520
rect 245746 73176 245752 73228
rect 245804 73216 245810 73228
rect 245838 73216 245844 73228
rect 245804 73188 245844 73216
rect 245804 73176 245810 73188
rect 245838 73176 245844 73188
rect 245896 73176 245902 73228
rect 247126 73216 247132 73228
rect 247087 73188 247132 73216
rect 247126 73176 247132 73188
rect 247184 73176 247190 73228
rect 267829 73219 267887 73225
rect 267829 73185 267841 73219
rect 267875 73216 267887 73219
rect 267918 73216 267924 73228
rect 267875 73188 267924 73216
rect 267875 73185 267887 73188
rect 267829 73179 267887 73185
rect 267918 73176 267924 73188
rect 267976 73176 267982 73228
rect 272153 70567 272211 70573
rect 272153 70533 272165 70567
rect 272199 70564 272211 70567
rect 272242 70564 272248 70576
rect 272199 70536 272248 70564
rect 272199 70533 272211 70536
rect 272153 70527 272211 70533
rect 272242 70524 272248 70536
rect 272300 70524 272306 70576
rect 270770 70496 270776 70508
rect 270696 70468 270776 70496
rect 270696 70372 270724 70468
rect 270770 70456 270776 70468
rect 270828 70456 270834 70508
rect 327258 70496 327264 70508
rect 327184 70468 327264 70496
rect 327184 70372 327212 70468
rect 327258 70456 327264 70468
rect 327316 70456 327322 70508
rect 375834 70456 375840 70508
rect 375892 70456 375898 70508
rect 377122 70496 377128 70508
rect 377083 70468 377128 70496
rect 377122 70456 377128 70468
rect 377180 70456 377186 70508
rect 375852 70372 375880 70456
rect 270678 70320 270684 70372
rect 270736 70320 270742 70372
rect 327166 70320 327172 70372
rect 327224 70320 327230 70372
rect 375834 70320 375840 70372
rect 375892 70320 375898 70372
rect 341061 70295 341119 70301
rect 341061 70261 341073 70295
rect 341107 70292 341119 70295
rect 341150 70292 341156 70304
rect 341107 70264 341156 70292
rect 341107 70261 341119 70264
rect 341061 70255 341119 70261
rect 341150 70252 341156 70264
rect 341208 70252 341214 70304
rect 245930 67668 245936 67720
rect 245988 67668 245994 67720
rect 357710 67708 357716 67720
rect 357636 67680 357716 67708
rect 235074 67572 235080 67584
rect 235035 67544 235080 67572
rect 235074 67532 235080 67544
rect 235132 67532 235138 67584
rect 236270 67572 236276 67584
rect 236231 67544 236276 67572
rect 236270 67532 236276 67544
rect 236328 67532 236334 67584
rect 245948 67516 245976 67668
rect 357636 67652 357664 67680
rect 357710 67668 357716 67680
rect 357768 67668 357774 67720
rect 265158 67600 265164 67652
rect 265216 67640 265222 67652
rect 265250 67640 265256 67652
rect 265216 67612 265256 67640
rect 265216 67600 265222 67612
rect 265250 67600 265256 67612
rect 265308 67600 265314 67652
rect 272150 67640 272156 67652
rect 272111 67612 272156 67640
rect 272150 67600 272156 67612
rect 272208 67600 272214 67652
rect 281718 67600 281724 67652
rect 281776 67640 281782 67652
rect 281810 67640 281816 67652
rect 281776 67612 281816 67640
rect 281776 67600 281782 67612
rect 281810 67600 281816 67612
rect 281868 67600 281874 67652
rect 291378 67600 291384 67652
rect 291436 67640 291442 67652
rect 291470 67640 291476 67652
rect 291436 67612 291476 67640
rect 291436 67600 291442 67612
rect 291470 67600 291476 67612
rect 291528 67600 291534 67652
rect 299750 67600 299756 67652
rect 299808 67640 299814 67652
rect 299842 67640 299848 67652
rect 299808 67612 299848 67640
rect 299808 67600 299814 67612
rect 299842 67600 299848 67612
rect 299900 67600 299906 67652
rect 301038 67600 301044 67652
rect 301096 67640 301102 67652
rect 301222 67640 301228 67652
rect 301096 67612 301228 67640
rect 301096 67600 301102 67612
rect 301222 67600 301228 67612
rect 301280 67600 301286 67652
rect 329926 67600 329932 67652
rect 329984 67640 329990 67652
rect 330110 67640 330116 67652
rect 329984 67612 330116 67640
rect 329984 67600 329990 67612
rect 330110 67600 330116 67612
rect 330168 67600 330174 67652
rect 357618 67600 357624 67652
rect 357676 67600 357682 67652
rect 377122 67640 377128 67652
rect 377083 67612 377128 67640
rect 377122 67600 377128 67612
rect 377180 67600 377186 67652
rect 431313 67643 431371 67649
rect 431313 67609 431325 67643
rect 431359 67640 431371 67643
rect 431402 67640 431408 67652
rect 431359 67612 431408 67640
rect 431359 67609 431371 67612
rect 431313 67603 431371 67609
rect 431402 67600 431408 67612
rect 431460 67600 431466 67652
rect 459922 67532 459928 67584
rect 459980 67572 459986 67584
rect 460198 67572 460204 67584
rect 459980 67544 460204 67572
rect 459980 67532 459986 67544
rect 460198 67532 460204 67544
rect 460256 67532 460262 67584
rect 245930 67464 245936 67516
rect 245988 67464 245994 67516
rect 389358 66280 389364 66292
rect 389319 66252 389364 66280
rect 389358 66240 389364 66252
rect 389416 66240 389422 66292
rect 232314 66172 232320 66224
rect 232372 66172 232378 66224
rect 244366 66212 244372 66224
rect 244327 66184 244372 66212
rect 244366 66172 244372 66184
rect 244424 66172 244430 66224
rect 245930 66172 245936 66224
rect 245988 66212 245994 66224
rect 245988 66184 246068 66212
rect 245988 66172 245994 66184
rect 232332 66085 232360 66172
rect 246040 66156 246068 66184
rect 265158 66172 265164 66224
rect 265216 66212 265222 66224
rect 265253 66215 265311 66221
rect 265253 66212 265265 66215
rect 265216 66184 265265 66212
rect 265216 66172 265222 66184
rect 265253 66181 265265 66184
rect 265299 66181 265311 66215
rect 273530 66212 273536 66224
rect 273491 66184 273536 66212
rect 265253 66175 265311 66181
rect 273530 66172 273536 66184
rect 273588 66172 273594 66224
rect 302510 66172 302516 66224
rect 302568 66212 302574 66224
rect 302694 66212 302700 66224
rect 302568 66184 302700 66212
rect 302568 66172 302574 66184
rect 302694 66172 302700 66184
rect 302752 66172 302758 66224
rect 306742 66172 306748 66224
rect 306800 66212 306806 66224
rect 306926 66212 306932 66224
rect 306800 66184 306932 66212
rect 306800 66172 306806 66184
rect 306926 66172 306932 66184
rect 306984 66172 306990 66224
rect 310790 66212 310796 66224
rect 310751 66184 310796 66212
rect 310790 66172 310796 66184
rect 310848 66172 310854 66224
rect 323394 66212 323400 66224
rect 323355 66184 323400 66212
rect 323394 66172 323400 66184
rect 323452 66172 323458 66224
rect 327166 66212 327172 66224
rect 327127 66184 327172 66212
rect 327166 66172 327172 66184
rect 327224 66172 327230 66224
rect 367002 66212 367008 66224
rect 366963 66184 367008 66212
rect 367002 66172 367008 66184
rect 367060 66172 367066 66224
rect 246022 66104 246028 66156
rect 246080 66104 246086 66156
rect 232317 66079 232375 66085
rect 232317 66045 232329 66079
rect 232363 66045 232375 66079
rect 232317 66039 232375 66045
rect 267918 64988 267924 65000
rect 267752 64960 267924 64988
rect 267752 64932 267780 64960
rect 267918 64948 267924 64960
rect 267976 64948 267982 65000
rect 251358 64920 251364 64932
rect 251319 64892 251364 64920
rect 251358 64880 251364 64892
rect 251416 64880 251422 64932
rect 267734 64880 267740 64932
rect 267792 64880 267798 64932
rect 294230 64920 294236 64932
rect 294191 64892 294236 64920
rect 294230 64880 294236 64892
rect 294288 64880 294294 64932
rect 295610 64880 295616 64932
rect 295668 64920 295674 64932
rect 295702 64920 295708 64932
rect 295668 64892 295708 64920
rect 295668 64880 295674 64892
rect 295702 64880 295708 64892
rect 295760 64880 295766 64932
rect 393685 64923 393743 64929
rect 393685 64889 393697 64923
rect 393731 64920 393743 64923
rect 393774 64920 393780 64932
rect 393731 64892 393780 64920
rect 393731 64889 393743 64892
rect 393685 64883 393743 64889
rect 393774 64880 393780 64892
rect 393832 64880 393838 64932
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 31018 64852 31024 64864
rect 3384 64824 31024 64852
rect 3384 64812 3390 64824
rect 31018 64812 31024 64824
rect 31076 64812 31082 64864
rect 378226 63860 378232 63912
rect 378284 63900 378290 63912
rect 386322 63900 386328 63912
rect 378284 63872 386328 63900
rect 378284 63860 378290 63872
rect 386322 63860 386328 63872
rect 386380 63860 386386 63912
rect 417878 63656 417884 63708
rect 417936 63696 417942 63708
rect 418154 63696 418160 63708
rect 417936 63668 418160 63696
rect 417936 63656 417942 63668
rect 418154 63656 418160 63668
rect 418212 63656 418218 63708
rect 437198 63656 437204 63708
rect 437256 63696 437262 63708
rect 437474 63696 437480 63708
rect 437256 63668 437480 63696
rect 437256 63656 437262 63668
rect 437474 63656 437480 63668
rect 437532 63656 437538 63708
rect 456518 63656 456524 63708
rect 456576 63696 456582 63708
rect 456886 63696 456892 63708
rect 456576 63668 456892 63696
rect 456576 63656 456582 63668
rect 456886 63656 456892 63668
rect 456944 63656 456950 63708
rect 303890 63492 303896 63504
rect 303851 63464 303896 63492
rect 303890 63452 303896 63464
rect 303948 63452 303954 63504
rect 235074 62744 235080 62756
rect 235035 62716 235080 62744
rect 235074 62704 235080 62716
rect 235132 62704 235138 62756
rect 259730 62636 259736 62688
rect 259788 62636 259794 62688
rect 259748 62608 259776 62636
rect 259914 62608 259920 62620
rect 259748 62580 259920 62608
rect 259914 62568 259920 62580
rect 259972 62568 259978 62620
rect 262766 61412 262772 61464
rect 262824 61452 262830 61464
rect 262950 61452 262956 61464
rect 262824 61424 262956 61452
rect 262824 61412 262830 61424
rect 262950 61412 262956 61424
rect 263008 61412 263014 61464
rect 281718 61452 281724 61464
rect 281679 61424 281724 61452
rect 281718 61412 281724 61424
rect 281776 61412 281782 61464
rect 295521 61455 295579 61461
rect 295521 61421 295533 61455
rect 295567 61452 295579 61455
rect 295610 61452 295616 61464
rect 295567 61424 295616 61452
rect 295567 61421 295579 61424
rect 295521 61415 295579 61421
rect 295610 61412 295616 61424
rect 295668 61412 295674 61464
rect 330110 61452 330116 61464
rect 330071 61424 330116 61452
rect 330110 61412 330116 61424
rect 330168 61412 330174 61464
rect 267734 60800 267740 60852
rect 267792 60800 267798 60852
rect 324590 60800 324596 60852
rect 324648 60800 324654 60852
rect 337194 60800 337200 60852
rect 337252 60800 337258 60852
rect 339770 60840 339776 60852
rect 339731 60812 339776 60840
rect 339770 60800 339776 60812
rect 339828 60800 339834 60852
rect 266630 60732 266636 60784
rect 266688 60732 266694 60784
rect 230753 60639 230811 60645
rect 230753 60605 230765 60639
rect 230799 60636 230811 60639
rect 230842 60636 230848 60648
rect 230799 60608 230848 60636
rect 230799 60605 230811 60608
rect 230753 60599 230811 60605
rect 230842 60596 230848 60608
rect 230900 60596 230906 60648
rect 266648 60636 266676 60732
rect 267752 60716 267780 60800
rect 324608 60716 324636 60800
rect 325878 60732 325884 60784
rect 325936 60732 325942 60784
rect 267734 60664 267740 60716
rect 267792 60664 267798 60716
rect 310790 60704 310796 60716
rect 310751 60676 310796 60704
rect 310790 60664 310796 60676
rect 310848 60664 310854 60716
rect 324590 60664 324596 60716
rect 324648 60664 324654 60716
rect 266722 60636 266728 60648
rect 266648 60608 266728 60636
rect 266722 60596 266728 60608
rect 266780 60596 266786 60648
rect 325896 60636 325924 60732
rect 337212 60648 337240 60800
rect 325970 60636 325976 60648
rect 325896 60608 325976 60636
rect 325970 60596 325976 60608
rect 326028 60596 326034 60648
rect 337194 60596 337200 60648
rect 337252 60596 337258 60648
rect 270678 58012 270684 58064
rect 270736 58012 270742 58064
rect 284754 58012 284760 58064
rect 284812 58012 284818 58064
rect 291470 58052 291476 58064
rect 291396 58024 291476 58052
rect 236270 57984 236276 57996
rect 236231 57956 236276 57984
rect 236270 57944 236276 57956
rect 236328 57944 236334 57996
rect 270696 57928 270724 58012
rect 272150 57944 272156 57996
rect 272208 57984 272214 57996
rect 272242 57984 272248 57996
rect 272208 57956 272248 57984
rect 272208 57944 272214 57956
rect 272242 57944 272248 57956
rect 272300 57944 272306 57996
rect 284772 57928 284800 58012
rect 291396 57928 291424 58024
rect 291470 58012 291476 58024
rect 291528 58012 291534 58064
rect 270678 57876 270684 57928
rect 270736 57876 270742 57928
rect 284754 57876 284760 57928
rect 284812 57876 284818 57928
rect 291378 57876 291384 57928
rect 291436 57876 291442 57928
rect 357621 57919 357679 57925
rect 357621 57885 357633 57919
rect 357667 57916 357679 57919
rect 357710 57916 357716 57928
rect 357667 57888 357716 57916
rect 357667 57885 357679 57888
rect 357621 57879 357679 57885
rect 357710 57876 357716 57888
rect 357768 57876 357774 57928
rect 460017 57919 460075 57925
rect 460017 57885 460029 57919
rect 460063 57916 460075 57919
rect 460106 57916 460112 57928
rect 460063 57888 460112 57916
rect 460063 57885 460075 57888
rect 460017 57879 460075 57885
rect 460106 57876 460112 57888
rect 460164 57876 460170 57928
rect 330113 57851 330171 57857
rect 330113 57817 330125 57851
rect 330159 57848 330171 57851
rect 330294 57848 330300 57860
rect 330159 57820 330300 57848
rect 330159 57817 330171 57820
rect 330113 57811 330171 57817
rect 330294 57808 330300 57820
rect 330352 57808 330358 57860
rect 389177 57579 389235 57585
rect 389177 57545 389189 57579
rect 389223 57576 389235 57579
rect 389358 57576 389364 57588
rect 389223 57548 389364 57576
rect 389223 57545 389235 57548
rect 389177 57539 389235 57545
rect 389358 57536 389364 57548
rect 389416 57536 389422 57588
rect 288710 57032 288716 57044
rect 288671 57004 288716 57032
rect 288710 56992 288716 57004
rect 288768 56992 288774 57044
rect 232314 56624 232320 56636
rect 232275 56596 232320 56624
rect 232314 56584 232320 56596
rect 232372 56584 232378 56636
rect 244369 56627 244427 56633
rect 244369 56593 244381 56627
rect 244415 56624 244427 56627
rect 244458 56624 244464 56636
rect 244415 56596 244464 56624
rect 244415 56593 244427 56596
rect 244369 56587 244427 56593
rect 244458 56584 244464 56596
rect 244516 56584 244522 56636
rect 250162 56624 250168 56636
rect 250123 56596 250168 56624
rect 250162 56584 250168 56596
rect 250220 56584 250226 56636
rect 273530 56624 273536 56636
rect 273491 56596 273536 56624
rect 273530 56584 273536 56596
rect 273588 56584 273594 56636
rect 323394 56624 323400 56636
rect 323355 56596 323400 56624
rect 323394 56584 323400 56596
rect 323452 56584 323458 56636
rect 327169 56627 327227 56633
rect 327169 56593 327181 56627
rect 327215 56624 327227 56627
rect 327442 56624 327448 56636
rect 327215 56596 327448 56624
rect 327215 56593 327227 56596
rect 327169 56587 327227 56593
rect 327442 56584 327448 56596
rect 327500 56584 327506 56636
rect 339770 56624 339776 56636
rect 339731 56596 339776 56624
rect 339770 56584 339776 56596
rect 339828 56584 339834 56636
rect 259914 56516 259920 56568
rect 259972 56556 259978 56568
rect 259972 56528 260017 56556
rect 259972 56516 259978 56528
rect 310790 56516 310796 56568
rect 310848 56556 310854 56568
rect 310882 56556 310888 56568
rect 310848 56528 310888 56556
rect 310848 56516 310854 56528
rect 310882 56516 310888 56528
rect 310940 56516 310946 56568
rect 341334 56556 341340 56568
rect 341295 56528 341340 56556
rect 341334 56516 341340 56528
rect 341392 56516 341398 56568
rect 317506 55224 317512 55276
rect 317564 55264 317570 55276
rect 317690 55264 317696 55276
rect 317564 55236 317696 55264
rect 317564 55224 317570 55236
rect 317690 55224 317696 55236
rect 317748 55224 317754 55276
rect 393498 55224 393504 55276
rect 393556 55264 393562 55276
rect 393774 55264 393780 55276
rect 393556 55236 393780 55264
rect 393556 55224 393562 55236
rect 393774 55224 393780 55236
rect 393832 55224 393838 55276
rect 247218 55196 247224 55208
rect 247179 55168 247224 55196
rect 247218 55156 247224 55168
rect 247276 55156 247282 55208
rect 250162 53836 250168 53848
rect 250123 53808 250168 53836
rect 250162 53796 250168 53808
rect 250220 53796 250226 53848
rect 303893 53839 303951 53845
rect 303893 53805 303905 53839
rect 303939 53836 303951 53839
rect 303982 53836 303988 53848
rect 303939 53808 303988 53836
rect 303939 53805 303951 53808
rect 303893 53799 303951 53805
rect 303982 53796 303988 53808
rect 304040 53796 304046 53848
rect 278866 51184 278872 51196
rect 278827 51156 278872 51184
rect 278866 51144 278872 51156
rect 278924 51144 278930 51196
rect 375834 51144 375840 51196
rect 375892 51144 375898 51196
rect 232314 51116 232320 51128
rect 232240 51088 232320 51116
rect 232240 51060 232268 51088
rect 232314 51076 232320 51088
rect 232372 51076 232378 51128
rect 273530 51076 273536 51128
rect 273588 51076 273594 51128
rect 337105 51119 337163 51125
rect 337105 51085 337117 51119
rect 337151 51116 337163 51119
rect 337194 51116 337200 51128
rect 337151 51088 337200 51116
rect 337151 51085 337163 51088
rect 337105 51079 337163 51085
rect 337194 51076 337200 51088
rect 337252 51076 337258 51128
rect 232222 51008 232228 51060
rect 232280 51008 232286 51060
rect 273548 50924 273576 51076
rect 375852 51060 375880 51144
rect 375834 51008 375840 51060
rect 375892 51008 375898 51060
rect 265158 50872 265164 50924
rect 265216 50912 265222 50924
rect 265253 50915 265311 50921
rect 265253 50912 265265 50915
rect 265216 50884 265265 50912
rect 265216 50872 265222 50884
rect 265253 50881 265265 50884
rect 265299 50881 265311 50915
rect 265253 50875 265311 50881
rect 273530 50872 273536 50924
rect 273588 50872 273594 50924
rect 341334 50640 341340 50652
rect 341295 50612 341340 50640
rect 341334 50600 341340 50612
rect 341392 50600 341398 50652
rect 2774 50464 2780 50516
rect 2832 50504 2838 50516
rect 4798 50504 4804 50516
rect 2832 50476 4804 50504
rect 2832 50464 2838 50476
rect 4798 50464 4804 50476
rect 4856 50464 4862 50516
rect 367002 48396 367008 48408
rect 366963 48368 367008 48396
rect 367002 48356 367008 48368
rect 367060 48356 367066 48408
rect 230750 48328 230756 48340
rect 230711 48300 230756 48328
rect 230750 48288 230756 48300
rect 230808 48288 230814 48340
rect 244366 48288 244372 48340
rect 244424 48328 244430 48340
rect 244550 48328 244556 48340
rect 244424 48300 244556 48328
rect 244424 48288 244430 48300
rect 244550 48288 244556 48300
rect 244608 48288 244614 48340
rect 278866 48328 278872 48340
rect 278827 48300 278872 48328
rect 278866 48288 278872 48300
rect 278924 48288 278930 48340
rect 281718 48328 281724 48340
rect 281679 48300 281724 48328
rect 281718 48288 281724 48300
rect 281776 48288 281782 48340
rect 284662 48288 284668 48340
rect 284720 48328 284726 48340
rect 284754 48328 284760 48340
rect 284720 48300 284760 48328
rect 284720 48288 284726 48300
rect 284754 48288 284760 48300
rect 284812 48288 284818 48340
rect 288710 48328 288716 48340
rect 288671 48300 288716 48328
rect 288710 48288 288716 48300
rect 288768 48288 288774 48340
rect 291378 48288 291384 48340
rect 291436 48328 291442 48340
rect 291470 48328 291476 48340
rect 291436 48300 291476 48328
rect 291436 48288 291442 48300
rect 291470 48288 291476 48300
rect 291528 48288 291534 48340
rect 295518 48328 295524 48340
rect 295479 48300 295524 48328
rect 295518 48288 295524 48300
rect 295576 48288 295582 48340
rect 299750 48288 299756 48340
rect 299808 48288 299814 48340
rect 301038 48288 301044 48340
rect 301096 48288 301102 48340
rect 325878 48288 325884 48340
rect 325936 48328 325942 48340
rect 326062 48328 326068 48340
rect 325936 48300 326068 48328
rect 325936 48288 325942 48300
rect 326062 48288 326068 48300
rect 326120 48288 326126 48340
rect 327350 48328 327356 48340
rect 327311 48300 327356 48328
rect 327350 48288 327356 48300
rect 327408 48288 327414 48340
rect 337102 48328 337108 48340
rect 337063 48300 337108 48328
rect 337102 48288 337108 48300
rect 337160 48288 337166 48340
rect 357618 48328 357624 48340
rect 357579 48300 357624 48328
rect 357618 48288 357624 48300
rect 357676 48288 357682 48340
rect 389177 48331 389235 48337
rect 389177 48297 389189 48331
rect 389223 48328 389235 48331
rect 389266 48328 389272 48340
rect 389223 48300 389272 48328
rect 389223 48297 389235 48300
rect 389177 48291 389235 48297
rect 389266 48288 389272 48300
rect 389324 48288 389330 48340
rect 460014 48328 460020 48340
rect 459975 48300 460020 48328
rect 460014 48288 460020 48300
rect 460072 48288 460078 48340
rect 236270 48260 236276 48272
rect 236231 48232 236276 48260
rect 236270 48220 236276 48232
rect 236328 48220 236334 48272
rect 299768 48192 299796 48288
rect 299842 48192 299848 48204
rect 299768 48164 299848 48192
rect 299842 48152 299848 48164
rect 299900 48152 299906 48204
rect 301056 48192 301084 48288
rect 323302 48220 323308 48272
rect 323360 48260 323366 48272
rect 323394 48260 323400 48272
rect 323360 48232 323400 48260
rect 323360 48220 323366 48232
rect 323394 48220 323400 48232
rect 323452 48220 323458 48272
rect 301130 48192 301136 48204
rect 301056 48164 301136 48192
rect 301130 48152 301136 48164
rect 301188 48152 301194 48204
rect 460014 48192 460020 48204
rect 459975 48164 460020 48192
rect 460014 48152 460020 48164
rect 460072 48152 460078 48204
rect 250162 47036 250168 47048
rect 250088 47008 250168 47036
rect 250088 46912 250116 47008
rect 250162 46996 250168 47008
rect 250220 46996 250226 47048
rect 327350 46968 327356 46980
rect 327311 46940 327356 46968
rect 327350 46928 327356 46940
rect 327408 46928 327414 46980
rect 250070 46860 250076 46912
rect 250128 46860 250134 46912
rect 265158 46900 265164 46912
rect 265119 46872 265164 46900
rect 265158 46860 265164 46872
rect 265216 46860 265222 46912
rect 266722 46900 266728 46912
rect 266683 46872 266728 46900
rect 266722 46860 266728 46872
rect 266780 46860 266786 46912
rect 284662 46860 284668 46912
rect 284720 46900 284726 46912
rect 284757 46903 284815 46909
rect 284757 46900 284769 46903
rect 284720 46872 284769 46900
rect 284720 46860 284726 46872
rect 284757 46869 284769 46872
rect 284803 46869 284815 46903
rect 284757 46863 284815 46869
rect 286042 46860 286048 46912
rect 286100 46900 286106 46912
rect 286134 46900 286140 46912
rect 286100 46872 286140 46900
rect 286100 46860 286106 46872
rect 286134 46860 286140 46872
rect 286192 46860 286198 46912
rect 291470 46900 291476 46912
rect 291431 46872 291476 46900
rect 291470 46860 291476 46872
rect 291528 46860 291534 46912
rect 323302 46900 323308 46912
rect 323263 46872 323308 46900
rect 323302 46860 323308 46872
rect 323360 46860 323366 46912
rect 339770 46900 339776 46912
rect 339731 46872 339776 46900
rect 339770 46860 339776 46872
rect 339828 46860 339834 46912
rect 366821 46903 366879 46909
rect 366821 46869 366833 46903
rect 366867 46900 366879 46903
rect 367002 46900 367008 46912
rect 366867 46872 367008 46900
rect 366867 46869 366879 46872
rect 366821 46863 366879 46869
rect 367002 46860 367008 46872
rect 367060 46860 367066 46912
rect 375742 46860 375748 46912
rect 375800 46900 375806 46912
rect 375834 46900 375840 46912
rect 375800 46872 375840 46900
rect 375800 46860 375806 46872
rect 375834 46860 375840 46872
rect 375892 46860 375898 46912
rect 377030 46860 377036 46912
rect 377088 46900 377094 46912
rect 377122 46900 377128 46912
rect 377088 46872 377128 46900
rect 377088 46860 377094 46872
rect 377122 46860 377128 46872
rect 377180 46860 377186 46912
rect 259917 45679 259975 45685
rect 259917 45676 259929 45679
rect 259748 45648 259929 45676
rect 259748 45620 259776 45648
rect 259917 45645 259929 45648
rect 259963 45645 259975 45679
rect 259917 45639 259975 45645
rect 247218 45608 247224 45620
rect 247179 45580 247224 45608
rect 247218 45568 247224 45580
rect 247276 45568 247282 45620
rect 259730 45568 259736 45620
rect 259788 45568 259794 45620
rect 393406 45568 393412 45620
rect 393464 45608 393470 45620
rect 393682 45608 393688 45620
rect 393464 45580 393688 45608
rect 393464 45568 393470 45580
rect 393682 45568 393688 45580
rect 393740 45568 393746 45620
rect 251358 45540 251364 45552
rect 251319 45512 251364 45540
rect 251358 45500 251364 45512
rect 251416 45500 251422 45552
rect 299753 45543 299811 45549
rect 299753 45509 299765 45543
rect 299799 45540 299811 45543
rect 299842 45540 299848 45552
rect 299799 45512 299848 45540
rect 299799 45509 299811 45512
rect 299753 45503 299811 45509
rect 299842 45500 299848 45512
rect 299900 45500 299906 45552
rect 310882 45500 310888 45552
rect 310940 45540 310946 45552
rect 311066 45540 311072 45552
rect 310940 45512 311072 45540
rect 310940 45500 310946 45512
rect 311066 45500 311072 45512
rect 311124 45500 311130 45552
rect 317506 45500 317512 45552
rect 317564 45540 317570 45552
rect 317690 45540 317696 45552
rect 317564 45512 317696 45540
rect 317564 45500 317570 45512
rect 317690 45500 317696 45512
rect 317748 45500 317754 45552
rect 245746 44112 245752 44124
rect 245707 44084 245752 44112
rect 245746 44072 245752 44084
rect 245804 44072 245810 44124
rect 303798 42372 303804 42424
rect 303856 42412 303862 42424
rect 304074 42412 304080 42424
rect 303856 42384 304080 42412
rect 303856 42372 303862 42384
rect 304074 42372 304080 42384
rect 304132 42372 304138 42424
rect 339770 42072 339776 42084
rect 339731 42044 339776 42072
rect 339770 42032 339776 42044
rect 339828 42032 339834 42084
rect 460017 41395 460075 41401
rect 460017 41361 460029 41395
rect 460063 41392 460075 41395
rect 460198 41392 460204 41404
rect 460063 41364 460204 41392
rect 460063 41361 460075 41364
rect 460017 41355 460075 41361
rect 460198 41352 460204 41364
rect 460256 41352 460262 41404
rect 306926 40780 306932 40792
rect 306887 40752 306932 40780
rect 306926 40740 306932 40752
rect 306984 40740 306990 40792
rect 245562 40332 245568 40384
rect 245620 40372 245626 40384
rect 245930 40372 245936 40384
rect 245620 40344 245936 40372
rect 245620 40332 245626 40344
rect 245930 40332 245936 40344
rect 245988 40332 245994 40384
rect 437198 40196 437204 40248
rect 437256 40236 437262 40248
rect 437566 40236 437572 40248
rect 437256 40208 437572 40236
rect 437256 40196 437262 40208
rect 437566 40196 437572 40208
rect 437624 40196 437630 40248
rect 456518 40196 456524 40248
rect 456576 40236 456582 40248
rect 456886 40236 456892 40248
rect 456576 40208 456892 40236
rect 456576 40196 456582 40208
rect 456886 40196 456892 40208
rect 456944 40196 456950 40248
rect 417878 40128 417884 40180
rect 417936 40168 417942 40180
rect 418154 40168 418160 40180
rect 417936 40140 418160 40168
rect 417936 40128 417942 40140
rect 418154 40128 418160 40140
rect 418212 40128 418218 40180
rect 230750 38740 230756 38752
rect 230711 38712 230756 38740
rect 230750 38700 230756 38712
rect 230808 38700 230814 38752
rect 244366 38700 244372 38752
rect 244424 38700 244430 38752
rect 267918 38700 267924 38752
rect 267976 38700 267982 38752
rect 325878 38700 325884 38752
rect 325936 38700 325942 38752
rect 366910 38700 366916 38752
rect 366968 38700 366974 38752
rect 236270 38672 236276 38684
rect 236231 38644 236276 38672
rect 236270 38632 236276 38644
rect 236328 38632 236334 38684
rect 244384 38672 244412 38700
rect 244458 38672 244464 38684
rect 244384 38644 244464 38672
rect 244458 38632 244464 38644
rect 244516 38632 244522 38684
rect 267936 38616 267964 38700
rect 270678 38632 270684 38684
rect 270736 38672 270742 38684
rect 270770 38672 270776 38684
rect 270736 38644 270776 38672
rect 270736 38632 270742 38644
rect 270770 38632 270776 38644
rect 270828 38632 270834 38684
rect 272150 38632 272156 38684
rect 272208 38672 272214 38684
rect 272242 38672 272248 38684
rect 272208 38644 272248 38672
rect 272208 38632 272214 38644
rect 272242 38632 272248 38644
rect 272300 38632 272306 38684
rect 324590 38632 324596 38684
rect 324648 38672 324654 38684
rect 324682 38672 324688 38684
rect 324648 38644 324688 38672
rect 324648 38632 324654 38644
rect 324682 38632 324688 38644
rect 324740 38632 324746 38684
rect 325896 38616 325924 38700
rect 327258 38632 327264 38684
rect 327316 38672 327322 38684
rect 327350 38672 327356 38684
rect 327316 38644 327356 38672
rect 327316 38632 327322 38644
rect 327350 38632 327356 38644
rect 327408 38632 327414 38684
rect 329926 38632 329932 38684
rect 329984 38672 329990 38684
rect 330202 38672 330208 38684
rect 329984 38644 330208 38672
rect 329984 38632 329990 38644
rect 330202 38632 330208 38644
rect 330260 38632 330266 38684
rect 331122 38632 331128 38684
rect 331180 38672 331186 38684
rect 331490 38672 331496 38684
rect 331180 38644 331496 38672
rect 331180 38632 331186 38644
rect 331490 38632 331496 38644
rect 331548 38632 331554 38684
rect 366928 38616 366956 38700
rect 267918 38564 267924 38616
rect 267976 38564 267982 38616
rect 281718 38604 281724 38616
rect 281679 38576 281724 38604
rect 281718 38564 281724 38576
rect 281776 38564 281782 38616
rect 325878 38564 325884 38616
rect 325936 38564 325942 38616
rect 366910 38564 366916 38616
rect 366968 38564 366974 38616
rect 372706 38564 372712 38616
rect 372764 38604 372770 38616
rect 372798 38604 372804 38616
rect 372764 38576 372804 38604
rect 372764 38564 372770 38576
rect 372798 38564 372804 38576
rect 372856 38564 372862 38616
rect 460109 38607 460167 38613
rect 460109 38573 460121 38607
rect 460155 38604 460167 38607
rect 460198 38604 460204 38616
rect 460155 38576 460204 38604
rect 460155 38573 460167 38576
rect 460109 38567 460167 38573
rect 460198 38564 460204 38576
rect 460256 38564 460262 38616
rect 232314 37380 232320 37392
rect 232240 37352 232320 37380
rect 232240 37324 232268 37352
rect 232314 37340 232320 37352
rect 232372 37340 232378 37392
rect 230750 37312 230756 37324
rect 230711 37284 230756 37312
rect 230750 37272 230756 37284
rect 230808 37272 230814 37324
rect 232222 37272 232228 37324
rect 232280 37272 232286 37324
rect 265158 37312 265164 37324
rect 265119 37284 265164 37312
rect 265158 37272 265164 37284
rect 265216 37272 265222 37324
rect 266722 37312 266728 37324
rect 266683 37284 266728 37312
rect 266722 37272 266728 37284
rect 266780 37272 266786 37324
rect 284754 37272 284760 37324
rect 284812 37312 284818 37324
rect 323302 37312 323308 37324
rect 284812 37284 284857 37312
rect 323263 37284 323308 37312
rect 284812 37272 284818 37284
rect 323302 37272 323308 37284
rect 323360 37272 323366 37324
rect 366818 37312 366824 37324
rect 366779 37284 366824 37312
rect 366818 37272 366824 37284
rect 366876 37272 366882 37324
rect 389174 37272 389180 37324
rect 389232 37312 389238 37324
rect 389358 37312 389364 37324
rect 389232 37284 389364 37312
rect 389232 37272 389238 37284
rect 389358 37272 389364 37284
rect 389416 37272 389422 37324
rect 270770 37204 270776 37256
rect 270828 37244 270834 37256
rect 270862 37244 270868 37256
rect 270828 37216 270868 37244
rect 270828 37204 270834 37216
rect 270862 37204 270868 37216
rect 270920 37204 270926 37256
rect 288802 37204 288808 37256
rect 288860 37244 288866 37256
rect 288894 37244 288900 37256
rect 288860 37216 288900 37244
rect 288860 37204 288866 37216
rect 288894 37204 288900 37216
rect 288952 37204 288958 37256
rect 393590 37244 393596 37256
rect 393551 37216 393596 37244
rect 393590 37204 393596 37216
rect 393648 37204 393654 37256
rect 232222 37176 232228 37188
rect 232183 37148 232228 37176
rect 232222 37136 232228 37148
rect 232280 37136 232286 37188
rect 259638 37136 259644 37188
rect 259696 37176 259702 37188
rect 259730 37176 259736 37188
rect 259696 37148 259736 37176
rect 259696 37136 259702 37148
rect 259730 37136 259736 37148
rect 259788 37136 259794 37188
rect 249978 35912 249984 35964
rect 250036 35952 250042 35964
rect 250070 35952 250076 35964
rect 250036 35924 250076 35952
rect 250036 35912 250042 35924
rect 250070 35912 250076 35924
rect 250128 35912 250134 35964
rect 251361 35955 251419 35961
rect 251361 35921 251373 35955
rect 251407 35952 251419 35955
rect 251450 35952 251456 35964
rect 251407 35924 251456 35952
rect 251407 35921 251419 35924
rect 251361 35915 251419 35921
rect 251450 35912 251456 35924
rect 251508 35912 251514 35964
rect 291473 35955 291531 35961
rect 291473 35921 291485 35955
rect 291519 35952 291531 35955
rect 291562 35952 291568 35964
rect 291519 35924 291568 35952
rect 291519 35921 291531 35924
rect 291473 35915 291531 35921
rect 291562 35912 291568 35924
rect 291620 35912 291626 35964
rect 299750 35952 299756 35964
rect 299711 35924 299756 35952
rect 299750 35912 299756 35924
rect 299808 35912 299814 35964
rect 306742 35912 306748 35964
rect 306800 35952 306806 35964
rect 306929 35955 306987 35961
rect 306929 35952 306941 35955
rect 306800 35924 306941 35952
rect 306800 35912 306806 35924
rect 306929 35921 306941 35924
rect 306975 35921 306987 35955
rect 306929 35915 306987 35921
rect 3142 35844 3148 35896
rect 3200 35884 3206 35896
rect 6178 35884 6184 35896
rect 3200 35856 6184 35884
rect 3200 35844 3206 35856
rect 6178 35844 6184 35856
rect 6236 35844 6242 35896
rect 247218 35884 247224 35896
rect 247179 35856 247224 35884
rect 247218 35844 247224 35856
rect 247276 35844 247282 35896
rect 259549 35887 259607 35893
rect 259549 35853 259561 35887
rect 259595 35884 259607 35887
rect 259638 35884 259644 35896
rect 259595 35856 259644 35884
rect 259595 35853 259607 35856
rect 259549 35847 259607 35853
rect 259638 35844 259644 35856
rect 259696 35844 259702 35896
rect 270773 35887 270831 35893
rect 270773 35853 270785 35887
rect 270819 35884 270831 35887
rect 270862 35884 270868 35896
rect 270819 35856 270868 35884
rect 270819 35853 270831 35856
rect 270773 35847 270831 35853
rect 270862 35844 270868 35856
rect 270920 35844 270926 35896
rect 294138 35844 294144 35896
rect 294196 35884 294202 35896
rect 294506 35884 294512 35896
rect 294196 35856 294512 35884
rect 294196 35844 294202 35856
rect 294506 35844 294512 35856
rect 294564 35844 294570 35896
rect 250070 35816 250076 35828
rect 250031 35788 250076 35816
rect 250070 35776 250076 35788
rect 250128 35776 250134 35828
rect 245746 34524 245752 34536
rect 245707 34496 245752 34524
rect 245746 34484 245752 34496
rect 245804 34484 245810 34536
rect 317506 31764 317512 31816
rect 317564 31804 317570 31816
rect 317690 31804 317696 31816
rect 317564 31776 317696 31804
rect 317564 31764 317570 31776
rect 317690 31764 317696 31776
rect 317748 31764 317754 31816
rect 339681 31807 339739 31813
rect 339681 31773 339693 31807
rect 339727 31804 339739 31807
rect 339770 31804 339776 31816
rect 339727 31776 339776 31804
rect 339727 31773 339739 31776
rect 339681 31767 339739 31773
rect 339770 31764 339776 31776
rect 339828 31764 339834 31816
rect 341150 31764 341156 31816
rect 341208 31764 341214 31816
rect 377122 31764 377128 31816
rect 377180 31764 377186 31816
rect 341168 31680 341196 31764
rect 377140 31680 377168 31764
rect 460106 31736 460112 31748
rect 460067 31708 460112 31736
rect 460106 31696 460112 31708
rect 460164 31696 460170 31748
rect 341150 31628 341156 31680
rect 341208 31628 341214 31680
rect 377122 31628 377128 31680
rect 377180 31628 377186 31680
rect 306653 31127 306711 31133
rect 306653 31093 306665 31127
rect 306699 31124 306711 31127
rect 306742 31124 306748 31136
rect 306699 31096 306748 31124
rect 306699 31093 306711 31096
rect 306653 31087 306711 31093
rect 306742 31084 306748 31096
rect 306800 31084 306806 31136
rect 253106 29180 253112 29232
rect 253164 29220 253170 29232
rect 257982 29220 257988 29232
rect 253164 29192 257988 29220
rect 253164 29180 253170 29192
rect 257982 29180 257988 29192
rect 258040 29180 258046 29232
rect 366818 29180 366824 29232
rect 366876 29220 366882 29232
rect 366876 29192 367048 29220
rect 366876 29180 366882 29192
rect 367020 29164 367048 29192
rect 437198 29180 437204 29232
rect 437256 29220 437262 29232
rect 437474 29220 437480 29232
rect 437256 29192 437480 29220
rect 437256 29180 437262 29192
rect 437474 29180 437480 29192
rect 437532 29180 437538 29232
rect 465258 29180 465264 29232
rect 465316 29220 465322 29232
rect 467926 29220 467932 29232
rect 465316 29192 467932 29220
rect 465316 29180 465322 29192
rect 467926 29180 467932 29192
rect 467984 29180 467990 29232
rect 367002 29112 367008 29164
rect 367060 29112 367066 29164
rect 417878 29112 417884 29164
rect 417936 29152 417942 29164
rect 418154 29152 418160 29164
rect 417936 29124 418160 29152
rect 417936 29112 417942 29124
rect 418154 29112 418160 29124
rect 418212 29112 418218 29164
rect 357710 29084 357716 29096
rect 357636 29056 357716 29084
rect 357636 29028 357664 29056
rect 357710 29044 357716 29056
rect 357768 29044 357774 29096
rect 492766 29044 492772 29096
rect 492824 29084 492830 29096
rect 502242 29084 502248 29096
rect 492824 29056 502248 29084
rect 492824 29044 492830 29056
rect 502242 29044 502248 29056
rect 502300 29044 502306 29096
rect 262674 28976 262680 29028
rect 262732 29016 262738 29028
rect 262766 29016 262772 29028
rect 262732 28988 262772 29016
rect 262732 28976 262738 28988
rect 262766 28976 262772 28988
rect 262824 28976 262830 29028
rect 265158 28976 265164 29028
rect 265216 29016 265222 29028
rect 265250 29016 265256 29028
rect 265216 28988 265256 29016
rect 265216 28976 265222 28988
rect 265250 28976 265256 28988
rect 265308 28976 265314 29028
rect 267826 28976 267832 29028
rect 267884 29016 267890 29028
rect 267918 29016 267924 29028
rect 267884 28988 267924 29016
rect 267884 28976 267890 28988
rect 267918 28976 267924 28988
rect 267976 28976 267982 29028
rect 281718 29016 281724 29028
rect 281679 28988 281724 29016
rect 281718 28976 281724 28988
rect 281776 28976 281782 29028
rect 301130 28976 301136 29028
rect 301188 29016 301194 29028
rect 301222 29016 301228 29028
rect 301188 28988 301228 29016
rect 301188 28976 301194 28988
rect 301222 28976 301228 28988
rect 301280 28976 301286 29028
rect 339678 29016 339684 29028
rect 339639 28988 339684 29016
rect 339678 28976 339684 28988
rect 339736 28976 339742 29028
rect 357618 28976 357624 29028
rect 357676 28976 357682 29028
rect 375742 28976 375748 29028
rect 375800 29016 375806 29028
rect 375834 29016 375840 29028
rect 375800 28988 375840 29016
rect 375800 28976 375806 28988
rect 375834 28976 375840 28988
rect 375892 28976 375898 29028
rect 284570 28908 284576 28960
rect 284628 28948 284634 28960
rect 284754 28948 284760 28960
rect 284628 28920 284760 28948
rect 284628 28908 284634 28920
rect 284754 28908 284760 28920
rect 284812 28908 284818 28960
rect 306282 28908 306288 28960
rect 306340 28948 306346 28960
rect 314562 28948 314568 28960
rect 306340 28920 314568 28948
rect 306340 28908 306346 28920
rect 314562 28908 314568 28920
rect 314620 28908 314626 28960
rect 323302 28908 323308 28960
rect 323360 28948 323366 28960
rect 323394 28948 323400 28960
rect 323360 28920 323400 28948
rect 323360 28908 323366 28920
rect 323394 28908 323400 28920
rect 323452 28908 323458 28960
rect 324590 28908 324596 28960
rect 324648 28948 324654 28960
rect 324682 28948 324688 28960
rect 324648 28920 324688 28948
rect 324648 28908 324654 28920
rect 324682 28908 324688 28920
rect 324740 28908 324746 28960
rect 325878 28908 325884 28960
rect 325936 28948 325942 28960
rect 325970 28948 325976 28960
rect 325936 28920 325976 28948
rect 325936 28908 325942 28920
rect 325970 28908 325976 28920
rect 326028 28908 326034 28960
rect 295610 27724 295616 27736
rect 295536 27696 295616 27724
rect 295536 27668 295564 27696
rect 295610 27684 295616 27696
rect 295668 27684 295674 27736
rect 389266 27684 389272 27736
rect 389324 27724 389330 27736
rect 389358 27724 389364 27736
rect 389324 27696 389364 27724
rect 389324 27684 389330 27696
rect 389358 27684 389364 27696
rect 389416 27684 389422 27736
rect 232225 27659 232283 27665
rect 232225 27625 232237 27659
rect 232271 27656 232283 27659
rect 232314 27656 232320 27668
rect 232271 27628 232320 27656
rect 232271 27625 232283 27628
rect 232225 27619 232283 27625
rect 232314 27616 232320 27628
rect 232372 27616 232378 27668
rect 291562 27616 291568 27668
rect 291620 27656 291626 27668
rect 291654 27656 291660 27668
rect 291620 27628 291660 27656
rect 291620 27616 291626 27628
rect 291654 27616 291660 27628
rect 291712 27616 291718 27668
rect 295518 27616 295524 27668
rect 295576 27616 295582 27668
rect 393593 27659 393651 27665
rect 393593 27625 393605 27659
rect 393639 27656 393651 27659
rect 393682 27656 393688 27668
rect 393639 27628 393688 27656
rect 393639 27625 393651 27628
rect 393593 27619 393651 27625
rect 393682 27616 393688 27628
rect 393740 27616 393746 27668
rect 230750 27588 230756 27600
rect 230711 27560 230756 27588
rect 230750 27548 230756 27560
rect 230808 27548 230814 27600
rect 265250 27588 265256 27600
rect 265211 27560 265256 27588
rect 265250 27548 265256 27560
rect 265308 27548 265314 27600
rect 302510 27548 302516 27600
rect 302568 27588 302574 27600
rect 302602 27588 302608 27600
rect 302568 27560 302608 27588
rect 302568 27548 302574 27560
rect 302602 27548 302608 27560
rect 302660 27548 302666 27600
rect 366821 27591 366879 27597
rect 366821 27557 366833 27591
rect 366867 27588 366879 27591
rect 367002 27588 367008 27600
rect 366867 27560 367008 27588
rect 366867 27557 366879 27560
rect 366821 27551 366879 27557
rect 367002 27548 367008 27560
rect 367060 27548 367066 27600
rect 375834 27588 375840 27600
rect 375795 27560 375840 27588
rect 375834 27548 375840 27560
rect 375892 27548 375898 27600
rect 247218 26364 247224 26376
rect 247179 26336 247224 26364
rect 247218 26324 247224 26336
rect 247276 26324 247282 26376
rect 259546 26364 259552 26376
rect 259507 26336 259552 26364
rect 259546 26324 259552 26336
rect 259604 26324 259610 26376
rect 306650 26364 306656 26376
rect 306611 26336 306656 26364
rect 306650 26324 306656 26336
rect 306708 26324 306714 26376
rect 250073 26299 250131 26305
rect 250073 26265 250085 26299
rect 250119 26296 250131 26299
rect 250162 26296 250168 26308
rect 250119 26268 250168 26296
rect 250119 26265 250131 26268
rect 250073 26259 250131 26265
rect 250162 26256 250168 26268
rect 250220 26256 250226 26308
rect 270770 26296 270776 26308
rect 270731 26268 270776 26296
rect 270770 26256 270776 26268
rect 270828 26256 270834 26308
rect 303982 26296 303988 26308
rect 303943 26268 303988 26296
rect 303982 26256 303988 26268
rect 304040 26256 304046 26308
rect 329926 26256 329932 26308
rect 329984 26296 329990 26308
rect 330202 26296 330208 26308
rect 329984 26268 330208 26296
rect 329984 26256 329990 26268
rect 330202 26256 330208 26268
rect 330260 26256 330266 26308
rect 245841 26231 245899 26237
rect 245841 26197 245853 26231
rect 245887 26228 245899 26231
rect 245930 26228 245936 26240
rect 245887 26200 245936 26228
rect 245887 26197 245899 26200
rect 245841 26191 245899 26197
rect 245930 26188 245936 26200
rect 245988 26188 245994 26240
rect 247129 26231 247187 26237
rect 247129 26197 247141 26231
rect 247175 26228 247187 26231
rect 247218 26228 247224 26240
rect 247175 26200 247224 26228
rect 247175 26197 247187 26200
rect 247129 26191 247187 26197
rect 247218 26188 247224 26200
rect 247276 26188 247282 26240
rect 259546 26228 259552 26240
rect 259507 26200 259552 26228
rect 259546 26188 259552 26200
rect 259604 26188 259610 26240
rect 272061 26231 272119 26237
rect 272061 26197 272073 26231
rect 272107 26228 272119 26231
rect 272242 26228 272248 26240
rect 272107 26200 272248 26228
rect 272107 26197 272119 26200
rect 272061 26191 272119 26197
rect 272242 26188 272248 26200
rect 272300 26188 272306 26240
rect 291565 26231 291623 26237
rect 291565 26197 291577 26231
rect 291611 26228 291623 26231
rect 291654 26228 291660 26240
rect 291611 26200 291660 26228
rect 291611 26197 291623 26200
rect 291565 26191 291623 26197
rect 291654 26188 291660 26200
rect 291712 26188 291718 26240
rect 310882 26228 310888 26240
rect 310843 26200 310888 26228
rect 310882 26188 310888 26200
rect 310940 26188 310946 26240
rect 331398 26228 331404 26240
rect 331359 26200 331404 26228
rect 331398 26188 331404 26200
rect 331456 26188 331462 26240
rect 389358 26228 389364 26240
rect 389319 26200 389364 26228
rect 389358 26188 389364 26200
rect 389416 26188 389422 26240
rect 329926 25848 329932 25900
rect 329984 25888 329990 25900
rect 330205 25891 330263 25897
rect 330205 25888 330217 25891
rect 329984 25860 330217 25888
rect 329984 25848 329990 25860
rect 330205 25857 330217 25860
rect 330251 25857 330263 25891
rect 330205 25851 330263 25857
rect 303982 24868 303988 24880
rect 303943 24840 303988 24868
rect 303982 24828 303988 24840
rect 304040 24828 304046 24880
rect 232133 22763 232191 22769
rect 232133 22729 232145 22763
rect 232179 22760 232191 22763
rect 232406 22760 232412 22772
rect 232179 22732 232412 22760
rect 232179 22729 232191 22732
rect 232133 22723 232191 22729
rect 232406 22720 232412 22732
rect 232464 22720 232470 22772
rect 267737 22627 267795 22633
rect 267737 22593 267749 22627
rect 267783 22624 267795 22627
rect 267826 22624 267832 22636
rect 267783 22596 267832 22624
rect 267783 22593 267795 22596
rect 267737 22587 267795 22593
rect 267826 22584 267832 22596
rect 267884 22584 267890 22636
rect 244185 22151 244243 22157
rect 244185 22117 244197 22151
rect 244231 22148 244243 22151
rect 244458 22148 244464 22160
rect 244231 22120 244464 22148
rect 244231 22117 244243 22120
rect 244185 22111 244243 22117
rect 244458 22108 244464 22120
rect 244516 22108 244522 22160
rect 249981 22151 250039 22157
rect 249981 22117 249993 22151
rect 250027 22148 250039 22151
rect 250162 22148 250168 22160
rect 250027 22120 250168 22148
rect 250027 22117 250039 22120
rect 249981 22111 250039 22117
rect 250162 22108 250168 22120
rect 250220 22108 250226 22160
rect 269850 22108 269856 22160
rect 269908 22148 269914 22160
rect 270678 22148 270684 22160
rect 269908 22120 270684 22148
rect 269908 22108 269914 22120
rect 270678 22108 270684 22120
rect 270736 22108 270742 22160
rect 377122 22108 377128 22160
rect 377180 22108 377186 22160
rect 377140 22024 377168 22108
rect 377122 21972 377128 22024
rect 377180 21972 377186 22024
rect 460106 21972 460112 22024
rect 460164 22012 460170 22024
rect 460382 22012 460388 22024
rect 460164 21984 460388 22012
rect 460164 21972 460170 21984
rect 460382 21972 460388 21984
rect 460440 21972 460446 22024
rect 375834 20856 375840 20868
rect 375795 20828 375840 20856
rect 375834 20816 375840 20828
rect 375892 20816 375898 20868
rect 266722 19428 266728 19440
rect 266648 19400 266728 19428
rect 251358 19320 251364 19372
rect 251416 19360 251422 19372
rect 251542 19360 251548 19372
rect 251416 19332 251548 19360
rect 251416 19320 251422 19332
rect 251542 19320 251548 19332
rect 251600 19320 251606 19372
rect 266648 19304 266676 19400
rect 266722 19388 266728 19400
rect 266780 19388 266786 19440
rect 281718 19428 281724 19440
rect 281644 19400 281724 19428
rect 281644 19372 281672 19400
rect 281718 19388 281724 19400
rect 281776 19388 281782 19440
rect 281626 19320 281632 19372
rect 281684 19320 281690 19372
rect 339678 19320 339684 19372
rect 339736 19360 339742 19372
rect 339770 19360 339776 19372
rect 339736 19332 339776 19360
rect 339736 19320 339742 19332
rect 339770 19320 339776 19332
rect 339828 19320 339834 19372
rect 341242 19320 341248 19372
rect 341300 19360 341306 19372
rect 341334 19360 341340 19372
rect 341300 19332 341340 19360
rect 341300 19320 341306 19332
rect 341334 19320 341340 19332
rect 341392 19320 341398 19372
rect 266630 19252 266636 19304
rect 266688 19252 266694 19304
rect 295518 19292 295524 19304
rect 295479 19264 295524 19292
rect 295518 19252 295524 19264
rect 295576 19252 295582 19304
rect 339681 19227 339739 19233
rect 339681 19193 339693 19227
rect 339727 19224 339739 19227
rect 339770 19224 339776 19236
rect 339727 19196 339776 19224
rect 339727 19193 339739 19196
rect 339681 19187 339739 19193
rect 339770 19184 339776 19196
rect 339828 19184 339834 19236
rect 265253 18071 265311 18077
rect 265253 18037 265265 18071
rect 265299 18037 265311 18071
rect 265253 18031 265311 18037
rect 230750 18000 230756 18012
rect 230711 17972 230756 18000
rect 230750 17960 230756 17972
rect 230808 17960 230814 18012
rect 259546 17932 259552 17944
rect 259507 17904 259552 17932
rect 259546 17892 259552 17904
rect 259604 17892 259610 17944
rect 264974 17892 264980 17944
rect 265032 17932 265038 17944
rect 265268 17932 265296 18031
rect 393682 18028 393688 18080
rect 393740 18028 393746 18080
rect 393700 17944 393728 18028
rect 273438 17932 273444 17944
rect 265032 17904 265296 17932
rect 273399 17904 273444 17932
rect 265032 17892 265038 17904
rect 273438 17892 273444 17904
rect 273496 17892 273502 17944
rect 393682 17892 393688 17944
rect 393740 17892 393746 17944
rect 299382 16940 299388 16992
rect 299440 16980 299446 16992
rect 311158 16980 311164 16992
rect 299440 16952 311164 16980
rect 299440 16940 299446 16952
rect 311158 16940 311164 16952
rect 311216 16940 311222 16992
rect 417878 16736 417884 16788
rect 417936 16776 417942 16788
rect 418154 16776 418160 16788
rect 417936 16748 418160 16776
rect 417936 16736 417942 16748
rect 418154 16736 418160 16748
rect 418212 16736 418218 16788
rect 437198 16736 437204 16788
rect 437256 16776 437262 16788
rect 437474 16776 437480 16788
rect 437256 16748 437480 16776
rect 437256 16736 437262 16748
rect 437474 16736 437480 16748
rect 437532 16736 437538 16788
rect 463786 16668 463792 16720
rect 463844 16708 463850 16720
rect 466546 16708 466552 16720
rect 463844 16680 466552 16708
rect 463844 16668 463850 16680
rect 466546 16668 466552 16680
rect 466604 16668 466610 16720
rect 244182 16640 244188 16652
rect 244143 16612 244188 16640
rect 244182 16600 244188 16612
rect 244240 16600 244246 16652
rect 245838 16640 245844 16652
rect 245799 16612 245844 16640
rect 245838 16600 245844 16612
rect 245896 16600 245902 16652
rect 249978 16640 249984 16652
rect 249939 16612 249984 16640
rect 249978 16600 249984 16612
rect 250036 16600 250042 16652
rect 291562 16640 291568 16652
rect 291523 16612 291568 16640
rect 291562 16600 291568 16612
rect 291620 16600 291626 16652
rect 310882 16640 310888 16652
rect 310843 16612 310888 16640
rect 310882 16600 310888 16612
rect 310940 16600 310946 16652
rect 389358 16640 389364 16652
rect 389319 16612 389364 16640
rect 389358 16600 389364 16612
rect 389416 16600 389422 16652
rect 306834 15172 306840 15224
rect 306892 15212 306898 15224
rect 307018 15212 307024 15224
rect 306892 15184 307024 15212
rect 306892 15172 306898 15184
rect 307018 15172 307024 15184
rect 307076 15172 307082 15224
rect 110322 15104 110328 15156
rect 110380 15144 110386 15156
rect 274726 15144 274732 15156
rect 110380 15116 274732 15144
rect 110380 15104 110386 15116
rect 274726 15104 274732 15116
rect 274784 15104 274790 15156
rect 107470 15036 107476 15088
rect 107528 15076 107534 15088
rect 273346 15076 273352 15088
rect 107528 15048 273352 15076
rect 107528 15036 107534 15048
rect 273346 15036 273352 15048
rect 273404 15036 273410 15088
rect 103422 14968 103428 15020
rect 103480 15008 103486 15020
rect 271966 15008 271972 15020
rect 103480 14980 271972 15008
rect 103480 14968 103486 14980
rect 271966 14968 271972 14980
rect 272024 14968 272030 15020
rect 99282 14900 99288 14952
rect 99340 14940 99346 14952
rect 270586 14940 270592 14952
rect 99340 14912 270592 14940
rect 99340 14900 99346 14912
rect 270586 14900 270592 14912
rect 270644 14900 270650 14952
rect 96522 14832 96528 14884
rect 96580 14872 96586 14884
rect 269206 14872 269212 14884
rect 96580 14844 269212 14872
rect 96580 14832 96586 14844
rect 269206 14832 269212 14844
rect 269264 14832 269270 14884
rect 92382 14764 92388 14816
rect 92440 14804 92446 14816
rect 266446 14804 266452 14816
rect 92440 14776 266452 14804
rect 92440 14764 92446 14776
rect 266446 14764 266452 14776
rect 266504 14764 266510 14816
rect 89622 14696 89628 14748
rect 89680 14736 89686 14748
rect 265066 14736 265072 14748
rect 89680 14708 265072 14736
rect 89680 14696 89686 14708
rect 265066 14696 265072 14708
rect 265124 14696 265130 14748
rect 85482 14628 85488 14680
rect 85540 14668 85546 14680
rect 263686 14668 263692 14680
rect 85540 14640 263692 14668
rect 85540 14628 85546 14640
rect 263686 14628 263692 14640
rect 263744 14628 263750 14680
rect 82722 14560 82728 14612
rect 82780 14600 82786 14612
rect 262582 14600 262588 14612
rect 82780 14572 262588 14600
rect 82780 14560 82786 14572
rect 262582 14560 262588 14572
rect 262640 14560 262646 14612
rect 78582 14492 78588 14544
rect 78640 14532 78646 14544
rect 260926 14532 260932 14544
rect 78640 14504 260932 14532
rect 78640 14492 78646 14504
rect 260926 14492 260932 14504
rect 260984 14492 260990 14544
rect 74442 14424 74448 14476
rect 74500 14464 74506 14476
rect 259546 14464 259552 14476
rect 74500 14436 259552 14464
rect 74500 14424 74506 14436
rect 259546 14424 259552 14436
rect 259604 14424 259610 14476
rect 114462 14356 114468 14408
rect 114520 14396 114526 14408
rect 276106 14396 276112 14408
rect 114520 14368 276112 14396
rect 114520 14356 114526 14368
rect 276106 14356 276112 14368
rect 276164 14356 276170 14408
rect 117222 14288 117228 14340
rect 117280 14328 117286 14340
rect 277670 14328 277676 14340
rect 117280 14300 277676 14328
rect 117280 14288 117286 14300
rect 277670 14288 277676 14300
rect 277728 14288 277734 14340
rect 121362 14220 121368 14272
rect 121420 14260 121426 14272
rect 278774 14260 278780 14272
rect 121420 14232 278780 14260
rect 121420 14220 121426 14232
rect 278774 14220 278780 14232
rect 278832 14220 278838 14272
rect 125410 14152 125416 14204
rect 125468 14192 125474 14204
rect 280246 14192 280252 14204
rect 125468 14164 280252 14192
rect 125468 14152 125474 14164
rect 280246 14152 280252 14164
rect 280304 14152 280310 14204
rect 232130 14124 232136 14136
rect 232091 14096 232136 14124
rect 232130 14084 232136 14096
rect 232188 14084 232194 14136
rect 183462 13744 183468 13796
rect 183520 13784 183526 13796
rect 303982 13784 303988 13796
rect 183520 13756 303988 13784
rect 183520 13744 183526 13756
rect 303982 13744 303988 13756
rect 304040 13744 304046 13796
rect 186222 13676 186228 13728
rect 186280 13716 186286 13728
rect 306558 13716 306564 13728
rect 186280 13688 306564 13716
rect 186280 13676 186286 13688
rect 306558 13676 306564 13688
rect 306616 13676 306622 13728
rect 179322 13608 179328 13660
rect 179380 13648 179386 13660
rect 302510 13648 302516 13660
rect 179380 13620 302516 13648
rect 179380 13608 179386 13620
rect 302510 13608 302516 13620
rect 302568 13608 302574 13660
rect 176562 13540 176568 13592
rect 176620 13580 176626 13592
rect 301038 13580 301044 13592
rect 176620 13552 301044 13580
rect 176620 13540 176626 13552
rect 301038 13540 301044 13552
rect 301096 13540 301102 13592
rect 172422 13472 172428 13524
rect 172480 13512 172486 13524
rect 299750 13512 299756 13524
rect 172480 13484 299756 13512
rect 172480 13472 172486 13484
rect 299750 13472 299756 13484
rect 299808 13472 299814 13524
rect 168282 13404 168288 13456
rect 168340 13444 168346 13456
rect 298278 13444 298284 13456
rect 168340 13416 298284 13444
rect 168340 13404 168346 13416
rect 298278 13404 298284 13416
rect 298336 13404 298342 13456
rect 165522 13336 165528 13388
rect 165580 13376 165586 13388
rect 296898 13376 296904 13388
rect 165580 13348 296904 13376
rect 165580 13336 165586 13348
rect 296898 13336 296904 13348
rect 296956 13336 296962 13388
rect 160002 13268 160008 13320
rect 160060 13308 160066 13320
rect 294414 13308 294420 13320
rect 160060 13280 294420 13308
rect 160060 13268 160066 13280
rect 294414 13268 294420 13280
rect 294472 13268 294478 13320
rect 155862 13200 155868 13252
rect 155920 13240 155926 13252
rect 292758 13240 292764 13252
rect 155920 13212 292764 13240
rect 155920 13200 155926 13212
rect 292758 13200 292764 13212
rect 292816 13200 292822 13252
rect 71682 13132 71688 13184
rect 71740 13172 71746 13184
rect 258166 13172 258172 13184
rect 71740 13144 258172 13172
rect 71740 13132 71746 13144
rect 258166 13132 258172 13144
rect 258224 13132 258230 13184
rect 31662 13064 31668 13116
rect 31720 13104 31726 13116
rect 241606 13104 241612 13116
rect 31720 13076 241612 13104
rect 31720 13064 31726 13076
rect 241606 13064 241612 13076
rect 241664 13064 241670 13116
rect 190362 12996 190368 13048
rect 190420 13036 190426 13048
rect 307938 13036 307944 13048
rect 190420 13008 307944 13036
rect 190420 12996 190426 13008
rect 307938 12996 307944 13008
rect 307996 12996 308002 13048
rect 206922 12928 206928 12980
rect 206980 12968 206986 12980
rect 314838 12968 314844 12980
rect 206980 12940 314844 12968
rect 206980 12928 206986 12940
rect 314838 12928 314844 12940
rect 314896 12928 314902 12980
rect 211062 12860 211068 12912
rect 211120 12900 211126 12912
rect 316218 12900 316224 12912
rect 211120 12872 316224 12900
rect 211120 12860 211126 12872
rect 316218 12860 316224 12872
rect 316276 12860 316282 12912
rect 213822 12792 213828 12844
rect 213880 12832 213886 12844
rect 317598 12832 317604 12844
rect 213880 12804 317604 12832
rect 213880 12792 213886 12804
rect 317598 12792 317604 12804
rect 317656 12792 317662 12844
rect 217962 12724 217968 12776
rect 218020 12764 218026 12776
rect 318978 12764 318984 12776
rect 218020 12736 318984 12764
rect 218020 12724 218026 12736
rect 318978 12724 318984 12736
rect 319036 12724 319042 12776
rect 220722 12656 220728 12708
rect 220780 12696 220786 12708
rect 320266 12696 320272 12708
rect 220780 12668 320272 12696
rect 220780 12656 220786 12668
rect 320266 12656 320272 12668
rect 320324 12656 320330 12708
rect 224862 12588 224868 12640
rect 224920 12628 224926 12640
rect 321738 12628 321744 12640
rect 224920 12600 321744 12628
rect 224920 12588 224926 12600
rect 321738 12588 321744 12600
rect 321796 12588 321802 12640
rect 229002 12520 229008 12572
rect 229060 12560 229066 12572
rect 323118 12560 323124 12572
rect 229060 12532 323124 12560
rect 229060 12520 229066 12532
rect 323118 12520 323124 12532
rect 323176 12520 323182 12572
rect 230661 12495 230719 12501
rect 230661 12461 230673 12495
rect 230707 12492 230719 12495
rect 230750 12492 230756 12504
rect 230707 12464 230756 12492
rect 230707 12461 230719 12464
rect 230661 12455 230719 12461
rect 230750 12452 230756 12464
rect 230808 12452 230814 12504
rect 366910 12452 366916 12504
rect 366968 12452 366974 12504
rect 173802 12384 173808 12436
rect 173860 12424 173866 12436
rect 300946 12424 300952 12436
rect 173860 12396 300952 12424
rect 173860 12384 173866 12396
rect 300946 12384 300952 12396
rect 301004 12384 301010 12436
rect 366928 12368 366956 12452
rect 169662 12316 169668 12368
rect 169720 12356 169726 12368
rect 299566 12356 299572 12368
rect 169720 12328 299572 12356
rect 169720 12316 169726 12328
rect 299566 12316 299572 12328
rect 299624 12316 299630 12368
rect 366910 12316 366916 12368
rect 366968 12316 366974 12368
rect 166902 12248 166908 12300
rect 166960 12288 166966 12300
rect 298186 12288 298192 12300
rect 166960 12260 298192 12288
rect 166960 12248 166966 12260
rect 298186 12248 298192 12260
rect 298244 12248 298250 12300
rect 162762 12180 162768 12232
rect 162820 12220 162826 12232
rect 295521 12223 295579 12229
rect 295521 12220 295533 12223
rect 162820 12192 295533 12220
rect 162820 12180 162826 12192
rect 295521 12189 295533 12192
rect 295567 12189 295579 12223
rect 295521 12183 295579 12189
rect 151722 12112 151728 12164
rect 151780 12152 151786 12164
rect 291562 12152 291568 12164
rect 151780 12124 291568 12152
rect 151780 12112 151786 12124
rect 291562 12112 291568 12124
rect 291620 12112 291626 12164
rect 148962 12044 148968 12096
rect 149020 12084 149026 12096
rect 289998 12084 290004 12096
rect 149020 12056 290004 12084
rect 149020 12044 149026 12056
rect 289998 12044 290004 12056
rect 290056 12044 290062 12096
rect 144822 11976 144828 12028
rect 144880 12016 144886 12028
rect 288894 12016 288900 12028
rect 144880 11988 288900 12016
rect 144880 11976 144886 11988
rect 288894 11976 288900 11988
rect 288952 11976 288958 12028
rect 142062 11908 142068 11960
rect 142120 11948 142126 11960
rect 287330 11948 287336 11960
rect 142120 11920 287336 11948
rect 142120 11908 142126 11920
rect 287330 11908 287336 11920
rect 287388 11908 287394 11960
rect 128262 11840 128268 11892
rect 128320 11880 128326 11892
rect 281626 11880 281632 11892
rect 128320 11852 281632 11880
rect 128320 11840 128326 11852
rect 281626 11840 281632 11852
rect 281684 11840 281690 11892
rect 126882 11772 126888 11824
rect 126940 11812 126946 11824
rect 281534 11812 281540 11824
rect 126940 11784 281540 11812
rect 126940 11772 126946 11784
rect 281534 11772 281540 11784
rect 281592 11772 281598 11824
rect 23382 11704 23388 11756
rect 23440 11744 23446 11756
rect 238938 11744 238944 11756
rect 23440 11716 238944 11744
rect 23440 11704 23446 11716
rect 238938 11704 238944 11716
rect 238996 11704 239002 11756
rect 468846 11704 468852 11756
rect 468904 11744 468910 11756
rect 469122 11744 469128 11756
rect 468904 11716 469128 11744
rect 468904 11704 468910 11716
rect 469122 11704 469128 11716
rect 469180 11704 469186 11756
rect 176470 11636 176476 11688
rect 176528 11676 176534 11688
rect 302326 11676 302332 11688
rect 176528 11648 302332 11676
rect 176528 11636 176534 11648
rect 302326 11636 302332 11648
rect 302384 11636 302390 11688
rect 180702 11568 180708 11620
rect 180760 11608 180766 11620
rect 303706 11608 303712 11620
rect 180760 11580 303712 11608
rect 180760 11568 180766 11580
rect 303706 11568 303712 11580
rect 303764 11568 303770 11620
rect 184842 11500 184848 11552
rect 184900 11540 184906 11552
rect 305086 11540 305092 11552
rect 184900 11512 305092 11540
rect 184900 11500 184906 11512
rect 305086 11500 305092 11512
rect 305144 11500 305150 11552
rect 187602 11432 187608 11484
rect 187660 11472 187666 11484
rect 306466 11472 306472 11484
rect 187660 11444 306472 11472
rect 187660 11432 187666 11444
rect 306466 11432 306472 11444
rect 306524 11432 306530 11484
rect 191742 11364 191748 11416
rect 191800 11404 191806 11416
rect 308030 11404 308036 11416
rect 191800 11376 308036 11404
rect 191800 11364 191806 11376
rect 308030 11364 308036 11376
rect 308088 11364 308094 11416
rect 194502 11296 194508 11348
rect 194560 11336 194566 11348
rect 309410 11336 309416 11348
rect 194560 11308 309416 11336
rect 194560 11296 194566 11308
rect 309410 11296 309416 11308
rect 309468 11296 309474 11348
rect 198642 11228 198648 11280
rect 198700 11268 198706 11280
rect 310882 11268 310888 11280
rect 198700 11240 310888 11268
rect 198700 11228 198706 11240
rect 310882 11228 310888 11240
rect 310940 11228 310946 11280
rect 230658 11200 230664 11212
rect 230619 11172 230664 11200
rect 230658 11160 230664 11172
rect 230716 11160 230722 11212
rect 113082 10956 113088 11008
rect 113140 10996 113146 11008
rect 276014 10996 276020 11008
rect 113140 10968 276020 10996
rect 113140 10956 113146 10968
rect 276014 10956 276020 10968
rect 276072 10956 276078 11008
rect 108942 10888 108948 10940
rect 109000 10928 109006 10940
rect 273441 10931 273499 10937
rect 273441 10928 273453 10931
rect 109000 10900 273453 10928
rect 109000 10888 109006 10900
rect 273441 10897 273453 10900
rect 273487 10897 273499 10931
rect 273441 10891 273499 10897
rect 106182 10820 106188 10872
rect 106240 10860 106246 10872
rect 272061 10863 272119 10869
rect 272061 10860 272073 10863
rect 106240 10832 272073 10860
rect 106240 10820 106246 10832
rect 272061 10829 272073 10832
rect 272107 10829 272119 10863
rect 272061 10823 272119 10829
rect 102042 10752 102048 10804
rect 102100 10792 102106 10804
rect 269850 10792 269856 10804
rect 102100 10764 269856 10792
rect 102100 10752 102106 10764
rect 269850 10752 269856 10764
rect 269908 10752 269914 10804
rect 99190 10684 99196 10736
rect 99248 10724 99254 10736
rect 269298 10724 269304 10736
rect 99248 10696 269304 10724
rect 99248 10684 99254 10696
rect 269298 10684 269304 10696
rect 269356 10684 269362 10736
rect 95142 10616 95148 10668
rect 95200 10656 95206 10668
rect 267737 10659 267795 10665
rect 267737 10656 267749 10659
rect 95200 10628 267749 10656
rect 95200 10616 95206 10628
rect 267737 10625 267749 10628
rect 267783 10625 267795 10659
rect 267737 10619 267795 10625
rect 91002 10548 91008 10600
rect 91060 10588 91066 10600
rect 266630 10588 266636 10600
rect 91060 10560 266636 10588
rect 91060 10548 91066 10560
rect 266630 10548 266636 10560
rect 266688 10548 266694 10600
rect 64782 10480 64788 10532
rect 64840 10520 64846 10532
rect 255590 10520 255596 10532
rect 64840 10492 255596 10520
rect 64840 10480 64846 10492
rect 255590 10480 255596 10492
rect 255648 10480 255654 10532
rect 60642 10412 60648 10464
rect 60700 10452 60706 10464
rect 254026 10452 254032 10464
rect 60700 10424 254032 10452
rect 60700 10412 60706 10424
rect 254026 10412 254032 10424
rect 254084 10412 254090 10464
rect 56502 10344 56508 10396
rect 56560 10384 56566 10396
rect 252646 10384 252652 10396
rect 56560 10356 252652 10384
rect 56560 10344 56566 10356
rect 252646 10344 252652 10356
rect 252704 10344 252710 10396
rect 53742 10276 53748 10328
rect 53800 10316 53806 10328
rect 251266 10316 251272 10328
rect 53800 10288 251272 10316
rect 53800 10276 53806 10288
rect 251266 10276 251272 10288
rect 251324 10276 251330 10328
rect 117130 10208 117136 10260
rect 117188 10248 117194 10260
rect 277578 10248 277584 10260
rect 117188 10220 277584 10248
rect 117188 10208 117194 10220
rect 277578 10208 277584 10220
rect 277636 10208 277642 10260
rect 119982 10140 119988 10192
rect 120040 10180 120046 10192
rect 278958 10180 278964 10192
rect 120040 10152 278964 10180
rect 120040 10140 120046 10152
rect 278958 10140 278964 10152
rect 279016 10140 279022 10192
rect 124122 10072 124128 10124
rect 124180 10112 124186 10124
rect 280338 10112 280344 10124
rect 124180 10084 280344 10112
rect 124180 10072 124186 10084
rect 280338 10072 280344 10084
rect 280396 10072 280402 10124
rect 143442 10004 143448 10056
rect 143500 10044 143506 10056
rect 288526 10044 288532 10056
rect 143500 10016 288532 10044
rect 143500 10004 143506 10016
rect 288526 10004 288532 10016
rect 288584 10004 288590 10056
rect 147582 9936 147588 9988
rect 147640 9976 147646 9988
rect 289814 9976 289820 9988
rect 147640 9948 289820 9976
rect 147640 9936 147646 9948
rect 289814 9936 289820 9948
rect 289872 9936 289878 9988
rect 151630 9868 151636 9920
rect 151688 9908 151694 9920
rect 291286 9908 291292 9920
rect 151688 9880 291292 9908
rect 151688 9868 151694 9880
rect 291286 9868 291292 9880
rect 291344 9868 291350 9920
rect 154482 9800 154488 9852
rect 154540 9840 154546 9852
rect 292850 9840 292856 9852
rect 154540 9812 292856 9840
rect 154540 9800 154546 9812
rect 292850 9800 292856 9812
rect 292908 9800 292914 9852
rect 158622 9732 158628 9784
rect 158680 9772 158686 9784
rect 294046 9772 294052 9784
rect 158680 9744 294052 9772
rect 158680 9732 158686 9744
rect 294046 9732 294052 9744
rect 294104 9732 294110 9784
rect 161382 9664 161388 9716
rect 161440 9704 161446 9716
rect 295426 9704 295432 9716
rect 161440 9676 295432 9704
rect 161440 9664 161446 9676
rect 295426 9664 295432 9676
rect 295484 9664 295490 9716
rect 330202 9704 330208 9716
rect 330163 9676 330208 9704
rect 330202 9664 330208 9676
rect 330260 9664 330266 9716
rect 331398 9704 331404 9716
rect 331359 9676 331404 9704
rect 331398 9664 331404 9676
rect 331456 9664 331462 9716
rect 339678 9704 339684 9716
rect 339639 9676 339684 9704
rect 339678 9664 339684 9676
rect 339736 9664 339742 9716
rect 366818 9704 366824 9716
rect 366779 9676 366824 9704
rect 366818 9664 366824 9676
rect 366876 9664 366882 9716
rect 203886 9596 203892 9648
rect 203944 9636 203950 9648
rect 313366 9636 313372 9648
rect 203944 9608 313372 9636
rect 203944 9596 203950 9608
rect 313366 9596 313372 9608
rect 313424 9596 313430 9648
rect 200390 9528 200396 9580
rect 200448 9568 200454 9580
rect 311986 9568 311992 9580
rect 200448 9540 311992 9568
rect 200448 9528 200454 9540
rect 311986 9528 311992 9540
rect 312044 9528 312050 9580
rect 196802 9460 196808 9512
rect 196860 9500 196866 9512
rect 310606 9500 310612 9512
rect 196860 9472 310612 9500
rect 196860 9460 196866 9472
rect 310606 9460 310612 9472
rect 310664 9460 310670 9512
rect 193214 9392 193220 9444
rect 193272 9432 193278 9444
rect 309226 9432 309232 9444
rect 193272 9404 309232 9432
rect 193272 9392 193278 9404
rect 309226 9392 309232 9404
rect 309284 9392 309290 9444
rect 139670 9324 139676 9376
rect 139728 9364 139734 9376
rect 287146 9364 287152 9376
rect 139728 9336 287152 9364
rect 139728 9324 139734 9336
rect 287146 9324 287152 9336
rect 287204 9324 287210 9376
rect 136082 9256 136088 9308
rect 136140 9296 136146 9308
rect 285858 9296 285864 9308
rect 136140 9268 285864 9296
rect 136140 9256 136146 9268
rect 285858 9256 285864 9268
rect 285916 9256 285922 9308
rect 49326 9188 49332 9240
rect 49384 9228 49390 9240
rect 249886 9228 249892 9240
rect 49384 9200 249892 9228
rect 49384 9188 49390 9200
rect 249886 9188 249892 9200
rect 249944 9188 249950 9240
rect 253842 9188 253848 9240
rect 253900 9228 253906 9240
rect 334158 9228 334164 9240
rect 253900 9200 334164 9228
rect 253900 9188 253906 9200
rect 334158 9188 334164 9200
rect 334216 9188 334222 9240
rect 44542 9120 44548 9172
rect 44600 9160 44606 9172
rect 247129 9163 247187 9169
rect 247129 9160 247141 9163
rect 44600 9132 247141 9160
rect 44600 9120 44606 9132
rect 247129 9129 247141 9132
rect 247175 9129 247187 9163
rect 247129 9123 247187 9129
rect 250346 9120 250352 9172
rect 250404 9160 250410 9172
rect 332778 9160 332784 9172
rect 250404 9132 332784 9160
rect 250404 9120 250410 9132
rect 332778 9120 332784 9132
rect 332836 9120 332842 9172
rect 27890 9052 27896 9104
rect 27948 9092 27954 9104
rect 233878 9092 233884 9104
rect 27948 9064 233884 9092
rect 27948 9052 27954 9064
rect 233878 9052 233884 9064
rect 233936 9052 233942 9104
rect 243170 9052 243176 9104
rect 243228 9092 243234 9104
rect 330018 9092 330024 9104
rect 243228 9064 330024 9092
rect 243228 9052 243234 9064
rect 330018 9052 330024 9064
rect 330076 9052 330082 9104
rect 18322 8984 18328 9036
rect 18380 9024 18386 9036
rect 236178 9024 236184 9036
rect 18380 8996 236184 9024
rect 18380 8984 18386 8996
rect 236178 8984 236184 8996
rect 236236 8984 236242 9036
rect 239582 8984 239588 9036
rect 239640 9024 239646 9036
rect 328638 9024 328644 9036
rect 239640 8996 328644 9024
rect 239640 8984 239646 8996
rect 328638 8984 328644 8996
rect 328696 8984 328702 9036
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 234798 8956 234804 8968
rect 13688 8928 234804 8956
rect 13688 8916 13694 8928
rect 234798 8916 234804 8928
rect 234856 8916 234862 8968
rect 235994 8916 236000 8968
rect 236052 8956 236058 8968
rect 325970 8956 325976 8968
rect 236052 8928 325976 8956
rect 236052 8916 236058 8928
rect 325970 8916 325976 8928
rect 326028 8916 326034 8968
rect 207474 8848 207480 8900
rect 207532 8888 207538 8900
rect 314930 8888 314936 8900
rect 207532 8860 314936 8888
rect 207532 8848 207538 8860
rect 314930 8848 314936 8860
rect 314988 8848 314994 8900
rect 210970 8780 210976 8832
rect 211028 8820 211034 8832
rect 316126 8820 316132 8832
rect 211028 8792 316132 8820
rect 211028 8780 211034 8792
rect 316126 8780 316132 8792
rect 316184 8780 316190 8832
rect 214650 8712 214656 8764
rect 214708 8752 214714 8764
rect 317506 8752 317512 8764
rect 214708 8724 317512 8752
rect 214708 8712 214714 8724
rect 317506 8712 317512 8724
rect 317564 8712 317570 8764
rect 218146 8644 218152 8696
rect 218204 8684 218210 8696
rect 318886 8684 318892 8696
rect 218204 8656 318892 8684
rect 218204 8644 218210 8656
rect 318886 8644 318892 8656
rect 318944 8644 318950 8696
rect 221734 8576 221740 8628
rect 221792 8616 221798 8628
rect 320174 8616 320180 8628
rect 221792 8588 320180 8616
rect 221792 8576 221798 8588
rect 320174 8576 320180 8588
rect 320232 8576 320238 8628
rect 225322 8508 225328 8560
rect 225380 8548 225386 8560
rect 321646 8548 321652 8560
rect 225380 8520 321652 8548
rect 225380 8508 225386 8520
rect 321646 8508 321652 8520
rect 321704 8508 321710 8560
rect 228910 8440 228916 8492
rect 228968 8480 228974 8492
rect 323302 8480 323308 8492
rect 228968 8452 323308 8480
rect 228968 8440 228974 8452
rect 323302 8440 323308 8452
rect 323360 8440 323366 8492
rect 232498 8372 232504 8424
rect 232556 8412 232562 8424
rect 324590 8412 324596 8424
rect 232556 8384 324596 8412
rect 232556 8372 232562 8384
rect 324590 8372 324596 8384
rect 324648 8372 324654 8424
rect 246758 8304 246764 8356
rect 246816 8344 246822 8356
rect 331398 8344 331404 8356
rect 246816 8316 331404 8344
rect 246816 8304 246822 8316
rect 331398 8304 331404 8316
rect 331456 8304 331462 8356
rect 87322 8236 87328 8288
rect 87380 8276 87386 8288
rect 265158 8276 265164 8288
rect 87380 8248 265164 8276
rect 87380 8236 87386 8248
rect 265158 8236 265164 8248
rect 265216 8236 265222 8288
rect 270494 8236 270500 8288
rect 270552 8276 270558 8288
rect 340966 8276 340972 8288
rect 270552 8248 340972 8276
rect 270552 8236 270558 8248
rect 340966 8236 340972 8248
rect 341024 8236 341030 8288
rect 445478 8236 445484 8288
rect 445536 8276 445542 8288
rect 523862 8276 523868 8288
rect 445536 8248 523868 8276
rect 445536 8236 445542 8248
rect 523862 8236 523868 8248
rect 523920 8236 523926 8288
rect 83826 8168 83832 8220
rect 83884 8208 83890 8220
rect 263870 8208 263876 8220
rect 83884 8180 263876 8208
rect 83884 8168 83890 8180
rect 263870 8168 263876 8180
rect 263928 8168 263934 8220
rect 266998 8168 267004 8220
rect 267056 8208 267062 8220
rect 339586 8208 339592 8220
rect 267056 8180 339592 8208
rect 267056 8168 267062 8180
rect 339586 8168 339592 8180
rect 339644 8168 339650 8220
rect 446950 8168 446956 8220
rect 447008 8208 447014 8220
rect 527450 8208 527456 8220
rect 447008 8180 527456 8208
rect 447008 8168 447014 8180
rect 527450 8168 527456 8180
rect 527508 8168 527514 8220
rect 80238 8100 80244 8152
rect 80296 8140 80302 8152
rect 262398 8140 262404 8152
rect 80296 8112 262404 8140
rect 80296 8100 80302 8112
rect 262398 8100 262404 8112
rect 262456 8100 262462 8152
rect 263410 8100 263416 8152
rect 263468 8140 263474 8152
rect 338298 8140 338304 8152
rect 263468 8112 338304 8140
rect 263468 8100 263474 8112
rect 338298 8100 338304 8112
rect 338356 8100 338362 8152
rect 448238 8100 448244 8152
rect 448296 8140 448302 8152
rect 531038 8140 531044 8152
rect 448296 8112 531044 8140
rect 448296 8100 448302 8112
rect 531038 8100 531044 8112
rect 531096 8100 531102 8152
rect 40954 8032 40960 8084
rect 41012 8072 41018 8084
rect 245930 8072 245936 8084
rect 41012 8044 245936 8072
rect 41012 8032 41018 8044
rect 245930 8032 245936 8044
rect 245988 8032 245994 8084
rect 259822 8032 259828 8084
rect 259880 8072 259886 8084
rect 336918 8072 336924 8084
rect 259880 8044 336924 8072
rect 259880 8032 259886 8044
rect 336918 8032 336924 8044
rect 336976 8032 336982 8084
rect 450998 8032 451004 8084
rect 451056 8072 451062 8084
rect 534534 8072 534540 8084
rect 451056 8044 534540 8072
rect 451056 8032 451062 8044
rect 534534 8032 534540 8044
rect 534592 8032 534598 8084
rect 37366 7964 37372 8016
rect 37424 8004 37430 8016
rect 244274 8004 244280 8016
rect 37424 7976 244280 8004
rect 37424 7964 37430 7976
rect 244274 7964 244280 7976
rect 244332 7964 244338 8016
rect 256234 7964 256240 8016
rect 256292 8004 256298 8016
rect 334066 8004 334072 8016
rect 256292 7976 334072 8004
rect 256292 7964 256298 7976
rect 334066 7964 334072 7976
rect 334124 7964 334130 8016
rect 452470 7964 452476 8016
rect 452528 8004 452534 8016
rect 538122 8004 538128 8016
rect 452528 7976 538128 8004
rect 452528 7964 452534 7976
rect 538122 7964 538128 7976
rect 538180 7964 538186 8016
rect 33870 7896 33876 7948
rect 33928 7936 33934 7948
rect 242986 7936 242992 7948
rect 33928 7908 242992 7936
rect 33928 7896 33934 7908
rect 242986 7896 242992 7908
rect 243044 7896 243050 7948
rect 252646 7896 252652 7948
rect 252704 7936 252710 7948
rect 332686 7936 332692 7948
rect 252704 7908 332692 7936
rect 252704 7896 252710 7908
rect 332686 7896 332692 7908
rect 332744 7896 332750 7948
rect 453758 7896 453764 7948
rect 453816 7936 453822 7948
rect 541710 7936 541716 7948
rect 453816 7908 541716 7936
rect 453816 7896 453822 7908
rect 541710 7896 541716 7908
rect 541768 7896 541774 7948
rect 30282 7828 30288 7880
rect 30340 7868 30346 7880
rect 241790 7868 241796 7880
rect 30340 7840 241796 7868
rect 30340 7828 30346 7840
rect 241790 7828 241796 7840
rect 241848 7828 241854 7880
rect 249150 7828 249156 7880
rect 249208 7868 249214 7880
rect 331306 7868 331312 7880
rect 249208 7840 331312 7868
rect 249208 7828 249214 7840
rect 331306 7828 331312 7840
rect 331364 7828 331370 7880
rect 455230 7828 455236 7880
rect 455288 7868 455294 7880
rect 545298 7868 545304 7880
rect 455288 7840 545304 7868
rect 455288 7828 455294 7840
rect 545298 7828 545304 7840
rect 545356 7828 545362 7880
rect 26694 7760 26700 7812
rect 26752 7800 26758 7812
rect 240410 7800 240416 7812
rect 26752 7772 240416 7800
rect 26752 7760 26758 7772
rect 240410 7760 240416 7772
rect 240468 7760 240474 7812
rect 245562 7760 245568 7812
rect 245620 7800 245626 7812
rect 330202 7800 330208 7812
rect 245620 7772 330208 7800
rect 245620 7760 245626 7772
rect 330202 7760 330208 7772
rect 330260 7760 330266 7812
rect 456610 7760 456616 7812
rect 456668 7800 456674 7812
rect 548886 7800 548892 7812
rect 456668 7772 548892 7800
rect 456668 7760 456674 7772
rect 548886 7760 548892 7772
rect 548944 7760 548950 7812
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 238846 7732 238852 7744
rect 21968 7704 238852 7732
rect 21968 7692 21974 7704
rect 238846 7692 238852 7704
rect 238904 7692 238910 7744
rect 241974 7692 241980 7744
rect 242032 7732 242038 7744
rect 328546 7732 328552 7744
rect 242032 7704 328552 7732
rect 242032 7692 242038 7704
rect 328546 7692 328552 7704
rect 328604 7692 328610 7744
rect 457990 7692 457996 7744
rect 458048 7732 458054 7744
rect 552382 7732 552388 7744
rect 458048 7704 552388 7732
rect 458048 7692 458054 7704
rect 552382 7692 552388 7704
rect 552440 7692 552446 7744
rect 8846 7624 8852 7676
rect 8904 7664 8910 7676
rect 227533 7667 227591 7673
rect 227533 7664 227545 7667
rect 8904 7636 227545 7664
rect 8904 7624 8910 7636
rect 227533 7633 227545 7636
rect 227579 7633 227591 7667
rect 230658 7664 230664 7676
rect 227533 7627 227591 7633
rect 227640 7636 230664 7664
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 227640 7596 227668 7636
rect 230658 7624 230664 7636
rect 230716 7624 230722 7676
rect 234798 7624 234804 7676
rect 234856 7664 234862 7676
rect 325786 7664 325792 7676
rect 234856 7636 325792 7664
rect 234856 7624 234862 7636
rect 325786 7624 325792 7636
rect 325844 7624 325850 7676
rect 459370 7624 459376 7676
rect 459428 7664 459434 7676
rect 555970 7664 555976 7676
rect 459428 7636 555976 7664
rect 459428 7624 459434 7636
rect 555970 7624 555976 7636
rect 556028 7624 556034 7676
rect 4120 7568 227668 7596
rect 4120 7556 4126 7568
rect 227714 7556 227720 7608
rect 227772 7596 227778 7608
rect 229002 7596 229008 7608
rect 227772 7568 229008 7596
rect 227772 7556 227778 7568
rect 229002 7556 229008 7568
rect 229060 7556 229066 7608
rect 231302 7556 231308 7608
rect 231360 7596 231366 7608
rect 324406 7596 324412 7608
rect 231360 7568 324412 7596
rect 231360 7556 231366 7568
rect 324406 7556 324412 7568
rect 324464 7556 324470 7608
rect 460750 7556 460756 7608
rect 460808 7596 460814 7608
rect 559558 7596 559564 7608
rect 460808 7568 559564 7596
rect 460808 7556 460814 7568
rect 559558 7556 559564 7568
rect 559616 7556 559622 7608
rect 134886 7488 134892 7540
rect 134944 7528 134950 7540
rect 284570 7528 284576 7540
rect 134944 7500 284576 7528
rect 134944 7488 134950 7500
rect 284570 7488 284576 7500
rect 284628 7488 284634 7540
rect 444190 7488 444196 7540
rect 444248 7528 444254 7540
rect 520274 7528 520280 7540
rect 444248 7500 520280 7528
rect 444248 7488 444254 7500
rect 520274 7488 520280 7500
rect 520332 7488 520338 7540
rect 138474 7420 138480 7472
rect 138532 7460 138538 7472
rect 285950 7460 285956 7472
rect 138532 7432 285956 7460
rect 138532 7420 138538 7432
rect 285950 7420 285956 7432
rect 286008 7420 286014 7472
rect 442810 7420 442816 7472
rect 442868 7460 442874 7472
rect 516778 7460 516784 7472
rect 442868 7432 516784 7460
rect 442868 7420 442874 7432
rect 516778 7420 516784 7432
rect 516836 7420 516842 7472
rect 141970 7352 141976 7404
rect 142028 7392 142034 7404
rect 287054 7392 287060 7404
rect 142028 7364 287060 7392
rect 142028 7352 142034 7364
rect 287054 7352 287060 7364
rect 287112 7352 287118 7404
rect 441430 7352 441436 7404
rect 441488 7392 441494 7404
rect 513190 7392 513196 7404
rect 441488 7364 513196 7392
rect 441488 7352 441494 7364
rect 513190 7352 513196 7364
rect 513248 7352 513254 7404
rect 145650 7284 145656 7336
rect 145708 7324 145714 7336
rect 288434 7324 288440 7336
rect 145708 7296 288440 7324
rect 145708 7284 145714 7296
rect 288434 7284 288440 7296
rect 288492 7284 288498 7336
rect 440050 7284 440056 7336
rect 440108 7324 440114 7336
rect 509602 7324 509608 7336
rect 440108 7296 509608 7324
rect 440108 7284 440114 7296
rect 509602 7284 509608 7296
rect 509660 7284 509666 7336
rect 149238 7216 149244 7268
rect 149296 7256 149302 7268
rect 291194 7256 291200 7268
rect 149296 7228 291200 7256
rect 149296 7216 149302 7228
rect 291194 7216 291200 7228
rect 291252 7216 291258 7268
rect 152734 7148 152740 7200
rect 152792 7188 152798 7200
rect 292574 7188 292580 7200
rect 152792 7160 292580 7188
rect 152792 7148 152798 7160
rect 292574 7148 292580 7160
rect 292632 7148 292638 7200
rect 156322 7080 156328 7132
rect 156380 7120 156386 7132
rect 293954 7120 293960 7132
rect 156380 7092 293960 7120
rect 156380 7080 156386 7092
rect 293954 7080 293960 7092
rect 294012 7080 294018 7132
rect 159910 7012 159916 7064
rect 159968 7052 159974 7064
rect 295334 7052 295340 7064
rect 159968 7024 295340 7052
rect 159968 7012 159974 7024
rect 295334 7012 295340 7024
rect 295392 7012 295398 7064
rect 227533 6987 227591 6993
rect 227533 6953 227545 6987
rect 227579 6984 227591 6987
rect 233418 6984 233424 6996
rect 227579 6956 233424 6984
rect 227579 6953 227591 6956
rect 227533 6947 227591 6953
rect 233418 6944 233424 6956
rect 233476 6944 233482 6996
rect 238386 6944 238392 6996
rect 238444 6984 238450 6996
rect 327258 6984 327264 6996
rect 238444 6956 327264 6984
rect 238444 6944 238450 6956
rect 327258 6944 327264 6956
rect 327316 6944 327322 6996
rect 306650 6876 306656 6928
rect 306708 6916 306714 6928
rect 306834 6916 306840 6928
rect 306708 6888 306840 6916
rect 306708 6876 306714 6888
rect 306834 6876 306840 6888
rect 306892 6876 306898 6928
rect 389358 6876 389364 6928
rect 389416 6916 389422 6928
rect 389542 6916 389548 6928
rect 389416 6888 389548 6916
rect 389416 6876 389422 6888
rect 389542 6876 389548 6888
rect 389600 6876 389606 6928
rect 393682 6876 393688 6928
rect 393740 6916 393746 6928
rect 394142 6916 394148 6928
rect 393740 6888 394148 6916
rect 393740 6876 393746 6888
rect 394142 6876 394148 6888
rect 394200 6876 394206 6928
rect 516686 6876 516692 6928
rect 516744 6916 516750 6928
rect 516870 6916 516876 6928
rect 516744 6888 516876 6916
rect 516744 6876 516750 6888
rect 516870 6876 516876 6888
rect 516928 6876 516934 6928
rect 170582 6808 170588 6860
rect 170640 6848 170646 6860
rect 299474 6848 299480 6860
rect 170640 6820 299480 6848
rect 170640 6808 170646 6820
rect 299474 6808 299480 6820
rect 299532 6808 299538 6860
rect 431862 6808 431868 6860
rect 431920 6848 431926 6860
rect 490558 6848 490564 6860
rect 431920 6820 490564 6848
rect 431920 6808 431926 6820
rect 490558 6808 490564 6820
rect 490616 6808 490622 6860
rect 167086 6740 167092 6792
rect 167144 6780 167150 6792
rect 298370 6780 298376 6792
rect 167144 6752 298376 6780
rect 167144 6740 167150 6752
rect 298370 6740 298376 6752
rect 298428 6740 298434 6792
rect 433150 6740 433156 6792
rect 433208 6780 433214 6792
rect 491754 6780 491760 6792
rect 433208 6752 491760 6780
rect 433208 6740 433214 6752
rect 491754 6740 491760 6752
rect 491812 6740 491818 6792
rect 163498 6672 163504 6724
rect 163556 6712 163562 6724
rect 296714 6712 296720 6724
rect 163556 6684 296720 6712
rect 163556 6672 163562 6684
rect 296714 6672 296720 6684
rect 296772 6672 296778 6724
rect 297358 6672 297364 6724
rect 297416 6712 297422 6724
rect 336826 6712 336832 6724
rect 297416 6684 336832 6712
rect 297416 6672 297422 6684
rect 336826 6672 336832 6684
rect 336884 6672 336890 6724
rect 434622 6672 434628 6724
rect 434680 6712 434686 6724
rect 495342 6712 495348 6724
rect 434680 6684 495348 6712
rect 434680 6672 434686 6684
rect 495342 6672 495348 6684
rect 495400 6672 495406 6724
rect 131390 6604 131396 6656
rect 131448 6644 131454 6656
rect 283006 6644 283012 6656
rect 131448 6616 283012 6644
rect 131448 6604 131454 6616
rect 283006 6604 283012 6616
rect 283064 6604 283070 6656
rect 295886 6604 295892 6656
rect 295944 6644 295950 6656
rect 335446 6644 335452 6656
rect 295944 6616 335452 6644
rect 295944 6604 295950 6616
rect 335446 6604 335452 6616
rect 335504 6604 335510 6656
rect 433242 6604 433248 6656
rect 433300 6644 433306 6656
rect 494146 6644 494152 6656
rect 433300 6616 494152 6644
rect 433300 6604 433306 6616
rect 494146 6604 494152 6616
rect 494204 6604 494210 6656
rect 76650 6536 76656 6588
rect 76708 6576 76714 6588
rect 261018 6576 261024 6588
rect 76708 6548 261024 6576
rect 76708 6536 76714 6548
rect 261018 6536 261024 6548
rect 261076 6536 261082 6588
rect 298094 6536 298100 6588
rect 298152 6576 298158 6588
rect 338390 6576 338396 6588
rect 298152 6548 338396 6576
rect 298152 6536 298158 6548
rect 338390 6536 338396 6548
rect 338448 6536 338454 6588
rect 435910 6536 435916 6588
rect 435968 6576 435974 6588
rect 497734 6576 497740 6588
rect 435968 6548 497740 6576
rect 435968 6536 435974 6548
rect 497734 6536 497740 6548
rect 497792 6536 497798 6588
rect 73062 6468 73068 6520
rect 73120 6508 73126 6520
rect 259454 6508 259460 6520
rect 73120 6480 259460 6508
rect 73120 6468 73126 6480
rect 259454 6468 259460 6480
rect 259512 6468 259518 6520
rect 289814 6468 289820 6520
rect 289872 6508 289878 6520
rect 339678 6508 339684 6520
rect 289872 6480 339684 6508
rect 289872 6468 289878 6480
rect 339678 6468 339684 6480
rect 339736 6468 339742 6520
rect 436002 6468 436008 6520
rect 436060 6508 436066 6520
rect 498930 6508 498936 6520
rect 436060 6480 498936 6508
rect 436060 6468 436066 6480
rect 498930 6468 498936 6480
rect 498988 6468 498994 6520
rect 69474 6400 69480 6452
rect 69532 6440 69538 6452
rect 258258 6440 258264 6452
rect 69532 6412 258264 6440
rect 69532 6400 69538 6412
rect 258258 6400 258264 6412
rect 258316 6400 258322 6452
rect 288434 6400 288440 6452
rect 288492 6440 288498 6452
rect 341242 6440 341248 6452
rect 288492 6412 341248 6440
rect 288492 6400 288498 6412
rect 341242 6400 341248 6412
rect 341300 6400 341306 6452
rect 437382 6400 437388 6452
rect 437440 6440 437446 6452
rect 501230 6440 501236 6452
rect 437440 6412 501236 6440
rect 437440 6400 437446 6412
rect 501230 6400 501236 6412
rect 501288 6400 501294 6452
rect 65978 6332 65984 6384
rect 66036 6372 66042 6384
rect 256786 6372 256792 6384
rect 66036 6344 256792 6372
rect 66036 6332 66042 6344
rect 256786 6332 256792 6344
rect 256844 6332 256850 6384
rect 288526 6332 288532 6384
rect 288584 6372 288590 6384
rect 343634 6372 343640 6384
rect 288584 6344 343640 6372
rect 288584 6332 288590 6344
rect 343634 6332 343640 6344
rect 343692 6332 343698 6384
rect 437290 6332 437296 6384
rect 437348 6372 437354 6384
rect 502426 6372 502432 6384
rect 437348 6344 502432 6372
rect 437348 6332 437354 6344
rect 502426 6332 502432 6344
rect 502484 6332 502490 6384
rect 62390 6264 62396 6316
rect 62448 6304 62454 6316
rect 255498 6304 255504 6316
rect 62448 6276 255504 6304
rect 62448 6264 62454 6276
rect 255498 6264 255504 6276
rect 255556 6264 255562 6316
rect 294322 6264 294328 6316
rect 294380 6304 294386 6316
rect 350626 6304 350632 6316
rect 294380 6276 350632 6304
rect 294380 6264 294386 6276
rect 350626 6264 350632 6276
rect 350684 6264 350690 6316
rect 438670 6264 438676 6316
rect 438728 6304 438734 6316
rect 504818 6304 504824 6316
rect 438728 6276 504824 6304
rect 438728 6264 438734 6276
rect 504818 6264 504824 6276
rect 504876 6264 504882 6316
rect 58802 6196 58808 6248
rect 58860 6236 58866 6248
rect 253934 6236 253940 6248
rect 58860 6208 253940 6236
rect 58860 6196 58866 6208
rect 253934 6196 253940 6208
rect 253992 6196 253998 6248
rect 280062 6196 280068 6248
rect 280120 6236 280126 6248
rect 345198 6236 345204 6248
rect 280120 6208 345204 6236
rect 280120 6196 280126 6208
rect 345198 6196 345204 6208
rect 345256 6196 345262 6248
rect 438762 6196 438768 6248
rect 438820 6236 438826 6248
rect 506014 6236 506020 6248
rect 438820 6208 506020 6236
rect 438820 6196 438826 6208
rect 506014 6196 506020 6208
rect 506072 6196 506078 6248
rect 55214 6128 55220 6180
rect 55272 6168 55278 6180
rect 251450 6168 251456 6180
rect 55272 6140 251456 6168
rect 55272 6128 55278 6140
rect 251450 6128 251456 6140
rect 251508 6128 251514 6180
rect 274082 6128 274088 6180
rect 274140 6168 274146 6180
rect 342346 6168 342352 6180
rect 274140 6140 342352 6168
rect 274140 6128 274146 6140
rect 342346 6128 342352 6140
rect 342404 6128 342410 6180
rect 440142 6128 440148 6180
rect 440200 6168 440206 6180
rect 508406 6168 508412 6180
rect 440200 6140 508412 6168
rect 440200 6128 440206 6140
rect 508406 6128 508412 6140
rect 508464 6128 508470 6180
rect 174170 6060 174176 6112
rect 174228 6100 174234 6112
rect 300854 6100 300860 6112
rect 174228 6072 300860 6100
rect 174228 6060 174234 6072
rect 300854 6060 300860 6072
rect 300912 6060 300918 6112
rect 431770 6060 431776 6112
rect 431828 6100 431834 6112
rect 488166 6100 488172 6112
rect 431828 6072 488172 6100
rect 431828 6060 431834 6072
rect 488166 6060 488172 6072
rect 488224 6060 488230 6112
rect 177758 5992 177764 6044
rect 177816 6032 177822 6044
rect 302234 6032 302240 6044
rect 177816 6004 302240 6032
rect 177816 5992 177822 6004
rect 302234 5992 302240 6004
rect 302292 5992 302298 6044
rect 430482 5992 430488 6044
rect 430540 6032 430546 6044
rect 486970 6032 486976 6044
rect 430540 6004 486976 6032
rect 430540 5992 430546 6004
rect 486970 5992 486976 6004
rect 487028 5992 487034 6044
rect 181346 5924 181352 5976
rect 181404 5964 181410 5976
rect 303614 5964 303620 5976
rect 181404 5936 303620 5964
rect 181404 5924 181410 5936
rect 303614 5924 303620 5936
rect 303672 5924 303678 5976
rect 430390 5924 430396 5976
rect 430448 5964 430454 5976
rect 484578 5964 484584 5976
rect 430448 5936 484584 5964
rect 430448 5924 430454 5936
rect 484578 5924 484584 5936
rect 484636 5924 484642 5976
rect 184842 5856 184848 5908
rect 184900 5896 184906 5908
rect 304994 5896 305000 5908
rect 184900 5868 305000 5896
rect 184900 5856 184906 5868
rect 304994 5856 305000 5868
rect 305052 5856 305058 5908
rect 429102 5856 429108 5908
rect 429160 5896 429166 5908
rect 483474 5896 483480 5908
rect 429160 5868 483480 5896
rect 429160 5856 429166 5868
rect 483474 5856 483480 5868
rect 483532 5856 483538 5908
rect 188430 5788 188436 5840
rect 188488 5828 188494 5840
rect 306650 5828 306656 5840
rect 188488 5800 306656 5828
rect 188488 5788 188494 5800
rect 306650 5788 306656 5800
rect 306708 5788 306714 5840
rect 427722 5788 427728 5840
rect 427780 5828 427786 5840
rect 479886 5828 479892 5840
rect 427780 5800 479892 5828
rect 427780 5788 427786 5800
rect 479886 5788 479892 5800
rect 479944 5788 479950 5840
rect 192018 5720 192024 5772
rect 192076 5760 192082 5772
rect 307754 5760 307760 5772
rect 192076 5732 307760 5760
rect 192076 5720 192082 5732
rect 307754 5720 307760 5732
rect 307812 5720 307818 5772
rect 426342 5720 426348 5772
rect 426400 5760 426406 5772
rect 476298 5760 476304 5772
rect 426400 5732 476304 5760
rect 426400 5720 426406 5732
rect 476298 5720 476304 5732
rect 476356 5720 476362 5772
rect 195606 5652 195612 5704
rect 195664 5692 195670 5704
rect 309134 5692 309140 5704
rect 195664 5664 309140 5692
rect 195664 5652 195670 5664
rect 309134 5652 309140 5664
rect 309192 5652 309198 5704
rect 202690 5584 202696 5636
rect 202748 5624 202754 5636
rect 313274 5624 313280 5636
rect 202748 5596 313280 5624
rect 202748 5584 202754 5596
rect 313274 5584 313280 5596
rect 313332 5584 313338 5636
rect 199194 5516 199200 5568
rect 199252 5556 199258 5568
rect 310514 5556 310520 5568
rect 199252 5528 310520 5556
rect 199252 5516 199258 5528
rect 310514 5516 310520 5528
rect 310572 5516 310578 5568
rect 137278 5448 137284 5500
rect 137336 5488 137342 5500
rect 285674 5488 285680 5500
rect 137336 5460 285680 5488
rect 137336 5448 137342 5460
rect 285674 5448 285680 5460
rect 285732 5448 285738 5500
rect 297818 5448 297824 5500
rect 297876 5488 297882 5500
rect 352098 5488 352104 5500
rect 297876 5460 352104 5488
rect 297876 5448 297882 5460
rect 352098 5448 352104 5460
rect 352156 5448 352162 5500
rect 452562 5448 452568 5500
rect 452620 5488 452626 5500
rect 540514 5488 540520 5500
rect 452620 5460 540520 5488
rect 452620 5448 452626 5460
rect 540514 5448 540520 5460
rect 540572 5448 540578 5500
rect 133782 5380 133788 5432
rect 133840 5420 133846 5432
rect 284294 5420 284300 5432
rect 133840 5392 284300 5420
rect 133840 5380 133846 5392
rect 284294 5380 284300 5392
rect 284352 5380 284358 5432
rect 290734 5380 290740 5432
rect 290792 5420 290798 5432
rect 349338 5420 349344 5432
rect 290792 5392 349344 5420
rect 290792 5380 290798 5392
rect 349338 5380 349344 5392
rect 349396 5380 349402 5432
rect 408402 5380 408408 5432
rect 408460 5420 408466 5432
rect 433518 5420 433524 5432
rect 408460 5392 433524 5420
rect 408460 5380 408466 5392
rect 433518 5380 433524 5392
rect 433576 5380 433582 5432
rect 453850 5380 453856 5432
rect 453908 5420 453914 5432
rect 544102 5420 544108 5432
rect 453908 5392 544108 5420
rect 453908 5380 453914 5392
rect 544102 5380 544108 5392
rect 544160 5380 544166 5432
rect 130194 5312 130200 5364
rect 130252 5352 130258 5364
rect 283190 5352 283196 5364
rect 130252 5324 283196 5352
rect 130252 5312 130258 5324
rect 283190 5312 283196 5324
rect 283248 5312 283254 5364
rect 287146 5312 287152 5364
rect 287204 5352 287210 5364
rect 347958 5352 347964 5364
rect 287204 5324 347964 5352
rect 287204 5312 287210 5324
rect 347958 5312 347964 5324
rect 348016 5312 348022 5364
rect 412450 5312 412456 5364
rect 412508 5352 412514 5364
rect 440602 5352 440608 5364
rect 412508 5324 440608 5352
rect 412508 5312 412514 5324
rect 440602 5312 440608 5324
rect 440660 5312 440666 5364
rect 455322 5312 455328 5364
rect 455380 5352 455386 5364
rect 547690 5352 547696 5364
rect 455380 5324 547696 5352
rect 455380 5312 455386 5324
rect 547690 5312 547696 5324
rect 547748 5312 547754 5364
rect 67174 5244 67180 5296
rect 67232 5284 67238 5296
rect 256970 5284 256976 5296
rect 67232 5256 256976 5284
rect 67232 5244 67238 5256
rect 256970 5244 256976 5256
rect 257028 5244 257034 5296
rect 283650 5244 283656 5296
rect 283708 5284 283714 5296
rect 346578 5284 346584 5296
rect 283708 5256 346584 5284
rect 283708 5244 283714 5256
rect 346578 5244 346584 5256
rect 346636 5244 346642 5296
rect 413830 5244 413836 5296
rect 413888 5284 413894 5296
rect 444190 5284 444196 5296
rect 413888 5256 444196 5284
rect 413888 5244 413894 5256
rect 444190 5244 444196 5256
rect 444248 5244 444254 5296
rect 459462 5244 459468 5296
rect 459520 5284 459526 5296
rect 466089 5287 466147 5293
rect 459520 5256 466040 5284
rect 459520 5244 459526 5256
rect 48130 5176 48136 5228
rect 48188 5216 48194 5228
rect 248506 5216 248512 5228
rect 48188 5188 248512 5216
rect 48188 5176 48194 5188
rect 248506 5176 248512 5188
rect 248564 5176 248570 5228
rect 251450 5176 251456 5228
rect 251508 5216 251514 5228
rect 332594 5216 332600 5228
rect 251508 5188 332600 5216
rect 251508 5176 251514 5188
rect 332594 5176 332600 5188
rect 332652 5176 332658 5228
rect 415302 5176 415308 5228
rect 415360 5216 415366 5228
rect 447778 5216 447784 5228
rect 415360 5188 447784 5216
rect 415360 5176 415366 5188
rect 447778 5176 447784 5188
rect 447836 5176 447842 5228
rect 460842 5176 460848 5228
rect 460900 5216 460906 5228
rect 466012 5216 466040 5256
rect 466089 5253 466101 5287
rect 466135 5284 466147 5287
rect 551186 5284 551192 5296
rect 466135 5256 551192 5284
rect 466135 5253 466147 5256
rect 466089 5247 466147 5253
rect 551186 5244 551192 5256
rect 551244 5244 551250 5296
rect 554774 5216 554780 5228
rect 460900 5188 465948 5216
rect 466012 5188 554780 5216
rect 460900 5176 460906 5188
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 236086 5148 236092 5160
rect 17276 5120 236092 5148
rect 17276 5108 17282 5120
rect 236086 5108 236092 5120
rect 236144 5108 236150 5160
rect 247954 5108 247960 5160
rect 248012 5148 248018 5160
rect 331214 5148 331220 5160
rect 248012 5120 331220 5148
rect 248012 5108 248018 5120
rect 331214 5108 331220 5120
rect 331272 5108 331278 5160
rect 416590 5108 416596 5160
rect 416648 5148 416654 5160
rect 451274 5148 451280 5160
rect 416648 5120 451280 5148
rect 416648 5108 416654 5120
rect 451274 5108 451280 5120
rect 451332 5108 451338 5160
rect 461213 5151 461271 5157
rect 461213 5117 461225 5151
rect 461259 5148 461271 5151
rect 461259 5120 462268 5148
rect 461259 5117 461271 5120
rect 461213 5111 461271 5117
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 234706 5080 234712 5092
rect 12492 5052 234712 5080
rect 12492 5040 12498 5052
rect 234706 5040 234712 5052
rect 234764 5040 234770 5092
rect 244366 5040 244372 5092
rect 244424 5080 244430 5092
rect 321557 5083 321615 5089
rect 321557 5080 321569 5083
rect 244424 5052 321569 5080
rect 244424 5040 244430 5052
rect 321557 5049 321569 5052
rect 321603 5049 321615 5083
rect 321557 5043 321615 5049
rect 321646 5040 321652 5092
rect 321704 5080 321710 5092
rect 327074 5080 327080 5092
rect 321704 5052 327080 5080
rect 321704 5040 321710 5052
rect 327074 5040 327080 5052
rect 327132 5040 327138 5092
rect 327169 5083 327227 5089
rect 327169 5049 327181 5083
rect 327215 5080 327227 5083
rect 329834 5080 329840 5092
rect 327215 5052 329840 5080
rect 327215 5049 327227 5052
rect 327169 5043 327227 5049
rect 329834 5040 329840 5052
rect 329892 5040 329898 5092
rect 337102 5040 337108 5092
rect 337160 5080 337166 5092
rect 368566 5080 368572 5092
rect 337160 5052 368572 5080
rect 337160 5040 337166 5052
rect 368566 5040 368572 5052
rect 368624 5040 368630 5092
rect 417970 5040 417976 5092
rect 418028 5080 418034 5092
rect 454862 5080 454868 5092
rect 418028 5052 454868 5080
rect 418028 5040 418034 5052
rect 454862 5040 454868 5052
rect 454920 5040 454926 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 232130 5012 232136 5024
rect 7708 4984 232136 5012
rect 7708 4972 7714 4984
rect 232130 4972 232136 4984
rect 232188 4972 232194 5024
rect 240778 4972 240784 5024
rect 240836 5012 240842 5024
rect 328730 5012 328736 5024
rect 240836 4984 328736 5012
rect 240836 4972 240842 4984
rect 328730 4972 328736 4984
rect 328788 4972 328794 5024
rect 333606 4972 333612 5024
rect 333664 5012 333670 5024
rect 367186 5012 367192 5024
rect 333664 4984 367192 5012
rect 333664 4972 333670 4984
rect 367186 4972 367192 4984
rect 367244 4972 367250 5024
rect 376849 5015 376907 5021
rect 376849 4981 376861 5015
rect 376895 5012 376907 5015
rect 380158 5012 380164 5024
rect 376895 4984 380164 5012
rect 376895 4981 376907 4984
rect 376849 4975 376907 4981
rect 380158 4972 380164 4984
rect 380216 4972 380222 5024
rect 419442 4972 419448 5024
rect 419500 5012 419506 5024
rect 458450 5012 458456 5024
rect 419500 4984 458456 5012
rect 419500 4972 419506 4984
rect 458450 4972 458456 4984
rect 458508 4972 458514 5024
rect 462240 5012 462268 5120
rect 463510 5108 463516 5160
rect 463568 5148 463574 5160
rect 465920 5148 465948 5188
rect 554774 5176 554780 5188
rect 554832 5176 554838 5228
rect 558362 5148 558368 5160
rect 463568 5120 465856 5148
rect 465920 5120 558368 5148
rect 463568 5108 463574 5120
rect 464982 5040 464988 5092
rect 465040 5080 465046 5092
rect 465828 5080 465856 5120
rect 558362 5108 558368 5120
rect 558420 5108 558426 5160
rect 469493 5083 469551 5089
rect 465040 5052 465764 5080
rect 465828 5052 469444 5080
rect 465040 5040 465046 5052
rect 465626 5012 465632 5024
rect 462240 4984 465632 5012
rect 465626 4972 465632 4984
rect 465684 4972 465690 5024
rect 465736 5012 465764 5052
rect 469416 5012 469444 5052
rect 469493 5049 469505 5083
rect 469539 5080 469551 5083
rect 561950 5080 561956 5092
rect 469539 5052 561956 5080
rect 469539 5049 469551 5052
rect 469493 5043 469551 5049
rect 561950 5040 561956 5052
rect 562008 5040 562014 5092
rect 565538 5012 565544 5024
rect 465736 4984 469352 5012
rect 469416 4984 565544 5012
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 224221 4947 224279 4953
rect 224221 4944 224233 4947
rect 2924 4916 224233 4944
rect 2924 4904 2930 4916
rect 224221 4913 224233 4916
rect 224267 4913 224279 4947
rect 229094 4944 229100 4956
rect 224221 4907 224279 4913
rect 224328 4916 229100 4944
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 224328 4876 224356 4916
rect 229094 4904 229100 4916
rect 229152 4904 229158 4956
rect 237190 4904 237196 4956
rect 237248 4944 237254 4956
rect 321646 4944 321652 4956
rect 237248 4916 321652 4944
rect 237248 4904 237254 4916
rect 321646 4904 321652 4916
rect 321704 4904 321710 4956
rect 321741 4947 321799 4953
rect 321741 4913 321753 4947
rect 321787 4944 321799 4947
rect 326985 4947 327043 4953
rect 326985 4944 326997 4947
rect 321787 4916 326997 4944
rect 321787 4913 321799 4916
rect 321741 4907 321799 4913
rect 326985 4913 326997 4916
rect 327031 4913 327043 4947
rect 326985 4907 327043 4913
rect 327074 4904 327080 4956
rect 327132 4944 327138 4956
rect 361666 4944 361672 4956
rect 327132 4916 361672 4944
rect 327132 4904 327138 4916
rect 361666 4904 361672 4916
rect 361724 4904 361730 4956
rect 376757 4947 376815 4953
rect 376757 4913 376769 4947
rect 376803 4944 376815 4947
rect 381538 4944 381544 4956
rect 376803 4916 381544 4944
rect 376803 4913 376815 4916
rect 376757 4907 376815 4913
rect 381538 4904 381544 4916
rect 381596 4904 381602 4956
rect 420730 4904 420736 4956
rect 420788 4944 420794 4956
rect 454681 4947 454739 4953
rect 454681 4944 454693 4947
rect 420788 4916 454693 4944
rect 420788 4904 420794 4916
rect 454681 4913 454693 4916
rect 454727 4913 454739 4947
rect 454681 4907 454739 4913
rect 458082 4904 458088 4956
rect 458140 4944 458146 4956
rect 466089 4947 466147 4953
rect 466089 4944 466101 4947
rect 458140 4916 466101 4944
rect 458140 4904 458146 4916
rect 466089 4913 466101 4916
rect 466135 4913 466147 4947
rect 466089 4907 466147 4913
rect 466178 4904 466184 4956
rect 466236 4944 466242 4956
rect 469324 4944 469352 4984
rect 565538 4972 565544 4984
rect 565596 4972 565602 5024
rect 569034 4944 569040 4956
rect 466236 4916 469260 4944
rect 469324 4916 569040 4944
rect 466236 4904 466242 4916
rect 624 4848 224356 4876
rect 624 4836 630 4848
rect 230106 4836 230112 4888
rect 230164 4876 230170 4888
rect 324314 4876 324320 4888
rect 230164 4848 324320 4876
rect 230164 4836 230170 4848
rect 324314 4836 324320 4848
rect 324372 4836 324378 4888
rect 326338 4836 326344 4888
rect 326396 4876 326402 4888
rect 360378 4876 360384 4888
rect 326396 4848 360384 4876
rect 326396 4836 326402 4848
rect 360378 4836 360384 4848
rect 360436 4836 360442 4888
rect 422202 4836 422208 4888
rect 422260 4876 422266 4888
rect 461213 4879 461271 4885
rect 461213 4876 461225 4879
rect 422260 4848 461225 4876
rect 422260 4836 422266 4848
rect 461213 4845 461225 4848
rect 461259 4845 461271 4879
rect 469122 4876 469128 4888
rect 461213 4839 461271 4845
rect 461596 4848 469128 4876
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 224129 4811 224187 4817
rect 224129 4808 224141 4811
rect 1728 4780 224141 4808
rect 1728 4768 1734 4780
rect 224129 4777 224141 4780
rect 224175 4777 224187 4811
rect 224129 4771 224187 4777
rect 224221 4811 224279 4817
rect 224221 4777 224233 4811
rect 224267 4808 224279 4811
rect 230566 4808 230572 4820
rect 224267 4780 230572 4808
rect 224267 4777 224279 4780
rect 224221 4771 224279 4777
rect 230566 4768 230572 4780
rect 230624 4768 230630 4820
rect 233694 4768 233700 4820
rect 233752 4808 233758 4820
rect 325694 4808 325700 4820
rect 233752 4780 325700 4808
rect 233752 4768 233758 4780
rect 325694 4768 325700 4780
rect 325752 4768 325758 4820
rect 328454 4768 328460 4820
rect 328512 4808 328518 4820
rect 363046 4808 363052 4820
rect 328512 4780 363052 4808
rect 328512 4768 328518 4780
rect 363046 4768 363052 4780
rect 363104 4768 363110 4820
rect 423582 4768 423588 4820
rect 423640 4808 423646 4820
rect 461596 4808 461624 4848
rect 469122 4836 469128 4848
rect 469180 4836 469186 4888
rect 469232 4876 469260 4916
rect 569034 4904 569040 4916
rect 569092 4904 569098 4956
rect 572622 4876 572628 4888
rect 469232 4848 572628 4876
rect 572622 4836 572628 4848
rect 572680 4836 572686 4888
rect 423640 4780 461624 4808
rect 423640 4768 423646 4780
rect 462130 4768 462136 4820
rect 462188 4808 462194 4820
rect 468849 4811 468907 4817
rect 468849 4808 468861 4811
rect 462188 4780 468861 4808
rect 462188 4768 462194 4780
rect 468849 4777 468861 4780
rect 468895 4777 468907 4811
rect 468849 4771 468907 4777
rect 468938 4768 468944 4820
rect 468996 4808 469002 4820
rect 579798 4808 579804 4820
rect 468996 4780 579804 4808
rect 468996 4768 469002 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 212258 4700 212264 4752
rect 212316 4740 212322 4752
rect 316034 4740 316040 4752
rect 212316 4712 316040 4740
rect 212316 4700 212322 4712
rect 316034 4700 316040 4712
rect 316092 4700 316098 4752
rect 318702 4700 318708 4752
rect 318760 4740 318766 4752
rect 318760 4712 323256 4740
rect 318760 4700 318766 4712
rect 215846 4632 215852 4684
rect 215904 4672 215910 4684
rect 317414 4672 317420 4684
rect 215904 4644 317420 4672
rect 215904 4632 215910 4644
rect 317414 4632 317420 4644
rect 317472 4632 317478 4684
rect 323228 4672 323256 4712
rect 323302 4700 323308 4752
rect 323360 4740 323366 4752
rect 358998 4740 359004 4752
rect 323360 4712 359004 4740
rect 323360 4700 323366 4712
rect 358998 4700 359004 4712
rect 359056 4700 359062 4752
rect 451090 4700 451096 4752
rect 451148 4740 451154 4752
rect 536926 4740 536932 4752
rect 451148 4712 536932 4740
rect 451148 4700 451154 4712
rect 536926 4700 536932 4712
rect 536984 4700 536990 4752
rect 333974 4672 333980 4684
rect 323228 4644 333980 4672
rect 333974 4632 333980 4644
rect 334032 4632 334038 4684
rect 365714 4632 365720 4684
rect 365772 4672 365778 4684
rect 366910 4672 366916 4684
rect 365772 4644 366916 4672
rect 365772 4632 365778 4644
rect 366910 4632 366916 4644
rect 366968 4632 366974 4684
rect 449802 4632 449808 4684
rect 449860 4672 449866 4684
rect 533430 4672 533436 4684
rect 449860 4644 533436 4672
rect 449860 4632 449866 4644
rect 533430 4632 533436 4644
rect 533488 4632 533494 4684
rect 219342 4564 219348 4616
rect 219400 4604 219406 4616
rect 318794 4604 318800 4616
rect 219400 4576 318800 4604
rect 219400 4564 219406 4576
rect 318794 4564 318800 4576
rect 318852 4564 318858 4616
rect 321370 4604 321376 4616
rect 318904 4576 321376 4604
rect 222930 4496 222936 4548
rect 222988 4536 222994 4548
rect 318904 4536 318932 4576
rect 321370 4564 321376 4576
rect 321428 4564 321434 4616
rect 322750 4564 322756 4616
rect 322808 4604 322814 4616
rect 337194 4604 337200 4616
rect 322808 4576 337200 4604
rect 322808 4564 322814 4576
rect 337194 4564 337200 4576
rect 337252 4564 337258 4616
rect 448330 4564 448336 4616
rect 448388 4604 448394 4616
rect 529842 4604 529848 4616
rect 448388 4576 529848 4604
rect 448388 4564 448394 4576
rect 529842 4564 529848 4576
rect 529900 4564 529906 4616
rect 222988 4508 318932 4536
rect 222988 4496 222994 4508
rect 320358 4496 320364 4548
rect 320416 4536 320422 4548
rect 335354 4536 335360 4548
rect 320416 4508 335360 4536
rect 320416 4496 320422 4508
rect 335354 4496 335360 4508
rect 335412 4496 335418 4548
rect 350537 4539 350595 4545
rect 350537 4505 350549 4539
rect 350583 4536 350595 4539
rect 353478 4536 353484 4548
rect 350583 4508 353484 4536
rect 350583 4505 350595 4508
rect 350537 4499 350595 4505
rect 353478 4496 353484 4508
rect 353536 4496 353542 4548
rect 447042 4496 447048 4548
rect 447100 4536 447106 4548
rect 526254 4536 526260 4548
rect 447100 4508 526260 4536
rect 447100 4496 447106 4508
rect 526254 4496 526260 4508
rect 526312 4496 526318 4548
rect 226518 4428 226524 4480
rect 226576 4468 226582 4480
rect 322934 4468 322940 4480
rect 226576 4440 322940 4468
rect 226576 4428 226582 4440
rect 322934 4428 322940 4440
rect 322992 4428 322998 4480
rect 325142 4428 325148 4480
rect 325200 4468 325206 4480
rect 338114 4468 338120 4480
rect 325200 4440 338120 4468
rect 325200 4428 325206 4440
rect 338114 4428 338120 4440
rect 338172 4428 338178 4480
rect 350169 4471 350227 4477
rect 350169 4437 350181 4471
rect 350215 4468 350227 4471
rect 352558 4468 352564 4480
rect 350215 4440 352564 4468
rect 350215 4437 350227 4440
rect 350169 4431 350227 4437
rect 352558 4428 352564 4440
rect 352616 4428 352622 4480
rect 445570 4428 445576 4480
rect 445628 4468 445634 4480
rect 522666 4468 522672 4480
rect 445628 4440 522672 4468
rect 445628 4428 445634 4440
rect 522666 4428 522672 4440
rect 522724 4428 522730 4480
rect 201494 4360 201500 4412
rect 201552 4400 201558 4412
rect 271138 4400 271144 4412
rect 201552 4372 271144 4400
rect 201552 4360 201558 4372
rect 271138 4360 271144 4372
rect 271196 4360 271202 4412
rect 301406 4360 301412 4412
rect 301464 4400 301470 4412
rect 350537 4403 350595 4409
rect 350537 4400 350549 4403
rect 301464 4372 350549 4400
rect 301464 4360 301470 4372
rect 350537 4369 350549 4372
rect 350583 4369 350595 4403
rect 350537 4363 350595 4369
rect 444282 4360 444288 4412
rect 444340 4400 444346 4412
rect 519078 4400 519084 4412
rect 444340 4372 519084 4400
rect 444340 4360 444346 4372
rect 519078 4360 519084 4372
rect 519136 4360 519142 4412
rect 205082 4292 205088 4344
rect 205140 4332 205146 4344
rect 272518 4332 272524 4344
rect 205140 4304 272524 4332
rect 205140 4292 205146 4304
rect 272518 4292 272524 4304
rect 272576 4292 272582 4344
rect 304994 4292 305000 4344
rect 305052 4332 305058 4344
rect 354950 4332 354956 4344
rect 305052 4304 354956 4332
rect 305052 4292 305058 4304
rect 354950 4292 354956 4304
rect 355008 4292 355014 4344
rect 442902 4292 442908 4344
rect 442960 4332 442966 4344
rect 515582 4332 515588 4344
rect 442960 4304 515588 4332
rect 442960 4292 442966 4304
rect 515582 4292 515588 4304
rect 515640 4292 515646 4344
rect 224129 4267 224187 4273
rect 224129 4233 224141 4267
rect 224175 4264 224187 4267
rect 230474 4264 230480 4276
rect 224175 4236 230480 4264
rect 224175 4233 224187 4236
rect 224129 4227 224187 4233
rect 230474 4224 230480 4236
rect 230532 4224 230538 4276
rect 269117 4267 269175 4273
rect 269117 4233 269129 4267
rect 269163 4264 269175 4267
rect 278685 4267 278743 4273
rect 278685 4264 278697 4267
rect 269163 4236 278697 4264
rect 269163 4233 269175 4236
rect 269117 4227 269175 4233
rect 278685 4233 278697 4236
rect 278731 4233 278743 4267
rect 278685 4227 278743 4233
rect 308582 4224 308588 4276
rect 308640 4264 308646 4276
rect 356146 4264 356152 4276
rect 308640 4236 356152 4264
rect 308640 4224 308646 4236
rect 356146 4224 356152 4236
rect 356204 4224 356210 4276
rect 441522 4224 441528 4276
rect 441580 4264 441586 4276
rect 511994 4264 512000 4276
rect 441580 4236 512000 4264
rect 441580 4224 441586 4236
rect 511994 4224 512000 4236
rect 512052 4224 512058 4276
rect 124214 4156 124220 4208
rect 124272 4196 124278 4208
rect 125410 4196 125416 4208
rect 124272 4168 125416 4196
rect 124272 4156 124278 4168
rect 125410 4156 125416 4168
rect 125468 4156 125474 4208
rect 140866 4156 140872 4208
rect 140924 4196 140930 4208
rect 142062 4196 142068 4208
rect 140924 4168 142068 4196
rect 140924 4156 140930 4168
rect 142062 4156 142068 4168
rect 142120 4156 142126 4208
rect 150434 4156 150440 4208
rect 150492 4196 150498 4208
rect 151630 4196 151636 4208
rect 150492 4168 151636 4196
rect 150492 4156 150498 4168
rect 151630 4156 151636 4168
rect 151688 4156 151694 4208
rect 158714 4156 158720 4208
rect 158772 4196 158778 4208
rect 160002 4196 160008 4208
rect 158772 4168 160008 4196
rect 158772 4156 158778 4168
rect 160002 4156 160008 4168
rect 160060 4156 160066 4208
rect 175366 4156 175372 4208
rect 175424 4196 175430 4208
rect 176562 4196 176568 4208
rect 175424 4168 176568 4196
rect 175424 4156 175430 4168
rect 176562 4156 176568 4168
rect 176620 4156 176626 4208
rect 209866 4156 209872 4208
rect 209924 4196 209930 4208
rect 211062 4196 211068 4208
rect 209924 4168 211068 4196
rect 209924 4156 209930 4168
rect 211062 4156 211068 4168
rect 211120 4156 211126 4208
rect 287609 4199 287667 4205
rect 284680 4168 285720 4196
rect 57606 4088 57612 4140
rect 57664 4128 57670 4140
rect 250438 4128 250444 4140
rect 57664 4100 250444 4128
rect 57664 4088 57670 4100
rect 250438 4088 250444 4100
rect 250496 4088 250502 4140
rect 268102 4088 268108 4140
rect 268160 4128 268166 4140
rect 269022 4128 269028 4140
rect 268160 4100 269028 4128
rect 268160 4088 268166 4100
rect 269022 4088 269028 4100
rect 269080 4088 269086 4140
rect 273441 4131 273499 4137
rect 273441 4097 273453 4131
rect 273487 4128 273499 4131
rect 284680 4128 284708 4168
rect 273487 4100 284708 4128
rect 273487 4097 273499 4100
rect 273441 4091 273499 4097
rect 284754 4088 284760 4140
rect 284812 4128 284818 4140
rect 285582 4128 285588 4140
rect 284812 4100 285588 4128
rect 284812 4088 284818 4100
rect 285582 4088 285588 4100
rect 285640 4088 285646 4140
rect 285692 4128 285720 4168
rect 287609 4165 287621 4199
rect 287655 4196 287667 4199
rect 287655 4168 287928 4196
rect 287655 4165 287667 4168
rect 287609 4159 287667 4165
rect 287900 4128 287928 4168
rect 312170 4156 312176 4208
rect 312228 4196 312234 4208
rect 357526 4196 357532 4208
rect 312228 4168 357532 4196
rect 312228 4156 312234 4168
rect 357526 4156 357532 4168
rect 357584 4156 357590 4208
rect 424962 4156 424968 4208
rect 425020 4196 425026 4208
rect 472710 4196 472716 4208
rect 425020 4168 472716 4196
rect 425020 4156 425026 4168
rect 472710 4156 472716 4168
rect 472768 4156 472774 4208
rect 295886 4128 295892 4140
rect 285692 4100 287836 4128
rect 287900 4100 295892 4128
rect 50522 4020 50528 4072
rect 50580 4060 50586 4072
rect 249058 4060 249064 4072
rect 50580 4032 249064 4060
rect 50580 4020 50586 4032
rect 249058 4020 249064 4032
rect 249116 4020 249122 4072
rect 264609 4063 264667 4069
rect 264609 4029 264621 4063
rect 264655 4060 264667 4063
rect 269117 4063 269175 4069
rect 269117 4060 269129 4063
rect 264655 4032 269129 4060
rect 264655 4029 264667 4032
rect 264609 4023 264667 4029
rect 269117 4029 269129 4032
rect 269163 4029 269175 4063
rect 269117 4023 269175 4029
rect 278685 4063 278743 4069
rect 278685 4029 278697 4063
rect 278731 4060 278743 4063
rect 282917 4063 282975 4069
rect 282917 4060 282929 4063
rect 278731 4032 282929 4060
rect 278731 4029 278743 4032
rect 278685 4023 278743 4029
rect 282917 4029 282929 4032
rect 282963 4029 282975 4063
rect 287808 4060 287836 4100
rect 295886 4088 295892 4100
rect 295944 4088 295950 4140
rect 296714 4088 296720 4140
rect 296772 4128 296778 4140
rect 297910 4128 297916 4140
rect 296772 4100 297916 4128
rect 296772 4088 296778 4100
rect 297910 4088 297916 4100
rect 297968 4088 297974 4140
rect 300302 4088 300308 4140
rect 300360 4128 300366 4140
rect 332321 4131 332379 4137
rect 332321 4128 332333 4131
rect 300360 4100 332333 4128
rect 300360 4088 300366 4100
rect 332321 4097 332333 4100
rect 332367 4097 332379 4131
rect 332321 4091 332379 4097
rect 332410 4088 332416 4140
rect 332468 4128 332474 4140
rect 333238 4128 333244 4140
rect 332468 4100 333244 4128
rect 332468 4088 332474 4100
rect 333238 4088 333244 4100
rect 333296 4088 333302 4140
rect 334710 4088 334716 4140
rect 334768 4128 334774 4140
rect 335262 4128 335268 4140
rect 334768 4100 335268 4128
rect 334768 4088 334774 4100
rect 335262 4088 335268 4100
rect 335320 4088 335326 4140
rect 335357 4131 335415 4137
rect 335357 4097 335369 4131
rect 335403 4128 335415 4131
rect 338758 4128 338764 4140
rect 335403 4100 338764 4128
rect 335403 4097 335415 4100
rect 335357 4091 335415 4097
rect 338758 4088 338764 4100
rect 338816 4088 338822 4140
rect 339494 4088 339500 4140
rect 339552 4128 339558 4140
rect 340782 4128 340788 4140
rect 339552 4100 340788 4128
rect 339552 4088 339558 4100
rect 340782 4088 340788 4100
rect 340840 4088 340846 4140
rect 340877 4131 340935 4137
rect 340877 4097 340889 4131
rect 340923 4128 340935 4131
rect 345658 4128 345664 4140
rect 340923 4100 345664 4128
rect 340923 4097 340935 4100
rect 340877 4091 340935 4097
rect 345658 4088 345664 4100
rect 345716 4088 345722 4140
rect 347866 4088 347872 4140
rect 347924 4128 347930 4140
rect 349062 4128 349068 4140
rect 347924 4100 349068 4128
rect 347924 4088 347930 4100
rect 349062 4088 349068 4100
rect 349120 4088 349126 4140
rect 349157 4131 349215 4137
rect 349157 4097 349169 4131
rect 349203 4128 349215 4131
rect 351178 4128 351184 4140
rect 349203 4100 351184 4128
rect 349203 4097 349215 4100
rect 349157 4091 349215 4097
rect 351178 4088 351184 4100
rect 351236 4088 351242 4140
rect 351362 4088 351368 4140
rect 351420 4128 351426 4140
rect 351822 4128 351828 4140
rect 351420 4100 351828 4128
rect 351420 4088 351426 4100
rect 351822 4088 351828 4100
rect 351880 4088 351886 4140
rect 352377 4131 352435 4137
rect 352377 4097 352389 4131
rect 352423 4128 352435 4131
rect 358906 4128 358912 4140
rect 352423 4100 358912 4128
rect 352423 4097 352435 4100
rect 352377 4091 352435 4097
rect 358906 4088 358912 4100
rect 358964 4088 358970 4140
rect 362126 4088 362132 4140
rect 362184 4128 362190 4140
rect 362862 4128 362868 4140
rect 362184 4100 362868 4128
rect 362184 4088 362190 4100
rect 362862 4088 362868 4100
rect 362920 4088 362926 4140
rect 363322 4088 363328 4140
rect 363380 4128 363386 4140
rect 364242 4128 364248 4140
rect 363380 4100 364248 4128
rect 363380 4088 363386 4100
rect 364242 4088 364248 4100
rect 364300 4088 364306 4140
rect 369210 4088 369216 4140
rect 369268 4128 369274 4140
rect 369762 4128 369768 4140
rect 369268 4100 369768 4128
rect 369268 4088 369274 4100
rect 369762 4088 369768 4100
rect 369820 4088 369826 4140
rect 370406 4088 370412 4140
rect 370464 4128 370470 4140
rect 371142 4128 371148 4140
rect 370464 4100 371148 4128
rect 370464 4088 370470 4100
rect 371142 4088 371148 4100
rect 371200 4088 371206 4140
rect 377582 4088 377588 4140
rect 377640 4128 377646 4140
rect 378042 4128 378048 4140
rect 377640 4100 378048 4128
rect 377640 4088 377646 4100
rect 378042 4088 378048 4100
rect 378100 4088 378106 4140
rect 378778 4088 378784 4140
rect 378836 4128 378842 4140
rect 385310 4128 385316 4140
rect 378836 4100 385316 4128
rect 378836 4088 378842 4100
rect 385310 4088 385316 4100
rect 385368 4088 385374 4140
rect 390830 4088 390836 4140
rect 390888 4128 390894 4140
rect 391842 4128 391848 4140
rect 390888 4100 391848 4128
rect 390888 4088 390894 4100
rect 391842 4088 391848 4100
rect 391900 4088 391906 4140
rect 393222 4088 393228 4140
rect 393280 4128 393286 4140
rect 395430 4128 395436 4140
rect 393280 4100 395436 4128
rect 393280 4088 393286 4100
rect 395430 4088 395436 4100
rect 395488 4088 395494 4140
rect 398098 4088 398104 4140
rect 398156 4128 398162 4140
rect 403710 4128 403716 4140
rect 398156 4100 403716 4128
rect 398156 4088 398162 4100
rect 403710 4088 403716 4100
rect 403768 4088 403774 4140
rect 409690 4088 409696 4140
rect 409748 4128 409754 4140
rect 437014 4128 437020 4140
rect 409748 4100 437020 4128
rect 409748 4088 409754 4100
rect 437014 4088 437020 4100
rect 437072 4088 437078 4140
rect 445662 4088 445668 4140
rect 445720 4128 445726 4140
rect 521470 4128 521476 4140
rect 445720 4100 521476 4128
rect 445720 4088 445726 4100
rect 521470 4088 521476 4100
rect 521528 4088 521534 4140
rect 529198 4088 529204 4140
rect 529256 4128 529262 4140
rect 575014 4128 575020 4140
rect 529256 4100 575020 4128
rect 529256 4088 529262 4100
rect 575014 4088 575020 4100
rect 575072 4088 575078 4140
rect 298094 4060 298100 4072
rect 287808 4032 298100 4060
rect 282917 4023 282975 4029
rect 298094 4020 298100 4032
rect 298152 4020 298158 4072
rect 302602 4020 302608 4072
rect 302660 4060 302666 4072
rect 309778 4060 309784 4072
rect 302660 4032 309784 4060
rect 302660 4020 302666 4032
rect 309778 4020 309784 4032
rect 309836 4020 309842 4072
rect 314562 4020 314568 4072
rect 314620 4060 314626 4072
rect 350537 4063 350595 4069
rect 350537 4060 350549 4063
rect 314620 4032 350549 4060
rect 314620 4020 314626 4032
rect 350537 4029 350549 4032
rect 350583 4029 350595 4063
rect 373994 4060 374000 4072
rect 350537 4023 350595 4029
rect 352760 4032 374000 4060
rect 46934 3952 46940 4004
rect 46992 3992 46998 4004
rect 248690 3992 248696 4004
rect 46992 3964 248696 3992
rect 46992 3952 46998 3964
rect 248690 3952 248696 3964
rect 248748 3952 248754 4004
rect 257430 3952 257436 4004
rect 257488 3992 257494 4004
rect 287609 3995 287667 4001
rect 287609 3992 287621 3995
rect 257488 3964 287621 3992
rect 257488 3952 257494 3964
rect 287609 3961 287621 3964
rect 287655 3961 287667 3995
rect 287609 3955 287667 3961
rect 287701 3995 287759 4001
rect 287701 3961 287713 3995
rect 287747 3992 287759 3995
rect 297358 3992 297364 4004
rect 287747 3964 297364 3992
rect 287747 3961 287759 3964
rect 287701 3955 287759 3961
rect 297358 3952 297364 3964
rect 297416 3952 297422 4004
rect 313366 3952 313372 4004
rect 313424 3992 313430 4004
rect 352377 3995 352435 4001
rect 352377 3992 352389 3995
rect 313424 3964 352389 3992
rect 313424 3952 313430 3964
rect 352377 3961 352389 3964
rect 352423 3961 352435 3995
rect 352377 3955 352435 3961
rect 352469 3995 352527 4001
rect 352469 3961 352481 3995
rect 352515 3992 352527 3995
rect 352760 3992 352788 4032
rect 373994 4020 374000 4032
rect 374052 4020 374058 4072
rect 383562 4020 383568 4072
rect 383620 4060 383626 4072
rect 384298 4060 384304 4072
rect 383620 4032 384304 4060
rect 383620 4020 383626 4032
rect 384298 4020 384304 4032
rect 384356 4020 384362 4072
rect 393130 4020 393136 4072
rect 393188 4060 393194 4072
rect 396626 4060 396632 4072
rect 393188 4032 396632 4060
rect 393188 4020 393194 4032
rect 396626 4020 396632 4032
rect 396684 4020 396690 4072
rect 411070 4020 411076 4072
rect 411128 4060 411134 4072
rect 439406 4060 439412 4072
rect 411128 4032 439412 4060
rect 411128 4020 411134 4032
rect 439406 4020 439412 4032
rect 439464 4020 439470 4072
rect 442258 4020 442264 4072
rect 442316 4060 442322 4072
rect 442316 4032 446720 4060
rect 442316 4020 442322 4032
rect 352515 3964 352788 3992
rect 352929 3995 352987 4001
rect 352515 3961 352527 3964
rect 352469 3955 352527 3961
rect 352929 3961 352941 3995
rect 352975 3992 352987 3995
rect 355318 3992 355324 4004
rect 352975 3964 355324 3992
rect 352975 3961 352987 3964
rect 352929 3955 352987 3961
rect 355318 3952 355324 3964
rect 355376 3952 355382 4004
rect 355413 3995 355471 4001
rect 355413 3961 355425 3995
rect 355459 3992 355471 3995
rect 359090 3992 359096 4004
rect 355459 3964 359096 3992
rect 355459 3961 355471 3964
rect 355413 3955 355471 3961
rect 359090 3952 359096 3964
rect 359148 3952 359154 4004
rect 359734 3952 359740 4004
rect 359792 3992 359798 4004
rect 377122 3992 377128 4004
rect 359792 3964 377128 3992
rect 359792 3952 359798 3964
rect 377122 3952 377128 3964
rect 377180 3952 377186 4004
rect 406378 3952 406384 4004
rect 406436 3992 406442 4004
rect 414474 3992 414480 4004
rect 406436 3964 414480 3992
rect 406436 3952 406442 3964
rect 414474 3952 414480 3964
rect 414532 3952 414538 4004
rect 420178 3952 420184 4004
rect 420236 3992 420242 4004
rect 423950 3992 423956 4004
rect 420236 3964 423956 3992
rect 420236 3952 420242 3964
rect 423950 3952 423956 3964
rect 424008 3952 424014 4004
rect 424410 3952 424416 4004
rect 424468 3992 424474 4004
rect 425241 3995 425299 4001
rect 425241 3992 425253 3995
rect 424468 3964 425253 3992
rect 424468 3952 424474 3964
rect 425241 3961 425253 3964
rect 425287 3961 425299 3995
rect 425241 3955 425299 3961
rect 426989 3995 427047 4001
rect 426989 3961 427001 3995
rect 427035 3992 427047 3995
rect 446582 3992 446588 4004
rect 427035 3964 446588 3992
rect 427035 3961 427047 3964
rect 426989 3955 427047 3961
rect 446582 3952 446588 3964
rect 446640 3952 446646 4004
rect 446692 3992 446720 4032
rect 448422 4020 448428 4072
rect 448480 4060 448486 4072
rect 528646 4060 528652 4072
rect 448480 4032 528652 4060
rect 448480 4020 448486 4032
rect 528646 4020 528652 4032
rect 528704 4020 528710 4072
rect 530578 4020 530584 4072
rect 530636 4060 530642 4072
rect 582190 4060 582196 4072
rect 530636 4032 582196 4060
rect 530636 4020 530642 4032
rect 582190 4020 582196 4032
rect 582248 4020 582254 4072
rect 449069 3995 449127 4001
rect 449069 3992 449081 3995
rect 446692 3964 449081 3992
rect 449069 3961 449081 3964
rect 449115 3961 449127 3995
rect 449069 3955 449127 3961
rect 451182 3952 451188 4004
rect 451240 3992 451246 4004
rect 535730 3992 535736 4004
rect 451240 3964 535736 3992
rect 451240 3952 451246 3964
rect 535730 3952 535736 3964
rect 535788 3952 535794 4004
rect 45738 3884 45744 3936
rect 45796 3924 45802 3936
rect 247678 3924 247684 3936
rect 45796 3896 247684 3924
rect 45796 3884 45802 3896
rect 247678 3884 247684 3896
rect 247736 3884 247742 3936
rect 282454 3884 282460 3936
rect 282512 3924 282518 3936
rect 320821 3927 320879 3933
rect 320821 3924 320833 3927
rect 282512 3896 320833 3924
rect 282512 3884 282518 3896
rect 320821 3893 320833 3896
rect 320867 3893 320879 3927
rect 320821 3887 320879 3893
rect 326341 3927 326399 3933
rect 326341 3893 326353 3927
rect 326387 3924 326399 3927
rect 332229 3927 332287 3933
rect 332229 3924 332241 3927
rect 326387 3896 332241 3924
rect 326387 3893 326399 3896
rect 326341 3887 326399 3893
rect 332229 3893 332241 3896
rect 332275 3893 332287 3927
rect 332229 3887 332287 3893
rect 332321 3927 332379 3933
rect 332321 3893 332333 3927
rect 332367 3924 332379 3927
rect 335909 3927 335967 3933
rect 332367 3896 335860 3924
rect 332367 3893 332379 3896
rect 332321 3887 332379 3893
rect 39758 3816 39764 3868
rect 39816 3856 39822 3868
rect 238110 3856 238116 3868
rect 39816 3828 238116 3856
rect 39816 3816 39822 3828
rect 238110 3816 238116 3828
rect 238168 3816 238174 3868
rect 264606 3816 264612 3868
rect 264664 3856 264670 3868
rect 273441 3859 273499 3865
rect 273441 3856 273453 3859
rect 264664 3828 273453 3856
rect 264664 3816 264670 3828
rect 273441 3825 273453 3828
rect 273487 3825 273499 3859
rect 288621 3859 288679 3865
rect 288621 3856 288633 3859
rect 273441 3819 273499 3825
rect 285876 3828 288633 3856
rect 20714 3748 20720 3800
rect 20772 3788 20778 3800
rect 35158 3788 35164 3800
rect 20772 3760 35164 3788
rect 20772 3748 20778 3760
rect 35158 3748 35164 3760
rect 35216 3748 35222 3800
rect 38562 3748 38568 3800
rect 38620 3788 38626 3800
rect 245654 3788 245660 3800
rect 38620 3760 245660 3788
rect 38620 3748 38626 3760
rect 245654 3748 245660 3760
rect 245712 3748 245718 3800
rect 278866 3748 278872 3800
rect 278924 3788 278930 3800
rect 285876 3788 285904 3828
rect 288621 3825 288633 3828
rect 288667 3825 288679 3859
rect 288621 3819 288679 3825
rect 289538 3816 289544 3868
rect 289596 3856 289602 3868
rect 335832 3856 335860 3896
rect 335909 3893 335921 3927
rect 335955 3924 335967 3927
rect 365806 3924 365812 3936
rect 335955 3896 365812 3924
rect 335955 3893 335967 3896
rect 335909 3887 335967 3893
rect 365806 3884 365812 3896
rect 365864 3884 365870 3936
rect 371602 3884 371608 3936
rect 371660 3924 371666 3936
rect 376757 3927 376815 3933
rect 376757 3924 376769 3927
rect 371660 3896 376769 3924
rect 371660 3884 371666 3896
rect 376757 3893 376769 3896
rect 376803 3893 376815 3927
rect 376757 3887 376815 3893
rect 404998 3884 405004 3936
rect 405056 3924 405062 3936
rect 416866 3924 416872 3936
rect 405056 3896 416872 3924
rect 405056 3884 405062 3896
rect 416866 3884 416872 3896
rect 416924 3884 416930 3936
rect 420270 3884 420276 3936
rect 420328 3924 420334 3936
rect 450170 3924 450176 3936
rect 420328 3896 450176 3924
rect 420328 3884 420334 3896
rect 450170 3884 450176 3896
rect 450228 3884 450234 3936
rect 453942 3884 453948 3936
rect 454000 3924 454006 3936
rect 542906 3924 542912 3936
rect 454000 3896 542912 3924
rect 454000 3884 454006 3896
rect 542906 3884 542912 3896
rect 542964 3884 542970 3936
rect 342898 3856 342904 3868
rect 289596 3828 335768 3856
rect 335832 3828 342904 3856
rect 289596 3816 289602 3828
rect 278924 3760 285904 3788
rect 278924 3748 278930 3760
rect 285950 3748 285956 3800
rect 286008 3788 286014 3800
rect 332137 3791 332195 3797
rect 332137 3788 332149 3791
rect 286008 3760 332149 3788
rect 286008 3748 286014 3760
rect 332137 3757 332149 3760
rect 332183 3757 332195 3791
rect 332137 3751 332195 3757
rect 332229 3791 332287 3797
rect 332229 3757 332241 3791
rect 332275 3788 332287 3791
rect 335538 3788 335544 3800
rect 332275 3760 335544 3788
rect 332275 3757 332287 3760
rect 332229 3751 332287 3757
rect 335538 3748 335544 3760
rect 335596 3748 335602 3800
rect 335740 3788 335768 3828
rect 342898 3816 342904 3828
rect 342956 3816 342962 3868
rect 343082 3816 343088 3868
rect 343140 3856 343146 3868
rect 369118 3856 369124 3868
rect 343140 3828 369124 3856
rect 343140 3816 343146 3828
rect 369118 3816 369124 3828
rect 369176 3816 369182 3868
rect 372798 3816 372804 3868
rect 372856 3856 372862 3868
rect 373902 3856 373908 3868
rect 372856 3828 373908 3856
rect 372856 3816 372862 3828
rect 373902 3816 373908 3828
rect 373960 3816 373966 3868
rect 399478 3816 399484 3868
rect 399536 3856 399542 3868
rect 407298 3856 407304 3868
rect 399536 3828 407304 3856
rect 399536 3816 399542 3828
rect 407298 3816 407304 3828
rect 407356 3816 407362 3868
rect 412542 3816 412548 3868
rect 412600 3856 412606 3868
rect 442994 3856 443000 3868
rect 412600 3828 443000 3856
rect 412600 3816 412606 3828
rect 442994 3816 443000 3828
rect 443052 3816 443058 3868
rect 453666 3856 453672 3868
rect 445496 3828 453672 3856
rect 341518 3788 341524 3800
rect 335740 3760 341524 3788
rect 341518 3748 341524 3760
rect 341576 3748 341582 3800
rect 341886 3748 341892 3800
rect 341944 3788 341950 3800
rect 370130 3788 370136 3800
rect 341944 3760 370136 3788
rect 341944 3748 341950 3760
rect 370130 3748 370136 3760
rect 370188 3748 370194 3800
rect 373994 3748 374000 3800
rect 374052 3788 374058 3800
rect 375282 3788 375288 3800
rect 374052 3760 375288 3788
rect 374052 3748 374058 3760
rect 375282 3748 375288 3760
rect 375340 3748 375346 3800
rect 399570 3748 399576 3800
rect 399628 3788 399634 3800
rect 408494 3788 408500 3800
rect 399628 3760 408500 3788
rect 399628 3748 399634 3760
rect 408494 3748 408500 3760
rect 408552 3748 408558 3800
rect 413278 3748 413284 3800
rect 413336 3788 413342 3800
rect 413462 3788 413468 3800
rect 413336 3760 413468 3788
rect 413336 3748 413342 3760
rect 413462 3748 413468 3760
rect 413520 3748 413526 3800
rect 413922 3748 413928 3800
rect 413980 3788 413986 3800
rect 445386 3788 445392 3800
rect 413980 3760 445392 3788
rect 413980 3748 413986 3760
rect 445386 3748 445392 3760
rect 445444 3748 445450 3800
rect 32674 3680 32680 3732
rect 32732 3720 32738 3732
rect 243078 3720 243084 3732
rect 32732 3692 243084 3720
rect 32732 3680 32738 3692
rect 243078 3680 243084 3692
rect 243136 3680 243142 3732
rect 282917 3723 282975 3729
rect 282917 3689 282929 3723
rect 282963 3720 282975 3723
rect 287701 3723 287759 3729
rect 287701 3720 287713 3723
rect 282963 3692 287713 3720
rect 282963 3689 282975 3692
rect 282917 3683 282975 3689
rect 287701 3689 287713 3692
rect 287747 3689 287759 3723
rect 287701 3683 287759 3689
rect 292485 3723 292543 3729
rect 292485 3689 292497 3723
rect 292531 3720 292543 3723
rect 326341 3723 326399 3729
rect 326341 3720 326353 3723
rect 292531 3692 326353 3720
rect 292531 3689 292543 3692
rect 292485 3683 292543 3689
rect 326341 3689 326353 3692
rect 326387 3689 326399 3723
rect 326341 3683 326399 3689
rect 326430 3680 326436 3732
rect 326488 3720 326494 3732
rect 328454 3720 328460 3732
rect 326488 3692 328460 3720
rect 326488 3680 326494 3692
rect 328454 3680 328460 3692
rect 328512 3680 328518 3732
rect 331214 3680 331220 3732
rect 331272 3720 331278 3732
rect 335909 3723 335967 3729
rect 335909 3720 335921 3723
rect 331272 3692 335921 3720
rect 331272 3680 331278 3692
rect 335909 3689 335921 3692
rect 335955 3689 335967 3723
rect 335909 3683 335967 3689
rect 338298 3680 338304 3732
rect 338356 3720 338362 3732
rect 368658 3720 368664 3732
rect 338356 3692 368664 3720
rect 338356 3680 338362 3692
rect 368658 3680 368664 3692
rect 368716 3680 368722 3732
rect 375190 3680 375196 3732
rect 375248 3720 375254 3732
rect 383838 3720 383844 3732
rect 375248 3692 383844 3720
rect 375248 3680 375254 3692
rect 383838 3680 383844 3692
rect 383896 3680 383902 3732
rect 402790 3680 402796 3732
rect 402848 3720 402854 3732
rect 419166 3720 419172 3732
rect 402848 3692 419172 3720
rect 402848 3680 402854 3692
rect 419166 3680 419172 3692
rect 419224 3680 419230 3732
rect 421558 3680 421564 3732
rect 421616 3720 421622 3732
rect 422297 3723 422355 3729
rect 422297 3720 422309 3723
rect 421616 3692 422309 3720
rect 421616 3680 421622 3692
rect 422297 3689 422309 3692
rect 422343 3689 422355 3723
rect 422297 3683 422355 3689
rect 428093 3723 428151 3729
rect 428093 3689 428105 3723
rect 428139 3720 428151 3723
rect 431865 3723 431923 3729
rect 428139 3692 431264 3720
rect 428139 3689 428151 3692
rect 428093 3683 428151 3689
rect 24302 3612 24308 3664
rect 24360 3652 24366 3664
rect 239030 3652 239036 3664
rect 24360 3624 239036 3652
rect 24360 3612 24366 3624
rect 239030 3612 239036 3624
rect 239088 3612 239094 3664
rect 262214 3612 262220 3664
rect 262272 3652 262278 3664
rect 320637 3655 320695 3661
rect 320637 3652 320649 3655
rect 262272 3624 320649 3652
rect 262272 3612 262278 3624
rect 320637 3621 320649 3624
rect 320683 3621 320695 3655
rect 325142 3652 325148 3664
rect 320637 3615 320695 3621
rect 320744 3624 325148 3652
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 19978 3584 19984 3596
rect 11296 3556 19984 3584
rect 11296 3544 11302 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 25498 3544 25504 3596
rect 25556 3584 25562 3596
rect 240318 3584 240324 3596
rect 25556 3556 240324 3584
rect 25556 3544 25562 3556
rect 240318 3544 240324 3556
rect 240376 3544 240382 3596
rect 265802 3544 265808 3596
rect 265860 3584 265866 3596
rect 320744 3584 320772 3624
rect 325142 3612 325148 3624
rect 325200 3612 325206 3664
rect 325234 3612 325240 3664
rect 325292 3652 325298 3664
rect 350537 3655 350595 3661
rect 350537 3652 350549 3655
rect 325292 3624 350549 3652
rect 325292 3612 325298 3624
rect 350537 3621 350549 3624
rect 350583 3621 350595 3655
rect 350537 3615 350595 3621
rect 350629 3655 350687 3661
rect 350629 3621 350641 3655
rect 350675 3652 350687 3655
rect 355045 3655 355103 3661
rect 355045 3652 355057 3655
rect 350675 3624 355057 3652
rect 350675 3621 350687 3624
rect 350629 3615 350687 3621
rect 355045 3621 355057 3624
rect 355091 3621 355103 3655
rect 355413 3655 355471 3661
rect 355413 3652 355425 3655
rect 355045 3615 355103 3621
rect 355152 3624 355425 3652
rect 265860 3556 320772 3584
rect 320821 3587 320879 3593
rect 265860 3544 265866 3556
rect 320821 3553 320833 3587
rect 320867 3584 320879 3587
rect 322753 3587 322811 3593
rect 322753 3584 322765 3587
rect 320867 3556 322765 3584
rect 320867 3553 320879 3556
rect 320821 3547 320879 3553
rect 322753 3553 322765 3556
rect 322799 3553 322811 3587
rect 322753 3547 322811 3553
rect 322842 3544 322848 3596
rect 322900 3584 322906 3596
rect 327074 3584 327080 3596
rect 322900 3556 327080 3584
rect 322900 3544 322906 3556
rect 327074 3544 327080 3556
rect 327132 3544 327138 3596
rect 332137 3587 332195 3593
rect 332137 3553 332149 3587
rect 332183 3584 332195 3587
rect 335357 3587 335415 3593
rect 335357 3584 335369 3587
rect 332183 3556 335369 3584
rect 332183 3553 332195 3556
rect 332137 3547 332195 3553
rect 335357 3553 335369 3556
rect 335403 3553 335415 3587
rect 335357 3547 335415 3553
rect 335725 3587 335783 3593
rect 335725 3553 335737 3587
rect 335771 3584 335783 3587
rect 355152 3584 355180 3624
rect 355413 3621 355425 3624
rect 355459 3621 355471 3655
rect 355413 3615 355471 3621
rect 355505 3655 355563 3661
rect 355505 3621 355517 3655
rect 355551 3652 355563 3655
rect 358078 3652 358084 3664
rect 355551 3624 358084 3652
rect 355551 3621 355563 3624
rect 355505 3615 355563 3621
rect 358078 3612 358084 3624
rect 358136 3612 358142 3664
rect 360930 3612 360936 3664
rect 360988 3652 360994 3664
rect 377398 3652 377404 3664
rect 360988 3624 377404 3652
rect 360988 3612 360994 3624
rect 377398 3612 377404 3624
rect 377456 3612 377462 3664
rect 400122 3612 400128 3664
rect 400180 3652 400186 3664
rect 412082 3652 412088 3664
rect 400180 3624 412088 3652
rect 400180 3612 400186 3624
rect 412082 3612 412088 3624
rect 412140 3612 412146 3664
rect 417418 3612 417424 3664
rect 417476 3652 417482 3664
rect 426989 3655 427047 3661
rect 426989 3652 427001 3655
rect 417476 3624 427001 3652
rect 417476 3612 417482 3624
rect 426989 3621 427001 3624
rect 427035 3621 427047 3655
rect 426989 3615 427047 3621
rect 427078 3612 427084 3664
rect 427136 3652 427142 3664
rect 431126 3652 431132 3664
rect 427136 3624 431132 3652
rect 427136 3612 427142 3624
rect 431126 3612 431132 3624
rect 431184 3612 431190 3664
rect 431236 3652 431264 3692
rect 431865 3689 431877 3723
rect 431911 3720 431923 3723
rect 445496 3720 445524 3828
rect 453666 3816 453672 3828
rect 453724 3816 453730 3868
rect 466365 3859 466423 3865
rect 466365 3825 466377 3859
rect 466411 3856 466423 3859
rect 550082 3856 550088 3868
rect 466411 3828 550088 3856
rect 466411 3825 466423 3828
rect 466365 3819 466423 3825
rect 550082 3816 550088 3828
rect 550140 3816 550146 3868
rect 460382 3748 460388 3800
rect 460440 3788 460446 3800
rect 463234 3788 463240 3800
rect 460440 3760 463240 3788
rect 460440 3748 460446 3760
rect 463234 3748 463240 3760
rect 463292 3748 463298 3800
rect 557166 3788 557172 3800
rect 463344 3760 557172 3788
rect 452470 3720 452476 3732
rect 431911 3692 445524 3720
rect 446416 3692 452476 3720
rect 431911 3689 431923 3692
rect 431865 3683 431923 3689
rect 446416 3652 446444 3692
rect 452470 3680 452476 3692
rect 452528 3680 452534 3732
rect 456702 3680 456708 3732
rect 456760 3720 456766 3732
rect 460201 3723 460259 3729
rect 460201 3720 460213 3723
rect 456760 3692 460213 3720
rect 456760 3680 456766 3692
rect 460201 3689 460213 3692
rect 460247 3689 460259 3723
rect 460201 3683 460259 3689
rect 460290 3680 460296 3732
rect 460348 3720 460354 3732
rect 460348 3692 461716 3720
rect 460348 3680 460354 3692
rect 431236 3624 446444 3652
rect 449158 3612 449164 3664
rect 449216 3652 449222 3664
rect 461581 3655 461639 3661
rect 461581 3652 461593 3655
rect 449216 3624 461593 3652
rect 449216 3612 449222 3624
rect 461581 3621 461593 3624
rect 461627 3621 461639 3655
rect 461688 3652 461716 3692
rect 463344 3652 463372 3760
rect 557166 3748 557172 3760
rect 557224 3748 557230 3800
rect 564342 3720 564348 3732
rect 461688 3624 463372 3652
rect 463436 3692 564348 3720
rect 461581 3615 461639 3621
rect 361850 3584 361856 3596
rect 335771 3556 355180 3584
rect 355244 3556 361856 3584
rect 335771 3553 335783 3556
rect 335725 3547 335783 3553
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 234890 3516 234896 3528
rect 14884 3488 234896 3516
rect 14884 3476 14890 3488
rect 234890 3476 234896 3488
rect 234948 3476 234954 3528
rect 258626 3476 258632 3528
rect 258684 3516 258690 3528
rect 320358 3516 320364 3528
rect 258684 3488 320364 3516
rect 258684 3476 258690 3488
rect 320358 3476 320364 3488
rect 320416 3476 320422 3528
rect 320450 3476 320456 3528
rect 320508 3516 320514 3528
rect 321186 3516 321192 3528
rect 320508 3488 321192 3516
rect 320508 3476 320514 3488
rect 321186 3476 321192 3488
rect 321244 3476 321250 3528
rect 321646 3476 321652 3528
rect 321704 3516 321710 3528
rect 355244 3516 355272 3556
rect 361850 3544 361856 3556
rect 361908 3544 361914 3596
rect 382366 3544 382372 3596
rect 382424 3584 382430 3596
rect 386598 3584 386604 3596
rect 382424 3556 386604 3584
rect 382424 3544 382430 3556
rect 386598 3544 386604 3556
rect 386656 3544 386662 3596
rect 402882 3544 402888 3596
rect 402940 3584 402946 3596
rect 420362 3584 420368 3596
rect 402940 3556 420368 3584
rect 402940 3544 402946 3556
rect 420362 3544 420368 3556
rect 420420 3544 420426 3596
rect 420822 3544 420828 3596
rect 420880 3584 420886 3596
rect 460842 3584 460848 3596
rect 420880 3556 460848 3584
rect 420880 3544 420886 3556
rect 460842 3544 460848 3556
rect 460900 3544 460906 3596
rect 462222 3544 462228 3596
rect 462280 3584 462286 3596
rect 463436 3584 463464 3692
rect 564342 3680 564348 3692
rect 564400 3680 564406 3732
rect 463602 3612 463608 3664
rect 463660 3652 463666 3664
rect 566734 3652 566740 3664
rect 463660 3624 566740 3652
rect 463660 3612 463666 3624
rect 566734 3612 566740 3624
rect 566792 3612 566798 3664
rect 462280 3556 463464 3584
rect 462280 3544 462286 3556
rect 466362 3544 466368 3596
rect 466420 3584 466426 3596
rect 571426 3584 571432 3596
rect 466420 3556 571432 3584
rect 466420 3544 466426 3556
rect 571426 3544 571432 3556
rect 571484 3544 571490 3596
rect 363138 3516 363144 3528
rect 321704 3488 355272 3516
rect 355336 3488 363144 3516
rect 321704 3476 321710 3488
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 16022 3408 16028 3460
rect 16080 3448 16086 3460
rect 236270 3448 236276 3460
rect 16080 3420 236276 3448
rect 16080 3408 16086 3420
rect 236270 3408 236276 3420
rect 236328 3408 236334 3460
rect 255038 3408 255044 3460
rect 255096 3448 255102 3460
rect 318702 3448 318708 3460
rect 255096 3420 318708 3448
rect 255096 3408 255102 3420
rect 318702 3408 318708 3420
rect 318760 3408 318766 3460
rect 320637 3451 320695 3457
rect 320637 3417 320649 3451
rect 320683 3448 320695 3451
rect 322750 3448 322756 3460
rect 320683 3420 322756 3448
rect 320683 3417 320695 3420
rect 320637 3411 320695 3417
rect 322750 3408 322756 3420
rect 322808 3408 322814 3460
rect 324038 3408 324044 3460
rect 324096 3448 324102 3460
rect 355336 3448 355364 3488
rect 363138 3476 363144 3488
rect 363196 3476 363202 3528
rect 376757 3519 376815 3525
rect 376757 3516 376769 3519
rect 370240 3488 376769 3516
rect 324096 3420 355364 3448
rect 355413 3451 355471 3457
rect 324096 3408 324102 3420
rect 355413 3417 355425 3451
rect 355459 3448 355471 3451
rect 363598 3448 363604 3460
rect 355459 3420 363604 3448
rect 355459 3417 355471 3420
rect 355413 3411 355471 3417
rect 363598 3408 363604 3420
rect 363656 3408 363662 3460
rect 368014 3408 368020 3460
rect 368072 3448 368078 3460
rect 370240 3448 370268 3488
rect 376757 3485 376769 3488
rect 376803 3485 376815 3519
rect 376757 3479 376815 3485
rect 379974 3476 379980 3528
rect 380032 3516 380038 3528
rect 380802 3516 380808 3528
rect 380032 3488 380808 3516
rect 380032 3476 380038 3488
rect 380802 3476 380808 3488
rect 380860 3476 380866 3528
rect 381170 3476 381176 3528
rect 381228 3516 381234 3528
rect 382182 3516 382188 3528
rect 381228 3488 382188 3516
rect 381228 3476 381234 3488
rect 382182 3476 382188 3488
rect 382240 3476 382246 3528
rect 388254 3476 388260 3528
rect 388312 3516 388318 3528
rect 389082 3516 389088 3528
rect 388312 3488 389088 3516
rect 388312 3476 388318 3488
rect 389082 3476 389088 3488
rect 389140 3476 389146 3528
rect 389266 3476 389272 3528
rect 389324 3516 389330 3528
rect 389453 3519 389511 3525
rect 389453 3516 389465 3519
rect 389324 3488 389465 3516
rect 389324 3476 389330 3488
rect 389453 3485 389465 3488
rect 389499 3485 389511 3519
rect 389453 3479 389511 3485
rect 394602 3476 394608 3528
rect 394660 3516 394666 3528
rect 399018 3516 399024 3528
rect 394660 3488 399024 3516
rect 394660 3476 394666 3488
rect 399018 3476 399024 3488
rect 399076 3476 399082 3528
rect 402238 3476 402244 3528
rect 402296 3516 402302 3528
rect 415670 3516 415676 3528
rect 402296 3488 415676 3516
rect 402296 3476 402302 3488
rect 415670 3476 415676 3488
rect 415728 3476 415734 3528
rect 418062 3476 418068 3528
rect 418120 3516 418126 3528
rect 457254 3516 457260 3528
rect 418120 3488 457260 3516
rect 418120 3476 418126 3488
rect 457254 3476 457260 3488
rect 457312 3476 457318 3528
rect 460201 3519 460259 3525
rect 460201 3485 460213 3519
rect 460247 3516 460259 3519
rect 466181 3519 466239 3525
rect 466181 3516 466193 3519
rect 460247 3488 466193 3516
rect 460247 3485 460259 3488
rect 460201 3479 460259 3485
rect 466181 3485 466193 3488
rect 466227 3485 466239 3519
rect 466181 3479 466239 3485
rect 466270 3476 466276 3528
rect 466328 3516 466334 3528
rect 573818 3516 573824 3528
rect 466328 3488 573824 3516
rect 466328 3476 466334 3488
rect 573818 3476 573824 3488
rect 573876 3476 573882 3528
rect 368072 3420 370268 3448
rect 370317 3451 370375 3457
rect 368072 3408 368078 3420
rect 370317 3417 370329 3451
rect 370363 3448 370375 3451
rect 379698 3448 379704 3460
rect 370363 3420 379704 3448
rect 370363 3417 370375 3420
rect 370317 3411 370375 3417
rect 379698 3408 379704 3420
rect 379756 3408 379762 3460
rect 404262 3408 404268 3460
rect 404320 3448 404326 3460
rect 422754 3448 422760 3460
rect 404320 3420 422760 3448
rect 404320 3408 404326 3420
rect 422754 3408 422760 3420
rect 422812 3408 422818 3460
rect 424318 3408 424324 3460
rect 424376 3448 424382 3460
rect 425146 3448 425152 3460
rect 424376 3420 425152 3448
rect 424376 3408 424382 3420
rect 425146 3408 425152 3420
rect 425204 3408 425210 3460
rect 425241 3451 425299 3457
rect 425241 3417 425253 3451
rect 425287 3448 425299 3451
rect 467926 3448 467932 3460
rect 425287 3420 467932 3448
rect 425287 3417 425299 3420
rect 425241 3411 425299 3417
rect 467926 3408 467932 3420
rect 467984 3408 467990 3460
rect 469030 3408 469036 3460
rect 469088 3448 469094 3460
rect 578602 3448 578608 3460
rect 469088 3420 578608 3448
rect 469088 3408 469094 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 28258 3380 28264 3392
rect 19576 3352 28264 3380
rect 19576 3340 19582 3352
rect 28258 3340 28264 3352
rect 28316 3340 28322 3392
rect 29086 3340 29092 3392
rect 29144 3380 29150 3392
rect 32398 3380 32404 3392
rect 29144 3352 32404 3380
rect 29144 3340 29150 3352
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 34974 3340 34980 3392
rect 35032 3380 35038 3392
rect 57238 3380 57244 3392
rect 35032 3352 57244 3380
rect 35032 3340 35038 3352
rect 57238 3340 57244 3352
rect 57296 3340 57302 3392
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 64690 3340 64696 3392
rect 64748 3380 64754 3392
rect 251818 3380 251824 3392
rect 64748 3352 251824 3380
rect 64748 3340 64754 3352
rect 251818 3340 251824 3352
rect 251876 3340 251882 3392
rect 282825 3383 282883 3389
rect 282825 3349 282837 3383
rect 282871 3380 282883 3383
rect 289814 3380 289820 3392
rect 282871 3352 289820 3380
rect 282871 3349 282883 3352
rect 282825 3343 282883 3349
rect 289814 3340 289820 3352
rect 289872 3340 289878 3392
rect 299106 3340 299112 3392
rect 299164 3380 299170 3392
rect 302878 3380 302884 3392
rect 299164 3352 302884 3380
rect 299164 3340 299170 3352
rect 302878 3340 302884 3352
rect 302936 3340 302942 3392
rect 310974 3340 310980 3392
rect 311032 3380 311038 3392
rect 345477 3383 345535 3389
rect 345477 3380 345489 3383
rect 311032 3352 345489 3380
rect 311032 3340 311038 3352
rect 345477 3349 345489 3352
rect 345523 3349 345535 3383
rect 345477 3343 345535 3349
rect 345937 3383 345995 3389
rect 345937 3349 345949 3383
rect 345983 3380 345995 3383
rect 352929 3383 352987 3389
rect 352929 3380 352941 3383
rect 345983 3352 352941 3380
rect 345983 3349 345995 3352
rect 345937 3343 345995 3349
rect 352929 3349 352941 3352
rect 352975 3349 352987 3383
rect 352929 3343 352987 3349
rect 353754 3340 353760 3392
rect 353812 3380 353818 3392
rect 375650 3380 375656 3392
rect 353812 3352 375656 3380
rect 353812 3340 353818 3352
rect 375650 3340 375656 3352
rect 375708 3340 375714 3392
rect 409782 3340 409788 3392
rect 409840 3380 409846 3392
rect 409840 3352 411024 3380
rect 409840 3340 409846 3352
rect 10042 3272 10048 3324
rect 10100 3312 10106 3324
rect 13078 3312 13084 3324
rect 10100 3284 13084 3312
rect 10100 3272 10106 3284
rect 13078 3272 13084 3284
rect 13136 3272 13142 3324
rect 42150 3272 42156 3324
rect 42208 3312 42214 3324
rect 66898 3312 66904 3324
rect 42208 3284 66904 3312
rect 42208 3272 42214 3284
rect 66898 3272 66904 3284
rect 66956 3272 66962 3324
rect 70670 3272 70676 3324
rect 70728 3312 70734 3324
rect 71682 3312 71688 3324
rect 70728 3284 71688 3312
rect 70728 3272 70734 3284
rect 71682 3272 71688 3284
rect 71740 3272 71746 3324
rect 71866 3272 71872 3324
rect 71924 3312 71930 3324
rect 253198 3312 253204 3324
rect 71924 3284 253204 3312
rect 71924 3272 71930 3284
rect 253198 3272 253204 3284
rect 253256 3272 253262 3324
rect 288434 3312 288440 3324
rect 276400 3284 288440 3312
rect 43346 3204 43352 3256
rect 43404 3244 43410 3256
rect 61378 3244 61384 3256
rect 43404 3216 61384 3244
rect 43404 3204 43410 3216
rect 61378 3204 61384 3216
rect 61436 3204 61442 3256
rect 63586 3204 63592 3256
rect 63644 3244 63650 3256
rect 64782 3244 64788 3256
rect 63644 3216 64788 3244
rect 63644 3204 63650 3216
rect 64782 3204 64788 3216
rect 64840 3204 64846 3256
rect 77846 3204 77852 3256
rect 77904 3244 77910 3256
rect 78582 3244 78588 3256
rect 77904 3216 78588 3244
rect 77904 3204 77910 3216
rect 78582 3204 78588 3216
rect 78640 3204 78646 3256
rect 81434 3204 81440 3256
rect 81492 3244 81498 3256
rect 82722 3244 82728 3256
rect 81492 3216 82728 3244
rect 81492 3204 81498 3216
rect 82722 3204 82728 3216
rect 82780 3204 82786 3256
rect 82817 3247 82875 3253
rect 82817 3213 82829 3247
rect 82863 3244 82875 3247
rect 84838 3244 84844 3256
rect 82863 3216 84844 3244
rect 82863 3213 82875 3216
rect 82817 3207 82875 3213
rect 84838 3204 84844 3216
rect 84896 3204 84902 3256
rect 84930 3204 84936 3256
rect 84988 3244 84994 3256
rect 85482 3244 85488 3256
rect 84988 3216 85488 3244
rect 84988 3204 84994 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 88518 3204 88524 3256
rect 88576 3244 88582 3256
rect 89622 3244 89628 3256
rect 88576 3216 89628 3244
rect 88576 3204 88582 3216
rect 89622 3204 89628 3216
rect 89680 3204 89686 3256
rect 254578 3244 254584 3256
rect 89732 3216 254584 3244
rect 52822 3136 52828 3188
rect 52880 3176 52886 3188
rect 53742 3176 53748 3188
rect 52880 3148 53748 3176
rect 52880 3136 52886 3148
rect 53742 3136 53748 3148
rect 53800 3136 53806 3188
rect 54018 3136 54024 3188
rect 54076 3176 54082 3188
rect 71038 3176 71044 3188
rect 54076 3148 71044 3176
rect 54076 3136 54082 3148
rect 71038 3136 71044 3148
rect 71096 3136 71102 3188
rect 79042 3136 79048 3188
rect 79100 3176 79106 3188
rect 89732 3176 89760 3216
rect 254578 3204 254584 3216
rect 254636 3204 254642 3256
rect 269298 3204 269304 3256
rect 269356 3244 269362 3256
rect 273257 3247 273315 3253
rect 273257 3244 273269 3247
rect 269356 3216 273269 3244
rect 269356 3204 269362 3216
rect 273257 3213 273269 3216
rect 273303 3213 273315 3247
rect 273257 3207 273315 3213
rect 255958 3176 255964 3188
rect 79100 3148 89760 3176
rect 94424 3148 255964 3176
rect 79100 3136 79106 3148
rect 61194 3068 61200 3120
rect 61252 3108 61258 3120
rect 77938 3108 77944 3120
rect 61252 3080 77944 3108
rect 61252 3068 61258 3080
rect 77938 3068 77944 3080
rect 77996 3068 78002 3120
rect 82630 3068 82636 3120
rect 82688 3108 82694 3120
rect 82688 3080 85896 3108
rect 82688 3068 82694 3080
rect 36170 3000 36176 3052
rect 36228 3040 36234 3052
rect 39298 3040 39304 3052
rect 36228 3012 39304 3040
rect 36228 3000 36234 3012
rect 39298 3000 39304 3012
rect 39356 3000 39362 3052
rect 68278 3000 68284 3052
rect 68336 3040 68342 3052
rect 68336 3012 74580 3040
rect 68336 3000 68342 3012
rect 74552 2904 74580 3012
rect 75454 3000 75460 3052
rect 75512 3040 75518 3052
rect 82817 3043 82875 3049
rect 82817 3040 82829 3043
rect 75512 3012 82829 3040
rect 75512 3000 75518 3012
rect 82817 3009 82829 3012
rect 82863 3009 82875 3043
rect 82817 3003 82875 3009
rect 79318 2904 79324 2916
rect 74552 2876 79324 2904
rect 79318 2864 79324 2876
rect 79376 2864 79382 2916
rect 85868 2836 85896 3080
rect 89714 3068 89720 3120
rect 89772 3108 89778 3120
rect 94424 3108 94452 3148
rect 255958 3136 255964 3148
rect 256016 3136 256022 3188
rect 272886 3136 272892 3188
rect 272944 3176 272950 3188
rect 276400 3176 276428 3284
rect 288434 3272 288440 3284
rect 288492 3272 288498 3324
rect 288621 3315 288679 3321
rect 288621 3281 288633 3315
rect 288667 3312 288679 3315
rect 292485 3315 292543 3321
rect 292485 3312 292497 3315
rect 288667 3284 292497 3312
rect 288667 3281 288679 3284
rect 288621 3275 288679 3281
rect 292485 3281 292497 3284
rect 292531 3281 292543 3315
rect 292485 3275 292543 3281
rect 303798 3272 303804 3324
rect 303856 3312 303862 3324
rect 344370 3312 344376 3324
rect 303856 3284 344376 3312
rect 303856 3272 303862 3284
rect 344370 3272 344376 3284
rect 344428 3272 344434 3324
rect 345750 3272 345756 3324
rect 345808 3312 345814 3324
rect 348418 3312 348424 3324
rect 345808 3284 348424 3312
rect 345808 3272 345814 3284
rect 348418 3272 348424 3284
rect 348476 3272 348482 3324
rect 349062 3272 349068 3324
rect 349120 3312 349126 3324
rect 364981 3315 365039 3321
rect 364981 3312 364993 3315
rect 349120 3284 364993 3312
rect 349120 3272 349126 3284
rect 364981 3281 364993 3284
rect 365027 3281 365039 3315
rect 364981 3275 365039 3281
rect 365530 3272 365536 3324
rect 365588 3312 365594 3324
rect 369857 3315 369915 3321
rect 369857 3312 369869 3315
rect 365588 3284 369869 3312
rect 365588 3272 365594 3284
rect 369857 3281 369869 3284
rect 369903 3281 369915 3315
rect 369857 3275 369915 3281
rect 394510 3272 394516 3324
rect 394568 3312 394574 3324
rect 400214 3312 400220 3324
rect 394568 3284 400220 3312
rect 394568 3272 394574 3284
rect 400214 3272 400220 3284
rect 400272 3272 400278 3324
rect 403618 3272 403624 3324
rect 403676 3312 403682 3324
rect 410886 3312 410892 3324
rect 403676 3284 410892 3312
rect 403676 3272 403682 3284
rect 410886 3272 410892 3284
rect 410944 3272 410950 3324
rect 410996 3312 411024 3352
rect 411162 3340 411168 3392
rect 411220 3380 411226 3392
rect 438210 3380 438216 3392
rect 411220 3352 438216 3380
rect 411220 3340 411226 3352
rect 438210 3340 438216 3352
rect 438268 3340 438274 3392
rect 443638 3340 443644 3392
rect 443696 3380 443702 3392
rect 443696 3352 510108 3380
rect 443696 3340 443702 3352
rect 410996 3284 427124 3312
rect 276474 3204 276480 3256
rect 276532 3244 276538 3256
rect 288526 3244 288532 3256
rect 276532 3216 288532 3244
rect 276532 3204 276538 3216
rect 288526 3204 288532 3216
rect 288584 3204 288590 3256
rect 291930 3204 291936 3256
rect 291988 3244 291994 3256
rect 316678 3244 316684 3256
rect 291988 3216 316684 3244
rect 291988 3204 291994 3216
rect 316678 3204 316684 3216
rect 316736 3204 316742 3256
rect 318058 3204 318064 3256
rect 318116 3244 318122 3256
rect 345569 3247 345627 3253
rect 345569 3244 345581 3247
rect 318116 3216 345581 3244
rect 318116 3204 318122 3216
rect 345569 3213 345581 3216
rect 345615 3213 345627 3247
rect 345569 3207 345627 3213
rect 345661 3247 345719 3253
rect 345661 3213 345673 3247
rect 345707 3244 345719 3247
rect 350169 3247 350227 3253
rect 350169 3244 350181 3247
rect 345707 3216 350181 3244
rect 345707 3213 345719 3216
rect 345661 3207 345719 3213
rect 350169 3213 350181 3216
rect 350215 3213 350227 3247
rect 350169 3207 350227 3213
rect 350258 3204 350264 3256
rect 350316 3244 350322 3256
rect 352469 3247 352527 3253
rect 352469 3244 352481 3247
rect 350316 3216 352481 3244
rect 350316 3204 350322 3216
rect 352469 3213 352481 3216
rect 352515 3213 352527 3247
rect 352469 3207 352527 3213
rect 352558 3204 352564 3256
rect 352616 3244 352622 3256
rect 356057 3247 356115 3253
rect 356057 3244 356069 3247
rect 352616 3216 356069 3244
rect 352616 3204 352622 3216
rect 356057 3213 356069 3216
rect 356103 3213 356115 3247
rect 356057 3207 356115 3213
rect 357342 3204 357348 3256
rect 357400 3244 357406 3256
rect 376018 3244 376024 3256
rect 357400 3216 376024 3244
rect 357400 3204 357406 3216
rect 376018 3204 376024 3216
rect 376076 3204 376082 3256
rect 407022 3204 407028 3256
rect 407080 3244 407086 3256
rect 426989 3247 427047 3253
rect 426989 3244 427001 3247
rect 407080 3216 427001 3244
rect 407080 3204 407086 3216
rect 426989 3213 427001 3216
rect 427035 3213 427047 3247
rect 426989 3207 427047 3213
rect 272944 3148 276428 3176
rect 272944 3136 272950 3148
rect 277670 3136 277676 3188
rect 277728 3176 277734 3188
rect 290458 3176 290464 3188
rect 277728 3148 290464 3176
rect 277728 3136 277734 3148
rect 290458 3136 290464 3148
rect 290516 3136 290522 3188
rect 309778 3136 309784 3188
rect 309836 3176 309842 3188
rect 335817 3179 335875 3185
rect 335817 3176 335829 3179
rect 309836 3148 335829 3176
rect 309836 3136 309842 3148
rect 335817 3145 335829 3148
rect 335863 3145 335875 3179
rect 335817 3139 335875 3145
rect 335906 3136 335912 3188
rect 335964 3176 335970 3188
rect 340601 3179 340659 3185
rect 340601 3176 340613 3179
rect 335964 3148 340613 3176
rect 335964 3136 335970 3148
rect 340601 3145 340613 3148
rect 340647 3145 340659 3179
rect 340601 3139 340659 3145
rect 340690 3136 340696 3188
rect 340748 3176 340754 3188
rect 345937 3179 345995 3185
rect 345937 3176 345949 3179
rect 340748 3148 345949 3176
rect 340748 3136 340754 3148
rect 345937 3145 345949 3148
rect 345983 3145 345995 3179
rect 345937 3139 345995 3145
rect 346670 3136 346676 3188
rect 346728 3176 346734 3188
rect 370498 3176 370504 3188
rect 346728 3148 370504 3176
rect 346728 3136 346734 3148
rect 370498 3136 370504 3148
rect 370556 3136 370562 3188
rect 405642 3136 405648 3188
rect 405700 3176 405706 3188
rect 426342 3176 426348 3188
rect 405700 3148 426348 3176
rect 405700 3136 405706 3148
rect 426342 3136 426348 3148
rect 426400 3136 426406 3188
rect 427096 3176 427124 3284
rect 428458 3272 428464 3324
rect 428516 3312 428522 3324
rect 432509 3315 432567 3321
rect 432509 3312 432521 3315
rect 428516 3284 432521 3312
rect 428516 3272 428522 3284
rect 432509 3281 432521 3284
rect 432555 3281 432567 3315
rect 432509 3275 432567 3281
rect 434070 3272 434076 3324
rect 434128 3312 434134 3324
rect 441798 3312 441804 3324
rect 434128 3284 441804 3312
rect 434128 3272 434134 3284
rect 441798 3272 441804 3284
rect 441856 3272 441862 3324
rect 442350 3272 442356 3324
rect 442408 3312 442414 3324
rect 503622 3312 503628 3324
rect 442408 3284 503628 3312
rect 442408 3272 442414 3284
rect 503622 3272 503628 3284
rect 503680 3272 503686 3324
rect 510080 3312 510108 3352
rect 514018 3340 514024 3392
rect 514076 3380 514082 3392
rect 517882 3380 517888 3392
rect 514076 3352 517888 3380
rect 514076 3340 514082 3352
rect 517882 3340 517888 3352
rect 517940 3340 517946 3392
rect 525058 3380 525064 3392
rect 517992 3352 525064 3380
rect 514386 3312 514392 3324
rect 510080 3284 514392 3312
rect 514386 3272 514392 3284
rect 514444 3272 514450 3324
rect 516870 3272 516876 3324
rect 516928 3312 516934 3324
rect 517992 3312 518020 3352
rect 525058 3340 525064 3352
rect 525116 3340 525122 3392
rect 527818 3340 527824 3392
rect 527876 3380 527882 3392
rect 567838 3380 567844 3392
rect 527876 3352 567844 3380
rect 527876 3340 527882 3352
rect 567838 3340 567844 3352
rect 567896 3340 567902 3392
rect 577406 3312 577412 3324
rect 516928 3284 518020 3312
rect 518084 3284 577412 3312
rect 516928 3272 516934 3284
rect 427173 3247 427231 3253
rect 427173 3213 427185 3247
rect 427219 3244 427231 3247
rect 429930 3244 429936 3256
rect 427219 3216 429936 3244
rect 427219 3213 427231 3216
rect 427173 3207 427231 3213
rect 429930 3204 429936 3216
rect 429988 3204 429994 3256
rect 430114 3204 430120 3256
rect 430172 3244 430178 3256
rect 433889 3247 433947 3253
rect 433889 3244 433901 3247
rect 430172 3216 433901 3244
rect 430172 3204 430178 3216
rect 433889 3213 433901 3216
rect 433935 3213 433947 3247
rect 433889 3207 433947 3213
rect 433978 3204 433984 3256
rect 434036 3244 434042 3256
rect 434809 3247 434867 3253
rect 434036 3216 434760 3244
rect 434036 3204 434042 3216
rect 434622 3176 434628 3188
rect 427096 3148 434628 3176
rect 434622 3136 434628 3148
rect 434680 3136 434686 3188
rect 434732 3176 434760 3216
rect 434809 3213 434821 3247
rect 434855 3244 434867 3247
rect 436005 3247 436063 3253
rect 436005 3244 436017 3247
rect 434855 3216 436017 3244
rect 434855 3213 434867 3216
rect 434809 3207 434867 3213
rect 436005 3213 436017 3216
rect 436051 3213 436063 3247
rect 436005 3207 436063 3213
rect 439498 3204 439504 3256
rect 439556 3244 439562 3256
rect 496538 3244 496544 3256
rect 439556 3216 496544 3244
rect 439556 3204 439562 3216
rect 496538 3204 496544 3216
rect 496596 3204 496602 3256
rect 512638 3204 512644 3256
rect 512696 3244 512702 3256
rect 518084 3244 518112 3284
rect 577406 3272 577412 3284
rect 577464 3272 577470 3324
rect 512696 3216 518112 3244
rect 518161 3247 518219 3253
rect 512696 3204 512702 3216
rect 518161 3213 518173 3247
rect 518207 3244 518219 3247
rect 570230 3244 570236 3256
rect 518207 3216 570236 3244
rect 518207 3213 518219 3216
rect 518161 3207 518219 3213
rect 570230 3204 570236 3216
rect 570288 3204 570294 3256
rect 489362 3176 489368 3188
rect 434732 3148 489368 3176
rect 489362 3136 489368 3148
rect 489420 3136 489426 3188
rect 505738 3136 505744 3188
rect 505796 3176 505802 3188
rect 563146 3176 563152 3188
rect 505796 3148 563152 3176
rect 505796 3136 505802 3148
rect 563146 3136 563152 3148
rect 563204 3136 563210 3188
rect 89772 3080 94452 3108
rect 89772 3068 89778 3080
rect 94498 3068 94504 3120
rect 94556 3108 94562 3120
rect 95142 3108 95148 3120
rect 94556 3080 95148 3108
rect 94556 3068 94562 3080
rect 95142 3068 95148 3080
rect 95200 3068 95206 3120
rect 95694 3068 95700 3120
rect 95752 3108 95758 3120
rect 96522 3108 96528 3120
rect 95752 3080 96528 3108
rect 95752 3068 95758 3080
rect 96522 3068 96528 3080
rect 96580 3068 96586 3120
rect 98086 3068 98092 3120
rect 98144 3108 98150 3120
rect 99190 3108 99196 3120
rect 98144 3080 99196 3108
rect 98144 3068 98150 3080
rect 99190 3068 99196 3080
rect 99248 3068 99254 3120
rect 101582 3068 101588 3120
rect 101640 3108 101646 3120
rect 102042 3108 102048 3120
rect 101640 3080 102048 3108
rect 101640 3068 101646 3080
rect 102042 3068 102048 3080
rect 102100 3068 102106 3120
rect 102778 3068 102784 3120
rect 102836 3108 102842 3120
rect 103422 3108 103428 3120
rect 102836 3080 103428 3108
rect 102836 3068 102842 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 105170 3068 105176 3120
rect 105228 3108 105234 3120
rect 106182 3108 106188 3120
rect 105228 3080 106188 3108
rect 105228 3068 105234 3080
rect 106182 3068 106188 3080
rect 106240 3068 106246 3120
rect 106366 3068 106372 3120
rect 106424 3108 106430 3120
rect 107470 3108 107476 3120
rect 106424 3080 107476 3108
rect 106424 3068 106430 3080
rect 107470 3068 107476 3080
rect 107528 3068 107534 3120
rect 257338 3108 257344 3120
rect 108316 3080 257344 3108
rect 86126 3000 86132 3052
rect 86184 3040 86190 3052
rect 95237 3043 95295 3049
rect 86184 3012 95188 3040
rect 86184 3000 86190 3012
rect 93302 2932 93308 2984
rect 93360 2972 93366 2984
rect 94961 2975 95019 2981
rect 94961 2972 94973 2975
rect 93360 2944 94973 2972
rect 93360 2932 93366 2944
rect 94961 2941 94973 2944
rect 95007 2941 95019 2975
rect 95160 2972 95188 3012
rect 95237 3009 95249 3043
rect 95283 3040 95295 3043
rect 97258 3040 97264 3052
rect 95283 3012 97264 3040
rect 95283 3009 95295 3012
rect 95237 3003 95295 3009
rect 97258 3000 97264 3012
rect 97316 3000 97322 3052
rect 95160 2944 96568 2972
rect 94961 2935 95019 2941
rect 95878 2836 95884 2848
rect 85868 2808 95884 2836
rect 95878 2796 95884 2808
rect 95936 2796 95942 2848
rect 96540 2836 96568 2944
rect 96890 2932 96896 2984
rect 96948 2972 96954 2984
rect 108316 2972 108344 3080
rect 257338 3068 257344 3080
rect 257396 3068 257402 3120
rect 295518 3068 295524 3120
rect 295576 3108 295582 3120
rect 319438 3108 319444 3120
rect 295576 3080 319444 3108
rect 295576 3068 295582 3080
rect 319438 3068 319444 3080
rect 319496 3068 319502 3120
rect 322753 3111 322811 3117
rect 322753 3077 322765 3111
rect 322799 3108 322811 3111
rect 327718 3108 327724 3120
rect 322799 3080 327724 3108
rect 322799 3077 322811 3080
rect 322753 3071 322811 3077
rect 327718 3068 327724 3080
rect 327776 3068 327782 3120
rect 328822 3068 328828 3120
rect 328880 3108 328886 3120
rect 355505 3111 355563 3117
rect 355505 3108 355517 3111
rect 328880 3080 355517 3108
rect 328880 3068 328886 3080
rect 355505 3077 355517 3080
rect 355551 3077 355563 3111
rect 355505 3071 355563 3077
rect 355597 3111 355655 3117
rect 355597 3077 355609 3111
rect 355643 3108 355655 3111
rect 359458 3108 359464 3120
rect 355643 3080 359464 3108
rect 355643 3077 355655 3080
rect 355597 3071 355655 3077
rect 359458 3068 359464 3080
rect 359516 3068 359522 3120
rect 364981 3111 365039 3117
rect 364981 3077 364993 3111
rect 365027 3108 365039 3111
rect 372982 3108 372988 3120
rect 365027 3080 372988 3108
rect 365027 3077 365039 3080
rect 364981 3071 365039 3077
rect 372982 3068 372988 3080
rect 373040 3068 373046 3120
rect 398190 3068 398196 3120
rect 398248 3108 398254 3120
rect 398248 3080 401456 3108
rect 398248 3068 398254 3080
rect 258810 3040 258816 3052
rect 96948 2944 108344 2972
rect 108408 3012 258816 3040
rect 96948 2932 96954 2944
rect 103974 2864 103980 2916
rect 104032 2904 104038 2916
rect 108408 2904 108436 3012
rect 258810 3000 258816 3012
rect 258868 3000 258874 3052
rect 273257 3043 273315 3049
rect 273257 3009 273269 3043
rect 273303 3040 273315 3043
rect 282825 3043 282883 3049
rect 282825 3040 282837 3043
rect 273303 3012 282837 3040
rect 273303 3009 273315 3012
rect 273257 3003 273315 3009
rect 282825 3009 282837 3012
rect 282871 3009 282883 3043
rect 282825 3003 282883 3009
rect 293126 3000 293132 3052
rect 293184 3040 293190 3052
rect 312538 3040 312544 3052
rect 293184 3012 312544 3040
rect 293184 3000 293190 3012
rect 312538 3000 312544 3012
rect 312596 3000 312602 3052
rect 315758 3000 315764 3052
rect 315816 3040 315822 3052
rect 323302 3040 323308 3052
rect 315816 3012 323308 3040
rect 315816 3000 315822 3012
rect 323302 3000 323308 3012
rect 323360 3000 323366 3052
rect 327626 3000 327632 3052
rect 327684 3040 327690 3052
rect 335725 3043 335783 3049
rect 335725 3040 335737 3043
rect 327684 3012 335737 3040
rect 327684 3000 327690 3012
rect 335725 3009 335737 3012
rect 335771 3009 335783 3043
rect 335725 3003 335783 3009
rect 335906 3000 335912 3052
rect 335964 3040 335970 3052
rect 360289 3043 360347 3049
rect 360289 3040 360301 3043
rect 335964 3012 360301 3040
rect 335964 3000 335970 3012
rect 360289 3009 360301 3012
rect 360335 3009 360347 3043
rect 360289 3003 360347 3009
rect 360396 3012 364472 3040
rect 112346 2932 112352 2984
rect 112404 2972 112410 2984
rect 113082 2972 113088 2984
rect 112404 2944 113088 2972
rect 112404 2932 112410 2944
rect 113082 2932 113088 2944
rect 113140 2932 113146 2984
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 115934 2932 115940 2984
rect 115992 2972 115998 2984
rect 116946 2972 116952 2984
rect 115992 2944 116952 2972
rect 115992 2932 115998 2944
rect 116946 2932 116952 2944
rect 117004 2932 117010 2984
rect 119430 2932 119436 2984
rect 119488 2972 119494 2984
rect 119982 2972 119988 2984
rect 119488 2944 119988 2972
rect 119488 2932 119494 2944
rect 119982 2932 119988 2944
rect 120040 2932 120046 2984
rect 120626 2932 120632 2984
rect 120684 2972 120690 2984
rect 121362 2972 121368 2984
rect 120684 2944 121368 2972
rect 120684 2932 120690 2944
rect 121362 2932 121368 2944
rect 121420 2932 121426 2984
rect 258718 2972 258724 2984
rect 121472 2944 258724 2972
rect 104032 2876 108436 2904
rect 104032 2864 104038 2876
rect 111150 2864 111156 2916
rect 111208 2904 111214 2916
rect 121472 2904 121500 2944
rect 258718 2932 258724 2944
rect 258776 2932 258782 2984
rect 316954 2932 316960 2984
rect 317012 2972 317018 2984
rect 335633 2975 335691 2981
rect 335633 2972 335645 2975
rect 317012 2944 335645 2972
rect 317012 2932 317018 2944
rect 335633 2941 335645 2944
rect 335679 2941 335691 2975
rect 335633 2935 335691 2941
rect 335817 2975 335875 2981
rect 335817 2941 335829 2975
rect 335863 2972 335875 2975
rect 344370 2972 344376 2984
rect 335863 2944 344376 2972
rect 335863 2941 335875 2944
rect 335817 2935 335875 2941
rect 344370 2932 344376 2944
rect 344428 2932 344434 2984
rect 345474 2932 345480 2984
rect 345532 2972 345538 2984
rect 349157 2975 349215 2981
rect 349157 2972 349169 2975
rect 345532 2944 349169 2972
rect 345532 2932 345538 2944
rect 349157 2941 349169 2944
rect 349203 2941 349215 2975
rect 354861 2975 354919 2981
rect 354861 2972 354873 2975
rect 349157 2935 349215 2941
rect 350644 2944 354873 2972
rect 260098 2904 260104 2916
rect 111208 2876 121500 2904
rect 121564 2876 260104 2904
rect 111208 2864 111214 2876
rect 102594 2836 102600 2848
rect 96540 2808 102600 2836
rect 102594 2796 102600 2808
rect 102652 2796 102658 2848
rect 114738 2796 114744 2848
rect 114796 2836 114802 2848
rect 121564 2836 121592 2876
rect 260098 2864 260104 2876
rect 260156 2864 260162 2916
rect 275278 2864 275284 2916
rect 275336 2904 275342 2916
rect 275922 2904 275928 2916
rect 275336 2876 275928 2904
rect 275336 2864 275342 2876
rect 275922 2864 275928 2876
rect 275980 2864 275986 2916
rect 319254 2864 319260 2916
rect 319312 2904 319318 2916
rect 326338 2904 326344 2916
rect 319312 2876 326344 2904
rect 319312 2864 319318 2876
rect 326338 2864 326344 2876
rect 326396 2864 326402 2916
rect 340693 2907 340751 2913
rect 340693 2873 340705 2907
rect 340739 2904 340751 2907
rect 340874 2904 340880 2916
rect 340739 2876 340880 2904
rect 340739 2873 340751 2876
rect 340693 2867 340751 2873
rect 340874 2864 340880 2876
rect 340932 2864 340938 2916
rect 344278 2864 344284 2916
rect 344336 2904 344342 2916
rect 350644 2904 350672 2944
rect 354861 2941 354873 2944
rect 354907 2941 354919 2975
rect 354861 2935 354919 2941
rect 354950 2932 354956 2984
rect 355008 2972 355014 2984
rect 355962 2972 355968 2984
rect 355008 2944 355968 2972
rect 355008 2932 355014 2944
rect 355962 2932 355968 2944
rect 356020 2932 356026 2984
rect 356057 2975 356115 2981
rect 356057 2941 356069 2975
rect 356103 2972 356115 2975
rect 360396 2972 360424 3012
rect 356103 2944 360424 2972
rect 360473 2975 360531 2981
rect 356103 2941 356115 2944
rect 356057 2935 356115 2941
rect 360473 2941 360485 2975
rect 360519 2972 360531 2975
rect 364444 2972 364472 3012
rect 364518 3000 364524 3052
rect 364576 3040 364582 3052
rect 365530 3040 365536 3052
rect 364576 3012 365536 3040
rect 364576 3000 364582 3012
rect 365530 3000 365536 3012
rect 365588 3000 365594 3052
rect 376386 3000 376392 3052
rect 376444 3040 376450 3052
rect 381630 3040 381636 3052
rect 376444 3012 381636 3040
rect 376444 3000 376450 3012
rect 381630 3000 381636 3012
rect 381688 3000 381694 3052
rect 395890 3000 395896 3052
rect 395948 3040 395954 3052
rect 401318 3040 401324 3052
rect 395948 3012 401324 3040
rect 395948 3000 395954 3012
rect 401318 3000 401324 3012
rect 401376 3000 401382 3052
rect 401428 3040 401456 3080
rect 411898 3068 411904 3120
rect 411956 3108 411962 3120
rect 428734 3108 428740 3120
rect 411956 3080 428740 3108
rect 411956 3068 411962 3080
rect 428734 3068 428740 3080
rect 428792 3068 428798 3120
rect 431218 3068 431224 3120
rect 431276 3108 431282 3120
rect 431276 3080 477632 3108
rect 431276 3068 431282 3080
rect 404906 3040 404912 3052
rect 401428 3012 404912 3040
rect 404906 3000 404912 3012
rect 404964 3000 404970 3052
rect 416682 3000 416688 3052
rect 416740 3040 416746 3052
rect 428093 3043 428151 3049
rect 428093 3040 428105 3043
rect 416740 3012 428105 3040
rect 416740 3000 416746 3012
rect 428093 3009 428105 3012
rect 428139 3009 428151 3043
rect 428093 3003 428151 3009
rect 428185 3043 428243 3049
rect 428185 3009 428197 3043
rect 428231 3040 428243 3043
rect 435818 3040 435824 3052
rect 428231 3012 435824 3040
rect 428231 3009 428243 3012
rect 428185 3003 428243 3009
rect 435818 3000 435824 3012
rect 435876 3000 435882 3052
rect 435913 3043 435971 3049
rect 435913 3009 435925 3043
rect 435959 3040 435971 3043
rect 475102 3040 475108 3052
rect 435959 3012 475108 3040
rect 435959 3009 435971 3012
rect 435913 3003 435971 3009
rect 475102 3000 475108 3012
rect 475160 3000 475166 3052
rect 475378 3000 475384 3052
rect 475436 3040 475442 3052
rect 477494 3040 477500 3052
rect 475436 3012 477500 3040
rect 475436 3000 475442 3012
rect 477494 3000 477500 3012
rect 477552 3000 477558 3052
rect 477604 3040 477632 3080
rect 524966 3068 524972 3120
rect 525024 3108 525030 3120
rect 560754 3108 560760 3120
rect 525024 3080 560760 3108
rect 525024 3068 525030 3080
rect 560754 3068 560760 3080
rect 560812 3068 560818 3120
rect 482278 3040 482284 3052
rect 477604 3012 482284 3040
rect 482278 3000 482284 3012
rect 482336 3000 482342 3052
rect 509878 3000 509884 3052
rect 509936 3040 509942 3052
rect 518161 3043 518219 3049
rect 518161 3040 518173 3043
rect 509936 3012 518173 3040
rect 509936 3000 509942 3012
rect 518161 3009 518173 3012
rect 518207 3009 518219 3043
rect 518161 3003 518219 3009
rect 523678 3000 523684 3052
rect 523736 3040 523742 3052
rect 553578 3040 553584 3052
rect 523736 3012 553584 3040
rect 523736 3000 523742 3012
rect 553578 3000 553584 3012
rect 553636 3000 553642 3052
rect 374086 2972 374092 2984
rect 360519 2944 362356 2972
rect 364444 2944 374092 2972
rect 360519 2941 360531 2944
rect 360473 2935 360531 2941
rect 344336 2876 350672 2904
rect 350813 2907 350871 2913
rect 344336 2864 344342 2876
rect 350813 2873 350825 2907
rect 350859 2904 350871 2907
rect 355597 2907 355655 2913
rect 355597 2904 355609 2907
rect 350859 2876 355609 2904
rect 350859 2873 350871 2876
rect 350813 2867 350871 2873
rect 355597 2873 355609 2876
rect 355643 2873 355655 2907
rect 362218 2904 362224 2916
rect 355597 2867 355655 2873
rect 355796 2876 362224 2904
rect 114796 2808 121592 2836
rect 114796 2796 114802 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 261478 2836 261484 2848
rect 121880 2808 261484 2836
rect 121880 2796 121886 2808
rect 261478 2796 261484 2808
rect 261536 2796 261542 2848
rect 330018 2796 330024 2848
rect 330076 2836 330082 2848
rect 335538 2836 335544 2848
rect 330076 2808 335544 2836
rect 330076 2796 330082 2808
rect 335538 2796 335544 2808
rect 335596 2796 335602 2848
rect 335633 2839 335691 2845
rect 335633 2805 335645 2839
rect 335679 2836 335691 2839
rect 340785 2839 340843 2845
rect 340785 2836 340797 2839
rect 335679 2808 340797 2836
rect 335679 2805 335691 2808
rect 335633 2799 335691 2805
rect 340785 2805 340797 2808
rect 340831 2805 340843 2839
rect 340785 2799 340843 2805
rect 345569 2839 345627 2845
rect 345569 2805 345581 2839
rect 345615 2836 345627 2839
rect 355689 2839 355747 2845
rect 355689 2836 355701 2839
rect 345615 2808 355701 2836
rect 345615 2805 345627 2808
rect 345569 2799 345627 2805
rect 355689 2805 355701 2808
rect 355735 2805 355747 2839
rect 355689 2799 355747 2805
rect 355505 2771 355563 2777
rect 355505 2737 355517 2771
rect 355551 2768 355563 2771
rect 355796 2768 355824 2876
rect 362218 2864 362224 2876
rect 362276 2864 362282 2916
rect 362328 2904 362356 2944
rect 374086 2932 374092 2944
rect 374144 2932 374150 2984
rect 395982 2932 395988 2984
rect 396040 2972 396046 2984
rect 402514 2972 402520 2984
rect 396040 2944 402520 2972
rect 396040 2932 396046 2944
rect 402514 2932 402520 2944
rect 402572 2932 402578 2984
rect 413462 2932 413468 2984
rect 413520 2972 413526 2984
rect 432322 2972 432328 2984
rect 413520 2944 432328 2972
rect 413520 2932 413526 2944
rect 432322 2932 432328 2944
rect 432380 2932 432386 2984
rect 459646 2972 459652 2984
rect 432432 2944 459652 2972
rect 367278 2904 367284 2916
rect 362328 2876 367284 2904
rect 367278 2864 367284 2876
rect 367336 2864 367342 2916
rect 385862 2864 385868 2916
rect 385920 2904 385926 2916
rect 387058 2904 387064 2916
rect 385920 2876 387064 2904
rect 385920 2864 385926 2876
rect 387058 2864 387064 2876
rect 387116 2864 387122 2916
rect 422297 2907 422355 2913
rect 422297 2873 422309 2907
rect 422343 2904 422355 2907
rect 422343 2876 428412 2904
rect 422343 2873 422355 2876
rect 422297 2867 422355 2873
rect 355965 2839 356023 2845
rect 355965 2805 355977 2839
rect 356011 2836 356023 2839
rect 356698 2836 356704 2848
rect 356011 2808 356704 2836
rect 356011 2805 356023 2808
rect 355965 2799 356023 2805
rect 356698 2796 356704 2808
rect 356756 2796 356762 2848
rect 375834 2836 375840 2848
rect 356900 2808 375840 2836
rect 355551 2740 355824 2768
rect 355551 2737 355563 2740
rect 355505 2731 355563 2737
rect 356146 2660 356152 2712
rect 356204 2700 356210 2712
rect 356900 2700 356928 2808
rect 375834 2796 375840 2808
rect 375892 2796 375898 2848
rect 388438 2836 388444 2848
rect 387076 2808 388444 2836
rect 387076 2780 387104 2808
rect 388438 2796 388444 2808
rect 388496 2796 388502 2848
rect 416038 2796 416044 2848
rect 416096 2836 416102 2848
rect 428185 2839 428243 2845
rect 428185 2836 428197 2839
rect 416096 2808 428197 2836
rect 416096 2796 416102 2808
rect 428185 2805 428197 2808
rect 428231 2805 428243 2839
rect 428185 2799 428243 2805
rect 387058 2728 387064 2780
rect 387116 2728 387122 2780
rect 428384 2768 428412 2876
rect 431310 2864 431316 2916
rect 431368 2904 431374 2916
rect 432432 2904 432460 2944
rect 459646 2932 459652 2944
rect 459704 2932 459710 2984
rect 461581 2975 461639 2981
rect 461581 2941 461593 2975
rect 461627 2972 461639 2975
rect 481082 2972 481088 2984
rect 461627 2944 481088 2972
rect 461627 2941 461639 2944
rect 461581 2935 461639 2941
rect 481082 2932 481088 2944
rect 481140 2932 481146 2984
rect 521010 2932 521016 2984
rect 521068 2972 521074 2984
rect 546494 2972 546500 2984
rect 521068 2944 546500 2972
rect 521068 2932 521074 2944
rect 546494 2932 546500 2944
rect 546552 2932 546558 2984
rect 431368 2876 432460 2904
rect 432509 2907 432567 2913
rect 431368 2864 431374 2876
rect 432509 2873 432521 2907
rect 432555 2904 432567 2907
rect 435913 2907 435971 2913
rect 435913 2904 435925 2907
rect 432555 2876 435925 2904
rect 432555 2873 432567 2876
rect 432509 2867 432567 2873
rect 435913 2873 435925 2876
rect 435959 2873 435971 2907
rect 435913 2867 435971 2873
rect 436005 2907 436063 2913
rect 436005 2873 436017 2907
rect 436051 2904 436063 2907
rect 448974 2904 448980 2916
rect 436051 2876 448980 2904
rect 436051 2873 436063 2876
rect 436005 2867 436063 2873
rect 448974 2864 448980 2876
rect 449032 2864 449038 2916
rect 449069 2907 449127 2913
rect 449069 2873 449081 2907
rect 449115 2904 449127 2907
rect 473906 2904 473912 2916
rect 449115 2876 473912 2904
rect 449115 2873 449127 2876
rect 449069 2867 449127 2873
rect 473906 2864 473912 2876
rect 473964 2864 473970 2916
rect 520918 2864 520924 2916
rect 520976 2904 520982 2916
rect 539318 2904 539324 2916
rect 520976 2876 539324 2904
rect 520976 2864 520982 2876
rect 539318 2864 539324 2876
rect 539376 2864 539382 2916
rect 438118 2796 438124 2848
rect 438176 2836 438182 2848
rect 466822 2836 466828 2848
rect 438176 2808 466828 2836
rect 438176 2796 438182 2808
rect 466822 2796 466828 2808
rect 466880 2796 466886 2848
rect 518158 2796 518164 2848
rect 518216 2836 518222 2848
rect 532234 2836 532240 2848
rect 518216 2808 532240 2836
rect 518216 2796 518222 2808
rect 532234 2796 532240 2808
rect 532292 2796 532298 2848
rect 431865 2771 431923 2777
rect 431865 2768 431877 2771
rect 428384 2740 431877 2768
rect 431865 2737 431877 2740
rect 431911 2737 431923 2771
rect 431865 2731 431923 2737
rect 454681 2771 454739 2777
rect 454681 2737 454693 2771
rect 454727 2768 454739 2771
rect 462038 2768 462044 2780
rect 454727 2740 462044 2768
rect 454727 2737 454739 2740
rect 454681 2731 454739 2737
rect 462038 2728 462044 2740
rect 462096 2728 462102 2780
rect 356204 2672 356928 2700
rect 356204 2660 356210 2672
rect 261018 1096 261024 1148
rect 261076 1136 261082 1148
rect 264609 1139 264667 1145
rect 264609 1136 264621 1139
rect 261076 1108 264621 1136
rect 261076 1096 261082 1108
rect 264609 1105 264621 1108
rect 264655 1105 264667 1139
rect 264609 1099 264667 1105
rect 394142 1028 394148 1080
rect 394200 1068 394206 1080
rect 394237 1071 394295 1077
rect 394237 1068 394249 1071
rect 394200 1040 394249 1068
rect 394200 1028 394206 1040
rect 394237 1037 394249 1040
rect 394283 1037 394295 1071
rect 394237 1031 394295 1037
rect 23106 552 23112 604
rect 23164 592 23170 604
rect 23382 592 23388 604
rect 23164 564 23388 592
rect 23164 552 23170 564
rect 23382 552 23388 564
rect 23440 552 23446 604
rect 164694 552 164700 604
rect 164752 592 164758 604
rect 165522 592 165528 604
rect 164752 564 165528 592
rect 164752 552 164758 564
rect 165522 552 165528 564
rect 165580 552 165586 604
rect 165890 552 165896 604
rect 165948 592 165954 604
rect 166902 592 166908 604
rect 165948 564 166908 592
rect 165948 552 165954 564
rect 166902 552 166908 564
rect 166960 552 166966 604
rect 169386 552 169392 604
rect 169444 592 169450 604
rect 169662 592 169668 604
rect 169444 564 169668 592
rect 169444 552 169450 564
rect 169662 552 169668 564
rect 169720 552 169726 604
rect 182542 552 182548 604
rect 182600 592 182606 604
rect 183462 592 183468 604
rect 182600 564 183468 592
rect 182600 552 182606 564
rect 183462 552 183468 564
rect 183520 552 183526 604
rect 183738 552 183744 604
rect 183796 592 183802 604
rect 184750 592 184756 604
rect 183796 564 184756 592
rect 183796 552 183802 564
rect 184750 552 184756 564
rect 184808 552 184814 604
rect 187234 552 187240 604
rect 187292 592 187298 604
rect 187602 592 187608 604
rect 187292 564 187608 592
rect 187292 552 187298 564
rect 187602 552 187608 564
rect 187660 552 187666 604
rect 189626 552 189632 604
rect 189684 592 189690 604
rect 190362 592 190368 604
rect 189684 564 190368 592
rect 189684 552 189690 564
rect 190362 552 190368 564
rect 190420 552 190426 604
rect 281258 552 281264 604
rect 281316 592 281322 604
rect 281442 592 281448 604
rect 281316 564 281448 592
rect 281316 552 281322 564
rect 281442 552 281448 564
rect 281500 552 281506 604
rect 358538 552 358544 604
rect 358596 592 358602 604
rect 358722 592 358728 604
rect 358596 564 358728 592
rect 358596 552 358602 564
rect 358722 552 358728 564
rect 358780 552 358786 604
rect 384666 552 384672 604
rect 384724 592 384730 604
rect 384942 592 384948 604
rect 384724 564 384948 592
rect 384724 552 384730 564
rect 384942 552 384948 564
rect 385000 552 385006 604
rect 389450 592 389456 604
rect 389411 564 389456 592
rect 389450 552 389456 564
rect 389508 552 389514 604
rect 394234 592 394240 604
rect 394195 564 394240 592
rect 394234 552 394240 564
rect 394292 552 394298 604
rect 405918 552 405924 604
rect 405976 592 405982 604
rect 406102 592 406108 604
rect 405976 564 406108 592
rect 405976 552 405982 564
rect 406102 552 406108 564
rect 406160 552 406166 604
rect 463694 552 463700 604
rect 463752 592 463758 604
rect 464430 592 464436 604
rect 463752 564 464436 592
rect 463752 552 463758 564
rect 464430 552 464436 564
rect 464488 552 464494 604
rect 469214 552 469220 604
rect 469272 592 469278 604
rect 470318 592 470324 604
rect 469272 564 470324 592
rect 469272 552 469278 564
rect 470318 552 470324 564
rect 470376 552 470382 604
<< via1 >>
rect 202788 700952 202840 701004
rect 358820 700952 358872 701004
rect 170312 700884 170364 700936
rect 362960 700884 363012 700936
rect 328368 700816 328420 700868
rect 527180 700816 527232 700868
rect 329748 700748 329800 700800
rect 543464 700748 543516 700800
rect 154120 700680 154172 700732
rect 367100 700680 367152 700732
rect 137836 700612 137888 700664
rect 364340 700612 364392 700664
rect 105452 700544 105504 700596
rect 368480 700544 368532 700596
rect 89168 700476 89220 700528
rect 374000 700476 374052 700528
rect 72976 700408 73028 700460
rect 371240 700408 371292 700460
rect 40500 700340 40552 700392
rect 375380 700340 375432 700392
rect 24308 700272 24360 700324
rect 379520 700272 379572 700324
rect 218980 700204 219032 700256
rect 360200 700204 360252 700256
rect 336648 700136 336700 700188
rect 478512 700136 478564 700188
rect 335268 700068 335320 700120
rect 462320 700068 462372 700120
rect 235172 700000 235224 700052
rect 356060 700000 356112 700052
rect 267648 699932 267700 699984
rect 351920 699932 351972 699984
rect 283840 699864 283892 699916
rect 354680 699864 354732 699916
rect 343548 699796 343600 699848
rect 413652 699796 413704 699848
rect 340788 699728 340840 699780
rect 397460 699728 397512 699780
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 332508 699660 332560 699712
rect 346400 699660 346452 699712
rect 347780 699660 347832 699712
rect 348792 699660 348844 699712
rect 321468 696940 321520 696992
rect 580172 696940 580224 696992
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 364616 687760 364668 687812
rect 365168 687760 365220 687812
rect 324228 685856 324280 685908
rect 580172 685856 580224 685908
rect 364616 685788 364668 685840
rect 429292 684428 429344 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 382280 681708 382332 681760
rect 364524 676243 364576 676252
rect 364524 676209 364533 676243
rect 364533 676209 364567 676243
rect 364567 676209 364576 676243
rect 364524 676200 364576 676209
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 320088 673480 320140 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 386420 667904 386472 667956
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 559380 666544 559432 666596
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 383660 652740 383712 652792
rect 315948 650020 316000 650072
rect 580172 650020 580224 650072
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 317328 638936 317380 638988
rect 580172 638936 580224 638988
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 313188 626560 313240 626612
rect 580172 626560 580224 626612
rect 3424 623772 3476 623824
rect 387800 623772 387852 623824
rect 364616 618196 364668 618248
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 3424 609968 3476 610020
rect 391940 609968 391992 610020
rect 364524 608651 364576 608660
rect 364524 608617 364533 608651
rect 364533 608617 364567 608651
rect 364567 608617 364576 608651
rect 364524 608608 364576 608617
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 309048 603100 309100 603152
rect 580172 603100 580224 603152
rect 429568 601672 429620 601724
rect 559288 601672 559340 601724
rect 364616 598927 364668 598936
rect 364616 598893 364625 598927
rect 364625 598893 364659 598927
rect 364659 598893 364668 598927
rect 364616 598884 364668 598893
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 390560 594804 390612 594856
rect 311808 592016 311860 592068
rect 580172 592016 580224 592068
rect 364708 589296 364760 589348
rect 429660 589296 429712 589348
rect 559380 589296 559432 589348
rect 344468 584672 344520 584724
rect 364708 584672 364760 584724
rect 300768 584604 300820 584656
rect 350816 584604 350868 584656
rect 338212 584536 338264 584588
rect 429660 584536 429712 584588
rect 331864 584468 331916 584520
rect 494244 584468 494296 584520
rect 325516 584400 325568 584452
rect 559380 584400 559432 584452
rect 304540 583652 304592 583704
rect 471244 583652 471296 583704
rect 298192 583584 298244 583636
rect 469772 583584 469824 583636
rect 262404 583516 262456 583568
rect 580724 583516 580776 583568
rect 256056 583448 256108 583500
rect 580448 583448 580500 583500
rect 251824 583380 251876 583432
rect 580356 583380 580408 583432
rect 6644 583312 6696 583364
rect 399208 583312 399260 583364
rect 6368 583244 6420 583296
rect 403440 583244 403492 583296
rect 4712 583176 4764 583228
rect 405556 583176 405608 583228
rect 5356 583108 5408 583160
rect 409788 583108 409840 583160
rect 3240 583040 3292 583092
rect 407672 583040 407724 583092
rect 5448 582972 5500 583024
rect 411904 582972 411956 583024
rect 14464 582904 14516 582956
rect 424508 582904 424560 582956
rect 5264 582836 5316 582888
rect 418160 582836 418212 582888
rect 15844 582768 15896 582820
rect 430856 582768 430908 582820
rect 4068 582700 4120 582752
rect 422392 582700 422444 582752
rect 17224 582632 17276 582684
rect 437112 582632 437164 582684
rect 24124 582564 24176 582616
rect 449808 582564 449860 582616
rect 5172 582496 5224 582548
rect 434996 582496 435048 582548
rect 3700 582428 3752 582480
rect 443460 582428 443512 582480
rect 5080 582360 5132 582412
rect 447692 582360 447744 582412
rect 302424 581544 302476 581596
rect 469588 581544 469640 581596
rect 296076 581476 296128 581528
rect 469680 581476 469732 581528
rect 289728 581408 289780 581460
rect 470508 581408 470560 581460
rect 287612 581340 287664 581392
rect 470416 581340 470468 581392
rect 283472 581272 283524 581324
rect 470324 581272 470376 581324
rect 281356 581204 281408 581256
rect 470140 581204 470192 581256
rect 275008 581136 275060 581188
rect 470048 581136 470100 581188
rect 264520 581068 264572 581120
rect 580908 581068 580960 581120
rect 258172 581000 258224 581052
rect 580632 581000 580684 581052
rect 268660 580252 268712 580304
rect 469864 580252 469916 580304
rect 306564 580184 306616 580236
rect 580172 580184 580224 580236
rect 6736 580116 6788 580168
rect 395068 580116 395120 580168
rect 6460 580048 6512 580100
rect 401324 580048 401376 580100
rect 6276 579980 6328 580032
rect 414112 579980 414164 580032
rect 3976 579912 4028 579964
rect 426440 579912 426492 579964
rect 3792 579844 3844 579896
rect 438860 579844 438912 579896
rect 4988 579776 5040 579828
rect 451556 579776 451608 579828
rect 4896 579708 4948 579760
rect 458272 579708 458324 579760
rect 6184 579640 6236 579692
rect 464252 579640 464304 579692
rect 271144 579368 271196 579420
rect 254124 579300 254176 579352
rect 260656 579300 260708 579352
rect 266820 579300 266872 579352
rect 273168 579300 273220 579352
rect 277308 579300 277360 579352
rect 279608 579300 279660 579352
rect 285772 579300 285824 579352
rect 292120 579343 292172 579352
rect 292120 579309 292129 579343
rect 292129 579309 292163 579343
rect 292163 579309 292172 579343
rect 292120 579300 292172 579309
rect 396724 579343 396776 579352
rect 396724 579309 396733 579343
rect 396733 579309 396767 579343
rect 396767 579309 396776 579343
rect 396724 579300 396776 579309
rect 415676 579343 415728 579352
rect 415676 579309 415685 579343
rect 415685 579309 415719 579343
rect 415719 579309 415728 579343
rect 415676 579300 415728 579309
rect 428372 579343 428424 579352
rect 428372 579309 428381 579343
rect 428381 579309 428415 579343
rect 428415 579309 428424 579343
rect 428372 579300 428424 579309
rect 441068 579343 441120 579352
rect 441068 579309 441077 579343
rect 441077 579309 441111 579343
rect 441111 579309 441120 579343
rect 441068 579300 441120 579309
rect 453580 579343 453632 579352
rect 453580 579309 453589 579343
rect 453589 579309 453623 579343
rect 453623 579309 453632 579343
rect 453580 579300 453632 579309
rect 455788 579343 455840 579352
rect 455788 579309 455797 579343
rect 455797 579309 455831 579343
rect 455831 579309 455840 579343
rect 455788 579300 455840 579309
rect 470232 579164 470284 579216
rect 469956 579096 470008 579148
rect 579896 579028 579948 579080
rect 580080 578960 580132 579012
rect 579988 578892 580040 578944
rect 580172 578824 580224 578876
rect 580816 578756 580868 578808
rect 580540 578688 580592 578740
rect 580264 578620 580316 578672
rect 6552 578552 6604 578604
rect 3332 578484 3384 578536
rect 3884 578416 3936 578468
rect 3608 578348 3660 578400
rect 3424 578280 3476 578332
rect 3516 578212 3568 578264
rect 3148 568284 3200 568336
rect 6736 568284 6788 568336
rect 579804 567128 579856 567180
rect 580908 567128 580960 567180
rect 579804 557608 579856 557660
rect 580908 557540 580960 557592
rect 469588 557472 469640 557524
rect 579804 557472 579856 557524
rect 3148 553324 3200 553376
rect 6644 553324 6696 553376
rect 579712 547816 579764 547868
rect 580908 547816 580960 547868
rect 471244 546388 471296 546440
rect 579804 546388 579856 546440
rect 3056 539044 3108 539096
rect 6552 539044 6604 539096
rect 579712 538228 579764 538280
rect 580908 538228 580960 538280
rect 579804 528504 579856 528556
rect 580908 528504 580960 528556
rect 579804 518916 579856 518968
rect 580908 518916 580960 518968
rect 469680 510552 469732 510604
rect 579804 510552 579856 510604
rect 3148 510212 3200 510264
rect 6460 510212 6512 510264
rect 579804 509192 579856 509244
rect 580908 509192 580960 509244
rect 579804 499604 579856 499656
rect 580908 499536 580960 499588
rect 469772 499468 469824 499520
rect 579804 499468 579856 499520
rect 2780 495728 2832 495780
rect 4712 495728 4764 495780
rect 579804 489812 579856 489864
rect 580908 489812 580960 489864
rect 3148 481244 3200 481296
rect 6368 481244 6420 481296
rect 579804 480224 579856 480276
rect 580908 480224 580960 480276
rect 579712 470500 579764 470552
rect 580908 470500 580960 470552
rect 470508 463632 470560 463684
rect 579804 463632 579856 463684
rect 579712 460912 579764 460964
rect 580908 460912 580960 460964
rect 470416 440172 470468 440224
rect 579896 440172 579948 440224
rect 2780 438540 2832 438592
rect 5448 438540 5500 438592
rect 2780 424804 2832 424856
rect 5356 424804 5408 424856
rect 470324 416712 470376 416764
rect 579896 416712 579948 416764
rect 579804 412564 579856 412616
rect 580908 412564 580960 412616
rect 470232 405628 470284 405680
rect 579896 405628 579948 405680
rect 579804 402976 579856 403028
rect 580908 402976 580960 403028
rect 3240 395836 3292 395888
rect 6276 395836 6328 395888
rect 470140 393252 470192 393304
rect 579896 393252 579948 393304
rect 579804 393184 579856 393236
rect 580908 393252 580960 393304
rect 579804 384276 579856 384328
rect 580908 384276 580960 384328
rect 2780 380740 2832 380792
rect 5264 380740 5316 380792
rect 579988 361224 580040 361276
rect 580908 361224 580960 361276
rect 579804 360136 579856 360188
rect 579988 360136 580040 360188
rect 470048 346332 470100 346384
rect 579804 346332 579856 346384
rect 580080 345040 580132 345092
rect 580908 345040 580960 345092
rect 580080 344904 580132 344956
rect 580908 344904 580960 344956
rect 341616 338784 341668 338836
rect 348516 338648 348568 338700
rect 327356 338376 327408 338428
rect 327908 338376 327960 338428
rect 79324 338036 79376 338088
rect 257896 338036 257948 338088
rect 309784 338036 309836 338088
rect 354404 338036 354456 338088
rect 358084 338036 358136 338088
rect 371516 338036 371568 338088
rect 378876 338036 378928 338088
rect 411260 338036 411312 338088
rect 412456 338036 412508 338088
rect 414664 338036 414716 338088
rect 429844 338036 429896 338088
rect 435732 338036 435784 338088
rect 499580 338036 499632 338088
rect 71044 337968 71096 338020
rect 252008 337968 252060 338020
rect 306196 337968 306248 338020
rect 355876 337968 355928 338020
rect 364248 337968 364300 338020
rect 379336 337968 379388 338020
rect 399484 337968 399536 338020
rect 400128 337968 400180 338020
rect 403348 337968 403400 338020
rect 415124 337968 415176 338020
rect 420276 337968 420328 338020
rect 420552 337968 420604 338020
rect 440148 338011 440200 338020
rect 440148 337977 440157 338011
rect 440157 337977 440191 338011
rect 440191 337977 440200 338011
rect 440148 337968 440200 337977
rect 454776 337968 454828 338020
rect 527824 337968 527876 338020
rect 66904 337900 66956 337952
rect 247132 337900 247184 337952
rect 303160 337900 303212 337952
rect 352932 337900 352984 337952
rect 355324 337900 355376 337952
rect 370044 337900 370096 337952
rect 371148 337900 371200 337952
rect 382280 337900 382332 337952
rect 409236 337900 409288 337952
rect 416044 337900 416096 337952
rect 416596 337900 416648 337952
rect 421564 337900 421616 337952
rect 422024 337900 422076 337952
rect 438124 337900 438176 337952
rect 438676 337900 438728 337952
rect 449164 337900 449216 337952
rect 450452 337900 450504 337952
rect 451188 337900 451240 337952
rect 451832 337900 451884 337952
rect 61384 337832 61436 337884
rect 247592 337832 247644 337884
rect 258816 337832 258868 337884
rect 272616 337832 272668 337884
rect 317420 337832 317472 337884
rect 326988 337832 327040 337884
rect 336096 337832 336148 337884
rect 344560 337832 344612 337884
rect 349988 337832 350040 337884
rect 57244 337764 57296 337816
rect 244188 337764 244240 337816
rect 259644 337764 259696 337816
rect 260104 337764 260156 337816
rect 288256 337764 288308 337816
rect 35164 337696 35216 337748
rect 238300 337696 238352 337748
rect 254584 337696 254636 337748
rect 262312 337696 262364 337748
rect 351920 337764 351972 337816
rect 327172 337696 327224 337748
rect 336188 337696 336240 337748
rect 39304 337628 39356 337680
rect 244648 337628 244700 337680
rect 260104 337628 260156 337680
rect 277032 337628 277084 337680
rect 285588 337628 285640 337680
rect 347044 337628 347096 337680
rect 348424 337628 348476 337680
rect 365628 337832 365680 337884
rect 380808 337832 380860 337884
rect 388444 337832 388496 337884
rect 389180 337832 389232 337884
rect 397460 337832 397512 337884
rect 399484 337832 399536 337884
rect 399944 337832 399996 337884
rect 412824 337832 412876 337884
rect 413652 337832 413704 337884
rect 417424 337832 417476 337884
rect 417608 337832 417660 337884
rect 455604 337832 455656 337884
rect 458732 337832 458784 337884
rect 459376 337832 459428 337884
rect 460664 337832 460716 337884
rect 525064 337900 525116 337952
rect 523684 337832 523736 337884
rect 358728 337764 358780 337816
rect 356704 337628 356756 337680
rect 360752 337628 360804 337680
rect 362868 337764 362920 337816
rect 361672 337696 361724 337748
rect 362316 337696 362368 337748
rect 363052 337696 363104 337748
rect 363788 337696 363840 337748
rect 377404 337764 377456 337816
rect 398012 337764 398064 337816
rect 399576 337764 399628 337816
rect 401876 337764 401928 337816
rect 416964 337764 417016 337816
rect 420000 337764 420052 337816
rect 420736 337764 420788 337816
rect 424968 337764 425020 337816
rect 442264 337764 442316 337816
rect 444564 337764 444616 337816
rect 445668 337764 445720 337816
rect 446036 337764 446088 337816
rect 453304 337764 453356 337816
rect 453948 337764 454000 337816
rect 463792 337764 463844 337816
rect 465632 337764 465684 337816
rect 466184 337764 466236 337816
rect 467104 337764 467156 337816
rect 467748 337764 467800 337816
rect 468024 337764 468076 337816
rect 469036 337764 469088 337816
rect 521016 337764 521068 337816
rect 375932 337696 375984 337748
rect 380164 337696 380216 337748
rect 381360 337696 381412 337748
rect 381544 337696 381596 337748
rect 382832 337696 382884 337748
rect 384948 337696 385000 337748
rect 388168 337696 388220 337748
rect 408776 337696 408828 337748
rect 409788 337696 409840 337748
rect 32404 337560 32456 337612
rect 241704 337560 241756 337612
rect 252192 337560 252244 337612
rect 256424 337560 256476 337612
rect 261392 337560 261444 337612
rect 279976 337560 280028 337612
rect 281448 337560 281500 337612
rect 345296 337560 345348 337612
rect 351460 337560 351512 337612
rect 351644 337560 351696 337612
rect 369124 337560 369176 337612
rect 371056 337560 371108 337612
rect 28264 337492 28316 337544
rect 19984 337424 20036 337476
rect 234344 337424 234396 337476
rect 253204 337492 253256 337544
rect 259368 337492 259420 337544
rect 237840 337424 237892 337476
rect 258724 337424 258776 337476
rect 275560 337492 275612 337544
rect 275928 337492 275980 337544
rect 342904 337492 342956 337544
rect 353392 337492 353444 337544
rect 357348 337492 357400 337544
rect 359464 337492 359516 337544
rect 363696 337492 363748 337544
rect 13084 337356 13136 337408
rect 233516 337356 233568 337408
rect 233884 337356 233936 337408
rect 241244 337356 241296 337408
rect 247684 337356 247736 337408
rect 248604 337356 248656 337408
rect 249064 337356 249116 337408
rect 250536 337356 250588 337408
rect 250720 337356 250772 337408
rect 253480 337356 253532 337408
rect 257344 337356 257396 337408
rect 269672 337424 269724 337476
rect 297916 337424 297968 337476
rect 314660 337424 314712 337476
rect 315396 337424 315448 337476
rect 316132 337424 316184 337476
rect 316316 337424 316368 337476
rect 317420 337424 317472 337476
rect 318340 337424 318392 337476
rect 318892 337424 318944 337476
rect 319260 337424 319312 337476
rect 320180 337424 320232 337476
rect 320732 337424 320784 337476
rect 338764 337424 338816 337476
rect 347504 337424 347556 337476
rect 349068 337424 349120 337476
rect 372988 337424 373040 337476
rect 77944 337288 77996 337340
rect 84844 337288 84896 337340
rect 260840 337288 260892 337340
rect 132500 337220 132552 337272
rect 142068 337220 142120 337272
rect 151820 337220 151872 337272
rect 161388 337220 161440 337272
rect 171140 337220 171192 337272
rect 180708 337220 180760 337272
rect 190460 337220 190512 337272
rect 200028 337220 200080 337272
rect 209780 337220 209832 337272
rect 219348 337220 219400 337272
rect 229192 337220 229244 337272
rect 234620 337220 234672 337272
rect 254952 337220 255004 337272
rect 255964 337220 256016 337272
rect 266728 337356 266780 337408
rect 269028 337356 269080 337408
rect 340236 337356 340288 337408
rect 340788 337356 340840 337408
rect 369584 337356 369636 337408
rect 369768 337356 369820 337408
rect 381820 337628 381872 337680
rect 384304 337628 384356 337680
rect 387708 337628 387760 337680
rect 404360 337628 404412 337680
rect 419540 337696 419592 337748
rect 420828 337696 420880 337748
rect 421472 337696 421524 337748
rect 422208 337696 422260 337748
rect 422484 337696 422536 337748
rect 424416 337696 424468 337748
rect 425428 337696 425480 337748
rect 428464 337696 428516 337748
rect 439136 337696 439188 337748
rect 440148 337696 440200 337748
rect 506480 337696 506532 337748
rect 420184 337628 420236 337680
rect 427912 337628 427964 337680
rect 442080 337628 442132 337680
rect 442908 337628 442960 337680
rect 443552 337628 443604 337680
rect 444288 337628 444340 337680
rect 445024 337628 445076 337680
rect 445576 337628 445628 337680
rect 446496 337628 446548 337680
rect 447048 337628 447100 337680
rect 448244 337628 448296 337680
rect 448428 337628 448480 337680
rect 449900 337628 449952 337680
rect 451004 337628 451056 337680
rect 451372 337628 451424 337680
rect 452476 337628 452528 337680
rect 452844 337628 452896 337680
rect 453764 337628 453816 337680
rect 454316 337628 454368 337680
rect 455236 337628 455288 337680
rect 455788 337628 455840 337680
rect 456616 337628 456668 337680
rect 456800 337628 456852 337680
rect 458088 337628 458140 337680
rect 458180 337628 458232 337680
rect 520924 337628 520976 337680
rect 373908 337560 373960 337612
rect 383292 337560 383344 337612
rect 404820 337560 404872 337612
rect 415584 337560 415636 337612
rect 416596 337560 416648 337612
rect 400404 337492 400456 337544
rect 406384 337492 406436 337544
rect 407304 337492 407356 337544
rect 375288 337424 375340 337476
rect 383752 337424 383804 337476
rect 387064 337424 387116 337476
rect 388720 337424 388772 337476
rect 398472 337424 398524 337476
rect 382188 337356 382240 337408
rect 386696 337356 386748 337408
rect 400956 337356 401008 337408
rect 402244 337356 402296 337408
rect 405832 337424 405884 337476
rect 426440 337424 426492 337476
rect 430120 337560 430172 337612
rect 436652 337560 436704 337612
rect 437296 337560 437348 337612
rect 437664 337560 437716 337612
rect 438676 337560 438728 337612
rect 440608 337560 440660 337612
rect 441528 337560 441580 337612
rect 441620 337560 441672 337612
rect 443644 337560 443696 337612
rect 427176 337492 427228 337544
rect 437204 337492 437256 337544
rect 442356 337492 442408 337544
rect 408684 337356 408736 337408
rect 411720 337356 411772 337408
rect 434260 337424 434312 337476
rect 439504 337424 439556 337476
rect 447508 337492 447560 337544
rect 448428 337492 448480 337544
rect 443092 337424 443144 337476
rect 448980 337560 449032 337612
rect 518164 337560 518216 337612
rect 514024 337492 514076 337544
rect 516784 337424 516836 337476
rect 510620 337356 510672 337408
rect 272800 337288 272852 337340
rect 314200 337288 314252 337340
rect 316040 337288 316092 337340
rect 316868 337288 316920 337340
rect 318800 337288 318852 337340
rect 319812 337288 319864 337340
rect 321468 337288 321520 337340
rect 361764 337288 361816 337340
rect 366916 337288 366968 337340
rect 380348 337288 380400 337340
rect 397000 337288 397052 337340
rect 405924 337288 405976 337340
rect 412732 337288 412784 337340
rect 413836 337288 413888 337340
rect 418528 337288 418580 337340
rect 419448 337288 419500 337340
rect 421012 337288 421064 337340
rect 470600 337288 470652 337340
rect 470692 337288 470744 337340
rect 529204 337288 529256 337340
rect 271328 337220 271380 337272
rect 312452 337220 312504 337272
rect 312544 337220 312596 337272
rect 350448 337220 350500 337272
rect 355968 337220 356020 337272
rect 414204 337220 414256 337272
rect 415308 337220 415360 337272
rect 423496 337220 423548 337272
rect 463608 337220 463660 337272
rect 469496 337220 469548 337272
rect 530584 337220 530636 337272
rect 97264 337152 97316 337204
rect 268200 337152 268252 337204
rect 271788 337152 271840 337204
rect 333244 337152 333296 337204
rect 366640 337152 366692 337204
rect 372068 337152 372120 337204
rect 424324 337152 424376 337204
rect 100668 337084 100720 337136
rect 271144 337084 271196 337136
rect 316684 337084 316736 337136
rect 341892 337084 341944 337136
rect 348976 337084 349028 337136
rect 351828 337084 351880 337136
rect 374460 337084 374512 337136
rect 406292 337084 406344 337136
rect 411904 337084 411956 337136
rect 417056 337084 417108 337136
rect 417976 337084 418028 337136
rect 419080 337084 419132 337136
rect 431500 337152 431552 337204
rect 434076 337152 434128 337204
rect 427084 337084 427136 337136
rect 432788 337084 432840 337136
rect 492680 337152 492732 337204
rect 485780 337084 485832 337136
rect 95884 337016 95936 337068
rect 263784 337016 263836 337068
rect 335268 337016 335320 337068
rect 367652 337016 367704 337068
rect 393596 337016 393648 337068
rect 397460 337016 397512 337068
rect 401416 337016 401468 337068
rect 405004 337016 405056 337068
rect 421104 337016 421156 337068
rect 444380 337016 444432 337068
rect 444748 337016 444800 337068
rect 477592 337016 477644 337068
rect 107568 336948 107620 337000
rect 274088 336948 274140 337000
rect 319444 336948 319496 337000
rect 378048 336948 378100 337000
rect 385224 336948 385276 337000
rect 398932 336948 398984 337000
rect 403624 336948 403676 337000
rect 407764 336948 407816 337000
rect 102784 336880 102836 336932
rect 265256 336880 265308 336932
rect 284300 336880 284352 336932
rect 284852 336880 284904 336932
rect 327724 336880 327776 336932
rect 345480 336880 345532 336932
rect 345664 336880 345716 336932
rect 360292 336880 360344 336932
rect 380808 336880 380860 336932
rect 386236 336880 386288 336932
rect 392124 336880 392176 336932
rect 393596 336880 393648 336932
rect 410248 336880 410300 336932
rect 411168 336880 411220 336932
rect 426808 336948 426860 337000
rect 475384 336948 475436 337000
rect 413284 336880 413336 336932
rect 444380 336880 444432 336932
rect 118608 336812 118660 336864
rect 278504 336812 278556 336864
rect 343088 336812 343140 336864
rect 344284 336812 344336 336864
rect 351184 336812 351236 336864
rect 351644 336812 351696 336864
rect 125508 336744 125560 336796
rect 281172 336744 281224 336796
rect 290464 336744 290516 336796
rect 344100 336744 344152 336796
rect 344376 336744 344428 336796
rect 354864 336812 354916 336864
rect 362224 336812 362276 336864
rect 365168 336812 365220 336864
rect 381636 336812 381688 336864
rect 384764 336812 384816 336864
rect 396080 336812 396132 336864
rect 398104 336812 398156 336864
rect 423956 336812 424008 336864
rect 428372 336812 428424 336864
rect 431224 336812 431276 336864
rect 431316 336812 431368 336864
rect 433984 336812 434036 336864
rect 434720 336812 434772 336864
rect 435916 336812 435968 336864
rect 352564 336744 352616 336796
rect 357808 336744 357860 336796
rect 363604 336744 363656 336796
rect 364708 336744 364760 336796
rect 370504 336744 370556 336796
rect 372528 336744 372580 336796
rect 376024 336744 376076 336796
rect 376944 336744 376996 336796
rect 377680 336744 377732 336796
rect 378416 336744 378468 336796
rect 392584 336744 392636 336796
rect 393228 336744 393280 336796
rect 394056 336744 394108 336796
rect 394608 336744 394660 336796
rect 395068 336744 395120 336796
rect 395896 336744 395948 336796
rect 396540 336744 396592 336796
rect 398196 336744 398248 336796
rect 429384 336744 429436 336796
rect 430396 336744 430448 336796
rect 430856 336744 430908 336796
rect 431776 336744 431828 336796
rect 432328 336744 432380 336796
rect 433156 336744 433208 336796
rect 433708 336744 433760 336796
rect 434628 336744 434680 336796
rect 435180 336744 435232 336796
rect 436008 336744 436060 336796
rect 436192 336744 436244 336796
rect 437388 336744 437440 336796
rect 444380 336744 444432 336796
rect 459192 336880 459244 336932
rect 460296 336880 460348 336932
rect 461676 336880 461728 336932
rect 465080 336880 465132 336932
rect 466368 336880 466420 336932
rect 466552 336880 466604 336932
rect 470508 336880 470560 336932
rect 459652 336812 459704 336864
rect 460204 336812 460256 336864
rect 460756 336812 460808 336864
rect 469220 336812 469272 336864
rect 457260 336744 457312 336796
rect 457996 336744 458048 336796
rect 458272 336744 458324 336796
rect 459468 336744 459520 336796
rect 459744 336744 459796 336796
rect 460848 336744 460900 336796
rect 461216 336744 461268 336796
rect 462136 336744 462188 336796
rect 462688 336744 462740 336796
rect 463516 336744 463568 336796
rect 464160 336744 464212 336796
rect 464988 336744 465040 336796
rect 509884 336812 509936 336864
rect 323676 336676 323728 336728
rect 464896 336676 464948 336728
rect 505744 336744 505796 336796
rect 236184 335656 236236 335708
rect 237012 335656 237064 335708
rect 302240 335656 302292 335708
rect 302700 335656 302752 335708
rect 331312 335656 331364 335708
rect 331956 335656 332008 335708
rect 334072 335656 334124 335708
rect 334900 335656 334952 335708
rect 236092 335588 236144 335640
rect 236552 335588 236604 335640
rect 241612 335588 241664 335640
rect 242348 335588 242400 335640
rect 260932 335588 260984 335640
rect 261484 335588 261536 335640
rect 262588 335588 262640 335640
rect 263048 335588 263100 335640
rect 263692 335588 263744 335640
rect 264428 335588 264480 335640
rect 265072 335588 265124 335640
rect 265900 335588 265952 335640
rect 266452 335588 266504 335640
rect 267372 335588 267424 335640
rect 280252 335588 280304 335640
rect 280620 335588 280672 335640
rect 283012 335588 283064 335640
rect 283564 335588 283616 335640
rect 285680 335588 285732 335640
rect 285956 335588 286008 335640
rect 287060 335588 287112 335640
rect 287980 335588 288032 335640
rect 288440 335588 288492 335640
rect 289452 335588 289504 335640
rect 292764 335588 292816 335640
rect 293316 335588 293368 335640
rect 298284 335588 298336 335640
rect 298652 335588 298704 335640
rect 300860 335588 300912 335640
rect 301228 335588 301280 335640
rect 303620 335588 303672 335640
rect 304172 335588 304224 335640
rect 305000 335588 305052 335640
rect 305644 335588 305696 335640
rect 307760 335588 307812 335640
rect 308588 335588 308640 335640
rect 309140 335588 309192 335640
rect 310060 335588 310112 335640
rect 310520 335588 310572 335640
rect 311532 335588 311584 335640
rect 321652 335588 321704 335640
rect 322204 335588 322256 335640
rect 329840 335588 329892 335640
rect 330116 335588 330168 335640
rect 331220 335588 331272 335640
rect 331588 335588 331640 335640
rect 332600 335588 332652 335640
rect 333060 335588 333112 335640
rect 333980 335588 334032 335640
rect 334532 335588 334584 335640
rect 338120 335588 338172 335640
rect 338948 335588 339000 335640
rect 356152 335588 356204 335640
rect 356612 335588 356664 335640
rect 359004 335588 359056 335640
rect 359372 335588 359424 335640
rect 250628 335520 250680 335572
rect 248512 335452 248564 335504
rect 249156 335452 249208 335504
rect 285956 335452 286008 335504
rect 286600 335452 286652 335504
rect 278872 335384 278924 335436
rect 580080 335384 580132 335436
rect 581000 335384 581052 335436
rect 367284 335316 367336 335368
rect 367928 335316 367980 335368
rect 580080 335248 580132 335300
rect 581000 335248 581052 335300
rect 278964 335180 279016 335232
rect 332692 335044 332744 335096
rect 333428 335044 333480 335096
rect 302516 334704 302568 334756
rect 303068 334704 303120 334756
rect 258172 334568 258224 334620
rect 258540 334568 258592 334620
rect 270776 334296 270828 334348
rect 271236 334296 271288 334348
rect 272248 334296 272300 334348
rect 272708 334296 272760 334348
rect 335360 333888 335412 333940
rect 336004 333888 336056 333940
rect 278872 333276 278924 333328
rect 279056 333276 279108 333328
rect 306472 333276 306524 333328
rect 306656 333276 306708 333328
rect 242992 332052 243044 332104
rect 243452 332052 243504 332104
rect 331404 331891 331456 331900
rect 331404 331857 331413 331891
rect 331413 331857 331447 331891
rect 331447 331857 331456 331891
rect 331404 331848 331456 331857
rect 336740 331848 336792 331900
rect 336924 331848 336976 331900
rect 328552 331644 328604 331696
rect 329012 331644 329064 331696
rect 341432 331304 341484 331356
rect 341708 331304 341760 331356
rect 299572 331236 299624 331288
rect 259644 331168 259696 331220
rect 259828 331168 259880 331220
rect 262588 331168 262640 331220
rect 262772 331168 262824 331220
rect 303896 331168 303948 331220
rect 304632 331168 304684 331220
rect 389272 331168 389324 331220
rect 389456 331168 389508 331220
rect 459652 331168 459704 331220
rect 460112 331168 460164 331220
rect 299572 331100 299624 331152
rect 299756 331100 299808 331152
rect 300308 331100 300360 331152
rect 299480 331032 299532 331084
rect 299664 331032 299716 331084
rect 301136 328448 301188 328500
rect 301688 328448 301740 328500
rect 339776 328448 339828 328500
rect 340328 328448 340380 328500
rect 367008 328448 367060 328500
rect 372712 328448 372764 328500
rect 373080 328448 373132 328500
rect 259828 328423 259880 328432
rect 259828 328389 259837 328423
rect 259837 328389 259871 328423
rect 259871 328389 259880 328423
rect 259828 328380 259880 328389
rect 265256 328380 265308 328432
rect 265348 328380 265400 328432
rect 294236 328380 294288 328432
rect 294420 328380 294472 328432
rect 295524 328380 295576 328432
rect 295708 328380 295760 328432
rect 296812 328380 296864 328432
rect 296996 328380 297048 328432
rect 341340 328423 341392 328432
rect 341340 328389 341349 328423
rect 341349 328389 341383 328423
rect 341383 328389 341392 328423
rect 341340 328380 341392 328389
rect 389456 328423 389508 328432
rect 389456 328389 389465 328423
rect 389465 328389 389499 328423
rect 389499 328389 389508 328423
rect 389456 328380 389508 328389
rect 393596 328380 393648 328432
rect 393688 328380 393740 328432
rect 367008 328355 367060 328364
rect 367008 328321 367017 328355
rect 367017 328321 367051 328355
rect 367051 328321 367060 328355
rect 367008 328312 367060 328321
rect 337016 327156 337068 327208
rect 250168 327131 250220 327140
rect 250168 327097 250177 327131
rect 250177 327097 250211 327131
rect 250211 327097 250220 327131
rect 250168 327088 250220 327097
rect 323308 327131 323360 327140
rect 323308 327097 323317 327131
rect 323317 327097 323351 327131
rect 323351 327097 323360 327131
rect 323308 327088 323360 327097
rect 324688 327088 324740 327140
rect 325056 327088 325108 327140
rect 325976 327088 326028 327140
rect 326620 327088 326672 327140
rect 336832 327088 336884 327140
rect 265348 327020 265400 327072
rect 301136 327020 301188 327072
rect 327264 327063 327316 327072
rect 327264 327029 327273 327063
rect 327273 327029 327307 327063
rect 327307 327029 327316 327063
rect 327264 327020 327316 327029
rect 288716 325660 288768 325712
rect 288808 325660 288860 325712
rect 580080 325660 580132 325712
rect 580908 325660 580960 325712
rect 3332 324232 3384 324284
rect 14464 324232 14516 324284
rect 469956 322872 470008 322924
rect 580080 322872 580132 322924
rect 273536 321759 273588 321768
rect 273536 321725 273545 321759
rect 273545 321725 273579 321759
rect 273579 321725 273588 321759
rect 273536 321716 273588 321725
rect 262772 321580 262824 321632
rect 266728 321580 266780 321632
rect 267832 321580 267884 321632
rect 281816 321580 281868 321632
rect 310796 321580 310848 321632
rect 375840 321580 375892 321632
rect 377128 321580 377180 321632
rect 230756 321512 230808 321564
rect 230940 321512 230992 321564
rect 232228 321512 232280 321564
rect 232412 321512 232464 321564
rect 262864 321444 262916 321496
rect 310888 321444 310940 321496
rect 375932 321376 375984 321428
rect 377220 321376 377272 321428
rect 331404 318903 331456 318912
rect 331404 318869 331413 318903
rect 331413 318869 331447 318903
rect 331447 318869 331456 318903
rect 331404 318860 331456 318869
rect 259920 318792 259972 318844
rect 266636 318835 266688 318844
rect 266636 318801 266645 318835
rect 266645 318801 266679 318835
rect 266679 318801 266688 318835
rect 266636 318792 266688 318801
rect 267740 318835 267792 318844
rect 267740 318801 267749 318835
rect 267749 318801 267783 318835
rect 267783 318801 267792 318835
rect 267740 318792 267792 318801
rect 299756 318792 299808 318844
rect 299848 318792 299900 318844
rect 302516 318792 302568 318844
rect 302608 318792 302660 318844
rect 306748 318792 306800 318844
rect 306840 318792 306892 318844
rect 341432 318792 341484 318844
rect 357624 318792 357676 318844
rect 357716 318792 357768 318844
rect 367008 318835 367060 318844
rect 367008 318801 367017 318835
rect 367017 318801 367051 318835
rect 367051 318801 367060 318835
rect 367008 318792 367060 318801
rect 389548 318792 389600 318844
rect 431408 318792 431460 318844
rect 431500 318792 431552 318844
rect 230940 318724 230992 318776
rect 235080 318767 235132 318776
rect 235080 318733 235089 318767
rect 235089 318733 235123 318767
rect 235123 318733 235132 318767
rect 235080 318724 235132 318733
rect 236276 318767 236328 318776
rect 236276 318733 236285 318767
rect 236285 318733 236319 318767
rect 236319 318733 236328 318767
rect 236276 318724 236328 318733
rect 372712 318767 372764 318776
rect 372712 318733 372721 318767
rect 372721 318733 372755 318767
rect 372755 318733 372764 318767
rect 372712 318724 372764 318733
rect 273536 317543 273588 317552
rect 273536 317509 273545 317543
rect 273545 317509 273579 317543
rect 273579 317509 273588 317543
rect 273536 317500 273588 317509
rect 265256 317475 265308 317484
rect 265256 317441 265265 317475
rect 265265 317441 265299 317475
rect 265299 317441 265308 317475
rect 265256 317432 265308 317441
rect 301044 317475 301096 317484
rect 301044 317441 301053 317475
rect 301053 317441 301087 317475
rect 301087 317441 301096 317475
rect 301044 317432 301096 317441
rect 327264 317475 327316 317484
rect 327264 317441 327273 317475
rect 327273 317441 327307 317475
rect 327307 317441 327316 317475
rect 327264 317432 327316 317441
rect 250168 317407 250220 317416
rect 250168 317373 250177 317407
rect 250177 317373 250211 317407
rect 250211 317373 250220 317407
rect 250168 317364 250220 317373
rect 251548 317407 251600 317416
rect 251548 317373 251557 317407
rect 251557 317373 251591 317407
rect 251591 317373 251600 317407
rect 251548 317364 251600 317373
rect 270776 317407 270828 317416
rect 270776 317373 270785 317407
rect 270785 317373 270819 317407
rect 270819 317373 270828 317407
rect 270776 317364 270828 317373
rect 272248 317407 272300 317416
rect 272248 317373 272257 317407
rect 272257 317373 272291 317407
rect 272291 317373 272300 317407
rect 272248 317364 272300 317373
rect 273536 317364 273588 317416
rect 290096 317364 290148 317416
rect 290188 317364 290240 317416
rect 291568 317364 291620 317416
rect 291660 317364 291712 317416
rect 296904 317364 296956 317416
rect 296996 317364 297048 317416
rect 306840 317407 306892 317416
rect 306840 317373 306849 317407
rect 306849 317373 306883 317407
rect 306883 317373 306892 317407
rect 306840 317364 306892 317373
rect 330208 317407 330260 317416
rect 330208 317373 330217 317407
rect 330217 317373 330251 317407
rect 330251 317373 330260 317407
rect 330208 317364 330260 317373
rect 331404 317407 331456 317416
rect 331404 317373 331413 317407
rect 331413 317373 331447 317407
rect 331447 317373 331456 317407
rect 331404 317364 331456 317373
rect 393596 317407 393648 317416
rect 393596 317373 393605 317407
rect 393605 317373 393639 317407
rect 393639 317373 393648 317407
rect 393596 317364 393648 317373
rect 460204 317407 460256 317416
rect 460204 317373 460213 317407
rect 460213 317373 460247 317407
rect 460247 317373 460256 317407
rect 460204 317364 460256 317373
rect 273628 317296 273680 317348
rect 579988 316072 580040 316124
rect 581000 316072 581052 316124
rect 281724 316047 281776 316056
rect 281724 316013 281733 316047
rect 281733 316013 281767 316047
rect 281767 316013 281776 316047
rect 281724 316004 281776 316013
rect 285772 316004 285824 316056
rect 286048 316004 286100 316056
rect 267740 315979 267792 315988
rect 267740 315945 267749 315979
rect 267749 315945 267783 315979
rect 267783 315945 267792 315979
rect 267740 315936 267792 315945
rect 580080 315936 580132 315988
rect 581000 315936 581052 315988
rect 250168 312579 250220 312588
rect 250168 312545 250177 312579
rect 250177 312545 250211 312579
rect 250211 312545 250220 312579
rect 250168 312536 250220 312545
rect 232412 311924 232464 311976
rect 244372 311924 244424 311976
rect 245844 311924 245896 311976
rect 284760 311924 284812 311976
rect 232320 311788 232372 311840
rect 235080 311831 235132 311840
rect 235080 311797 235089 311831
rect 235089 311797 235123 311831
rect 235123 311797 235132 311831
rect 235080 311788 235132 311797
rect 244464 311720 244516 311772
rect 259736 311856 259788 311908
rect 259920 311856 259972 311908
rect 299848 311924 299900 311976
rect 302608 311924 302660 311976
rect 310888 311967 310940 311976
rect 310888 311933 310897 311967
rect 310897 311933 310931 311967
rect 310931 311933 310940 311967
rect 310888 311924 310940 311933
rect 323308 311924 323360 311976
rect 337108 311967 337160 311976
rect 337108 311933 337117 311967
rect 337117 311933 337151 311967
rect 337151 311933 337160 311967
rect 337108 311924 337160 311933
rect 431408 311924 431460 311976
rect 431500 311924 431552 311976
rect 323216 311856 323268 311908
rect 341248 311856 341300 311908
rect 341432 311856 341484 311908
rect 389364 311856 389416 311908
rect 389548 311856 389600 311908
rect 284760 311788 284812 311840
rect 299756 311788 299808 311840
rect 302516 311788 302568 311840
rect 245936 311720 245988 311772
rect 239128 311652 239180 311704
rect 239128 311516 239180 311568
rect 267832 311108 267884 311160
rect 266636 309247 266688 309256
rect 266636 309213 266645 309247
rect 266645 309213 266679 309247
rect 266679 309213 266688 309247
rect 266636 309204 266688 309213
rect 230848 309179 230900 309188
rect 230848 309145 230857 309179
rect 230857 309145 230891 309179
rect 230891 309145 230900 309179
rect 230848 309136 230900 309145
rect 236276 309179 236328 309188
rect 236276 309145 236285 309179
rect 236285 309145 236319 309179
rect 236319 309145 236328 309179
rect 236276 309136 236328 309145
rect 327172 309136 327224 309188
rect 372712 309179 372764 309188
rect 372712 309145 372721 309179
rect 372721 309145 372755 309179
rect 372755 309145 372764 309179
rect 372712 309136 372764 309145
rect 265256 309111 265308 309120
rect 265256 309077 265265 309111
rect 265265 309077 265299 309111
rect 265299 309077 265308 309111
rect 265256 309068 265308 309077
rect 337200 309068 337252 309120
rect 341248 309068 341300 309120
rect 367008 309111 367060 309120
rect 367008 309077 367017 309111
rect 367017 309077 367051 309111
rect 367051 309077 367060 309111
rect 367008 309068 367060 309077
rect 327172 309000 327224 309052
rect 310704 307844 310756 307896
rect 251548 307819 251600 307828
rect 251548 307785 251557 307819
rect 251557 307785 251591 307819
rect 251591 307785 251600 307819
rect 251548 307776 251600 307785
rect 270776 307819 270828 307828
rect 270776 307785 270785 307819
rect 270785 307785 270819 307819
rect 270819 307785 270828 307819
rect 270776 307776 270828 307785
rect 272248 307819 272300 307828
rect 272248 307785 272257 307819
rect 272257 307785 272291 307819
rect 272291 307785 272300 307819
rect 272248 307776 272300 307785
rect 330208 307819 330260 307828
rect 330208 307785 330217 307819
rect 330217 307785 330251 307819
rect 330251 307785 330260 307819
rect 330208 307776 330260 307785
rect 393596 307819 393648 307828
rect 393596 307785 393605 307819
rect 393605 307785 393639 307819
rect 393639 307785 393648 307819
rect 393596 307776 393648 307785
rect 460204 307819 460256 307828
rect 460204 307785 460213 307819
rect 460213 307785 460247 307819
rect 460247 307785 460256 307819
rect 460204 307776 460256 307785
rect 288808 307708 288860 307760
rect 310704 307751 310756 307760
rect 310704 307717 310713 307751
rect 310713 307717 310747 307751
rect 310747 307717 310756 307751
rect 310704 307708 310756 307717
rect 337108 307751 337160 307760
rect 337108 307717 337117 307751
rect 337117 307717 337151 307751
rect 337151 307717 337160 307751
rect 337108 307708 337160 307717
rect 286140 306348 286192 306400
rect 286232 306348 286284 306400
rect 288716 306391 288768 306400
rect 288716 306357 288725 306391
rect 288725 306357 288759 306391
rect 288759 306357 288768 306391
rect 288716 306348 288768 306357
rect 317512 306348 317564 306400
rect 317696 306348 317748 306400
rect 463700 306348 463752 306400
rect 463884 306348 463936 306400
rect 580080 306348 580132 306400
rect 580908 306348 580960 306400
rect 266636 305031 266688 305040
rect 266636 304997 266645 305031
rect 266645 304997 266679 305031
rect 266679 304997 266688 305031
rect 266636 304988 266688 304997
rect 291752 304920 291804 304972
rect 291844 304920 291896 304972
rect 294236 304240 294288 304292
rect 294420 304240 294472 304292
rect 295524 304240 295576 304292
rect 295708 304240 295760 304292
rect 323216 304283 323268 304292
rect 323216 304249 323225 304283
rect 323225 304249 323259 304283
rect 323259 304249 323268 304283
rect 323216 304240 323268 304249
rect 291752 303560 291804 303612
rect 259736 302268 259788 302320
rect 357532 302200 357584 302252
rect 357716 302200 357768 302252
rect 389180 302200 389232 302252
rect 389364 302200 389416 302252
rect 431316 302200 431368 302252
rect 431500 302200 431552 302252
rect 296812 301112 296864 301164
rect 296996 301112 297048 301164
rect 265348 300092 265400 300144
rect 262680 299616 262732 299668
rect 331404 299591 331456 299600
rect 331404 299557 331413 299591
rect 331413 299557 331447 299591
rect 331447 299557 331456 299591
rect 331404 299548 331456 299557
rect 266636 299480 266688 299532
rect 266728 299480 266780 299532
rect 299756 299480 299808 299532
rect 299848 299480 299900 299532
rect 302516 299480 302568 299532
rect 302608 299480 302660 299532
rect 306840 299523 306892 299532
rect 306840 299489 306849 299523
rect 306849 299489 306883 299523
rect 306883 299489 306892 299523
rect 306840 299480 306892 299489
rect 323308 299480 323360 299532
rect 341156 299523 341208 299532
rect 341156 299489 341165 299523
rect 341165 299489 341199 299523
rect 341199 299489 341208 299523
rect 341156 299480 341208 299489
rect 367008 299523 367060 299532
rect 367008 299489 367017 299523
rect 367017 299489 367051 299523
rect 367051 299489 367060 299523
rect 367008 299480 367060 299489
rect 235080 299455 235132 299464
rect 235080 299421 235089 299455
rect 235089 299421 235123 299455
rect 235123 299421 235132 299455
rect 235080 299412 235132 299421
rect 236276 299455 236328 299464
rect 236276 299421 236285 299455
rect 236285 299421 236319 299455
rect 236319 299421 236328 299455
rect 236276 299412 236328 299421
rect 270776 299455 270828 299464
rect 270776 299421 270785 299455
rect 270785 299421 270819 299455
rect 270819 299421 270828 299455
rect 270776 299412 270828 299421
rect 272248 299455 272300 299464
rect 272248 299421 272257 299455
rect 272257 299421 272291 299455
rect 272291 299421 272300 299455
rect 272248 299412 272300 299421
rect 273536 299412 273588 299464
rect 281724 299412 281776 299464
rect 281816 299412 281868 299464
rect 284668 299412 284720 299464
rect 284760 299412 284812 299464
rect 324688 299455 324740 299464
rect 324688 299421 324697 299455
rect 324697 299421 324731 299455
rect 324731 299421 324740 299455
rect 324688 299412 324740 299421
rect 325884 299412 325936 299464
rect 372712 299455 372764 299464
rect 372712 299421 372721 299455
rect 372721 299421 372755 299455
rect 372755 299421 372764 299455
rect 372712 299412 372764 299421
rect 469864 299412 469916 299464
rect 580172 299412 580224 299464
rect 325976 299344 326028 299396
rect 273536 299276 273588 299328
rect 286048 298188 286100 298240
rect 286140 298188 286192 298240
rect 247040 298120 247092 298172
rect 247316 298120 247368 298172
rect 288900 298120 288952 298172
rect 310888 298120 310940 298172
rect 337292 298120 337344 298172
rect 251548 298052 251600 298104
rect 266728 298095 266780 298104
rect 266728 298061 266737 298095
rect 266737 298061 266771 298095
rect 266771 298061 266780 298095
rect 266728 298052 266780 298061
rect 281724 298052 281776 298104
rect 281816 298052 281868 298104
rect 284668 298052 284720 298104
rect 284760 298052 284812 298104
rect 286048 298052 286100 298104
rect 286140 298052 286192 298104
rect 301044 298095 301096 298104
rect 301044 298061 301053 298095
rect 301053 298061 301087 298095
rect 301087 298061 301096 298095
rect 301044 298052 301096 298061
rect 393596 298095 393648 298104
rect 393596 298061 393605 298095
rect 393605 298061 393639 298095
rect 393639 298061 393648 298095
rect 393596 298052 393648 298061
rect 460020 298095 460072 298104
rect 460020 298061 460029 298095
rect 460029 298061 460063 298095
rect 460063 298061 460072 298095
rect 460020 298052 460072 298061
rect 288900 297984 288952 298036
rect 580080 296760 580132 296812
rect 581000 296760 581052 296812
rect 259644 296735 259696 296744
rect 259644 296701 259653 296735
rect 259653 296701 259687 296735
rect 259687 296701 259696 296735
rect 259644 296692 259696 296701
rect 262588 296735 262640 296744
rect 262588 296701 262597 296735
rect 262597 296701 262631 296735
rect 262631 296701 262640 296735
rect 262588 296692 262640 296701
rect 267740 296692 267792 296744
rect 268016 296692 268068 296744
rect 580172 296624 580224 296676
rect 581000 296624 581052 296676
rect 267740 296556 267792 296608
rect 291568 296531 291620 296540
rect 291568 296497 291577 296531
rect 291577 296497 291611 296531
rect 291611 296497 291620 296531
rect 291568 296488 291620 296497
rect 290004 294584 290056 294636
rect 290188 294584 290240 294636
rect 265348 293904 265400 293956
rect 265532 293904 265584 293956
rect 310888 293063 310940 293072
rect 310888 293029 310897 293063
rect 310897 293029 310931 293063
rect 310931 293029 310940 293063
rect 310888 293020 310940 293029
rect 299848 292612 299900 292664
rect 306840 292612 306892 292664
rect 295524 292544 295576 292596
rect 239128 292476 239180 292528
rect 291568 292476 291620 292528
rect 295616 292476 295668 292528
rect 299848 292476 299900 292528
rect 301044 292519 301096 292528
rect 301044 292485 301053 292519
rect 301053 292485 301087 292519
rect 301087 292485 301096 292519
rect 301044 292476 301096 292485
rect 306840 292476 306892 292528
rect 239128 292340 239180 292392
rect 337108 290368 337160 290420
rect 337292 290368 337344 290420
rect 235080 289867 235132 289876
rect 235080 289833 235089 289867
rect 235089 289833 235123 289867
rect 235123 289833 235132 289867
rect 235080 289824 235132 289833
rect 236276 289867 236328 289876
rect 236276 289833 236285 289867
rect 236285 289833 236319 289867
rect 236319 289833 236328 289867
rect 236276 289824 236328 289833
rect 247040 289824 247092 289876
rect 247224 289824 247276 289876
rect 270776 289867 270828 289876
rect 270776 289833 270785 289867
rect 270785 289833 270819 289867
rect 270819 289833 270828 289867
rect 270776 289824 270828 289833
rect 324688 289867 324740 289876
rect 324688 289833 324697 289867
rect 324697 289833 324731 289867
rect 324731 289833 324740 289867
rect 324688 289824 324740 289833
rect 372712 289867 372764 289876
rect 372712 289833 372721 289867
rect 372721 289833 372755 289867
rect 372755 289833 372764 289867
rect 372712 289824 372764 289833
rect 375840 289824 375892 289876
rect 375932 289824 375984 289876
rect 377128 289824 377180 289876
rect 377220 289824 377272 289876
rect 290004 289756 290056 289808
rect 290188 289756 290240 289808
rect 341248 289756 341300 289808
rect 367008 289799 367060 289808
rect 367008 289765 367017 289799
rect 367017 289765 367051 289799
rect 367051 289765 367060 289799
rect 367008 289756 367060 289765
rect 389456 289756 389508 289808
rect 272248 289323 272300 289332
rect 272248 289289 272257 289323
rect 272257 289289 272291 289323
rect 272291 289289 272300 289323
rect 272248 289280 272300 289289
rect 244464 288396 244516 288448
rect 244556 288396 244608 288448
rect 251364 288439 251416 288448
rect 251364 288405 251373 288439
rect 251373 288405 251407 288439
rect 251407 288405 251416 288439
rect 251364 288396 251416 288405
rect 266820 288396 266872 288448
rect 330116 288396 330168 288448
rect 330208 288396 330260 288448
rect 331404 288396 331456 288448
rect 331496 288396 331548 288448
rect 460112 288396 460164 288448
rect 272248 288328 272300 288380
rect 272340 288328 272392 288380
rect 337108 288371 337160 288380
rect 337108 288337 337117 288371
rect 337117 288337 337151 288371
rect 337151 288337 337160 288371
rect 337108 288328 337160 288337
rect 267740 287036 267792 287088
rect 323308 287036 323360 287088
rect 323492 287036 323544 287088
rect 580172 287036 580224 287088
rect 580908 287036 580960 287088
rect 325976 286968 326028 287020
rect 326068 286968 326120 287020
rect 288992 284248 289044 284300
rect 270776 282956 270828 283008
rect 295616 282956 295668 283008
rect 460112 282956 460164 283008
rect 357532 282888 357584 282940
rect 357716 282888 357768 282940
rect 431316 282888 431368 282940
rect 431500 282888 431552 282940
rect 270684 282820 270736 282872
rect 295524 282820 295576 282872
rect 310888 282795 310940 282804
rect 310888 282761 310897 282795
rect 310897 282761 310931 282795
rect 310931 282761 310940 282795
rect 310888 282752 310940 282761
rect 460112 282752 460164 282804
rect 266728 280168 266780 280220
rect 266820 280168 266872 280220
rect 294236 280168 294288 280220
rect 294328 280168 294380 280220
rect 327172 280211 327224 280220
rect 327172 280177 327181 280211
rect 327181 280177 327215 280211
rect 327215 280177 327224 280211
rect 327172 280168 327224 280177
rect 341156 280211 341208 280220
rect 341156 280177 341165 280211
rect 341165 280177 341199 280211
rect 341199 280177 341208 280211
rect 341156 280168 341208 280177
rect 367008 280211 367060 280220
rect 367008 280177 367017 280211
rect 367017 280177 367051 280211
rect 367051 280177 367060 280211
rect 367008 280168 367060 280177
rect 389364 280211 389416 280220
rect 389364 280177 389373 280211
rect 389373 280177 389407 280211
rect 389407 280177 389416 280211
rect 389364 280168 389416 280177
rect 393596 280211 393648 280220
rect 393596 280177 393605 280211
rect 393605 280177 393639 280211
rect 393639 280177 393648 280211
rect 393596 280168 393648 280177
rect 3332 280100 3384 280152
rect 15844 280100 15896 280152
rect 235080 280143 235132 280152
rect 235080 280109 235089 280143
rect 235089 280109 235123 280143
rect 235123 280109 235132 280143
rect 235080 280100 235132 280109
rect 236276 280143 236328 280152
rect 236276 280109 236285 280143
rect 236285 280109 236319 280143
rect 236319 280109 236328 280143
rect 236276 280100 236328 280109
rect 250076 280100 250128 280152
rect 250168 280100 250220 280152
rect 270684 280143 270736 280152
rect 270684 280109 270693 280143
rect 270693 280109 270727 280143
rect 270727 280109 270736 280143
rect 270684 280100 270736 280109
rect 273536 280143 273588 280152
rect 273536 280109 273545 280143
rect 273545 280109 273579 280143
rect 273579 280109 273588 280143
rect 273536 280100 273588 280109
rect 281724 280100 281776 280152
rect 281816 280100 281868 280152
rect 284760 280100 284812 280152
rect 284852 280100 284904 280152
rect 372712 280143 372764 280152
rect 372712 280109 372721 280143
rect 372721 280109 372755 280143
rect 372755 280109 372764 280143
rect 372712 280100 372764 280109
rect 375840 280143 375892 280152
rect 375840 280109 375849 280143
rect 375849 280109 375883 280143
rect 375883 280109 375892 280143
rect 375840 280100 375892 280109
rect 377128 280143 377180 280152
rect 377128 280109 377137 280143
rect 377137 280109 377171 280143
rect 377171 280109 377180 280143
rect 377128 280100 377180 280109
rect 460112 280143 460164 280152
rect 460112 280109 460121 280143
rect 460121 280109 460155 280143
rect 460155 280109 460164 280143
rect 460112 280100 460164 280109
rect 329932 278876 329984 278928
rect 330208 278876 330260 278928
rect 327172 278783 327224 278792
rect 327172 278749 327181 278783
rect 327181 278749 327215 278783
rect 327215 278749 327224 278783
rect 327172 278740 327224 278749
rect 331496 278808 331548 278860
rect 337200 278740 337252 278792
rect 310888 278715 310940 278724
rect 310888 278681 310897 278715
rect 310897 278681 310931 278715
rect 310931 278681 310940 278715
rect 310888 278672 310940 278681
rect 331404 278672 331456 278724
rect 393596 278715 393648 278724
rect 393596 278681 393605 278715
rect 393605 278681 393639 278715
rect 393639 278681 393648 278715
rect 393596 278672 393648 278681
rect 296812 277380 296864 277432
rect 296904 277380 296956 277432
rect 331404 277355 331456 277364
rect 331404 277321 331413 277355
rect 331413 277321 331447 277355
rect 331447 277321 331456 277355
rect 331404 277312 331456 277321
rect 580172 277312 580224 277364
rect 580908 277312 580960 277364
rect 294236 275952 294288 276004
rect 294328 275952 294380 276004
rect 297088 275952 297140 276004
rect 270684 275315 270736 275324
rect 270684 275281 270693 275315
rect 270693 275281 270727 275315
rect 270727 275281 270736 275315
rect 270684 275272 270736 275281
rect 463792 275315 463844 275324
rect 463792 275281 463801 275315
rect 463801 275281 463835 275315
rect 463835 275281 463844 275315
rect 463792 275272 463844 275281
rect 288900 274703 288952 274712
rect 288900 274669 288909 274703
rect 288909 274669 288943 274703
rect 288943 274669 288952 274703
rect 288900 274660 288952 274669
rect 291384 274703 291436 274712
rect 291384 274669 291393 274703
rect 291393 274669 291427 274703
rect 291427 274669 291436 274703
rect 291384 274660 291436 274669
rect 250076 273912 250128 273964
rect 250260 273912 250312 273964
rect 323308 273343 323360 273352
rect 323308 273309 323317 273343
rect 323317 273309 323351 273343
rect 323351 273309 323360 273343
rect 323308 273300 323360 273309
rect 301044 273232 301096 273284
rect 239128 273164 239180 273216
rect 337200 273300 337252 273352
rect 301136 273164 301188 273216
rect 337108 273164 337160 273216
rect 460112 273139 460164 273148
rect 460112 273105 460121 273139
rect 460121 273105 460155 273139
rect 460155 273105 460164 273139
rect 460112 273096 460164 273105
rect 239128 273028 239180 273080
rect 299848 270580 299900 270632
rect 235080 270555 235132 270564
rect 235080 270521 235089 270555
rect 235089 270521 235123 270555
rect 235123 270521 235132 270555
rect 235080 270512 235132 270521
rect 236276 270555 236328 270564
rect 236276 270521 236285 270555
rect 236285 270521 236319 270555
rect 236319 270521 236328 270555
rect 236276 270512 236328 270521
rect 247040 270512 247092 270564
rect 247224 270512 247276 270564
rect 251180 270512 251232 270564
rect 251456 270512 251508 270564
rect 273536 270555 273588 270564
rect 273536 270521 273545 270555
rect 273545 270521 273579 270555
rect 273579 270521 273588 270555
rect 273536 270512 273588 270521
rect 299756 270512 299808 270564
rect 302516 270512 302568 270564
rect 302700 270512 302752 270564
rect 327172 270512 327224 270564
rect 327264 270512 327316 270564
rect 372712 270555 372764 270564
rect 372712 270521 372721 270555
rect 372721 270521 372755 270555
rect 372755 270521 372764 270555
rect 372712 270512 372764 270521
rect 375840 270555 375892 270564
rect 375840 270521 375849 270555
rect 375849 270521 375883 270555
rect 375883 270521 375892 270555
rect 375840 270512 375892 270521
rect 377128 270555 377180 270564
rect 377128 270521 377137 270555
rect 377137 270521 377171 270555
rect 377171 270521 377180 270555
rect 377128 270512 377180 270521
rect 463884 270512 463936 270564
rect 286048 270444 286100 270496
rect 286140 270444 286192 270496
rect 341248 270444 341300 270496
rect 367008 270487 367060 270496
rect 367008 270453 367017 270487
rect 367017 270453 367051 270487
rect 367051 270453 367060 270487
rect 367008 270444 367060 270453
rect 389456 270444 389508 270496
rect 460112 270444 460164 270496
rect 245936 269084 245988 269136
rect 246120 269084 246172 269136
rect 259644 269084 259696 269136
rect 259736 269084 259788 269136
rect 265256 269084 265308 269136
rect 290096 269084 290148 269136
rect 290188 269084 290240 269136
rect 295524 269084 295576 269136
rect 295800 269084 295852 269136
rect 265164 269016 265216 269068
rect 324504 267792 324556 267844
rect 324688 267792 324740 267844
rect 323308 267767 323360 267776
rect 323308 267733 323317 267767
rect 323317 267733 323351 267767
rect 323351 267733 323360 267767
rect 323308 267724 323360 267733
rect 325976 267724 326028 267776
rect 326068 267724 326120 267776
rect 329932 267724 329984 267776
rect 330116 267724 330168 267776
rect 331404 267767 331456 267776
rect 331404 267733 331413 267767
rect 331413 267733 331447 267767
rect 331447 267733 331456 267767
rect 331404 267724 331456 267733
rect 296996 266407 297048 266416
rect 296996 266373 297005 266407
rect 297005 266373 297039 266407
rect 297039 266373 297048 266407
rect 296996 266364 297048 266373
rect 294328 266296 294380 266348
rect 294420 266296 294472 266348
rect 250168 264299 250220 264308
rect 250168 264265 250177 264299
rect 250177 264265 250211 264299
rect 250211 264265 250220 264299
rect 250168 264256 250220 264265
rect 266728 263619 266780 263628
rect 266728 263585 266737 263619
rect 266737 263585 266771 263619
rect 266771 263585 266780 263619
rect 266728 263576 266780 263585
rect 270684 263576 270736 263628
rect 357532 263576 357584 263628
rect 357716 263576 357768 263628
rect 431316 263576 431368 263628
rect 431500 263576 431552 263628
rect 270684 263440 270736 263492
rect 310888 263483 310940 263492
rect 310888 263449 310897 263483
rect 310897 263449 310931 263483
rect 310931 263449 310940 263483
rect 310888 263440 310940 263449
rect 296812 262896 296864 262948
rect 296996 262896 297048 262948
rect 247132 260856 247184 260908
rect 235080 260831 235132 260840
rect 235080 260797 235089 260831
rect 235089 260797 235123 260831
rect 235123 260797 235132 260831
rect 235080 260788 235132 260797
rect 236276 260831 236328 260840
rect 236276 260797 236285 260831
rect 236285 260797 236319 260831
rect 236319 260797 236328 260831
rect 236276 260788 236328 260797
rect 270684 260831 270736 260840
rect 270684 260797 270693 260831
rect 270693 260797 270727 260831
rect 270727 260797 270736 260831
rect 270684 260788 270736 260797
rect 272340 260924 272392 260976
rect 281816 260899 281868 260908
rect 281816 260865 281825 260899
rect 281825 260865 281859 260899
rect 281859 260865 281868 260899
rect 281816 260856 281868 260865
rect 324596 260899 324648 260908
rect 324596 260865 324605 260899
rect 324605 260865 324639 260899
rect 324639 260865 324648 260899
rect 324596 260856 324648 260865
rect 273536 260831 273588 260840
rect 273536 260797 273545 260831
rect 273545 260797 273579 260831
rect 273579 260797 273588 260831
rect 273536 260788 273588 260797
rect 327264 260924 327316 260976
rect 460020 260967 460072 260976
rect 460020 260933 460029 260967
rect 460029 260933 460063 260967
rect 460063 260933 460072 260967
rect 460020 260924 460072 260933
rect 341156 260899 341208 260908
rect 341156 260865 341165 260899
rect 341165 260865 341199 260899
rect 341199 260865 341208 260899
rect 341156 260856 341208 260865
rect 367008 260899 367060 260908
rect 367008 260865 367017 260899
rect 367017 260865 367051 260899
rect 367051 260865 367060 260899
rect 367008 260856 367060 260865
rect 389364 260899 389416 260908
rect 389364 260865 389373 260899
rect 389373 260865 389407 260899
rect 389407 260865 389416 260899
rect 389364 260856 389416 260865
rect 393596 260899 393648 260908
rect 393596 260865 393605 260899
rect 393605 260865 393639 260899
rect 393639 260865 393648 260899
rect 393596 260856 393648 260865
rect 372712 260831 372764 260840
rect 372712 260797 372721 260831
rect 372721 260797 372755 260831
rect 372755 260797 372764 260831
rect 372712 260788 372764 260797
rect 375840 260831 375892 260840
rect 375840 260797 375849 260831
rect 375849 260797 375883 260831
rect 375883 260797 375892 260831
rect 375840 260788 375892 260797
rect 377128 260831 377180 260840
rect 377128 260797 377137 260831
rect 377137 260797 377171 260831
rect 377171 260797 377180 260831
rect 377128 260788 377180 260797
rect 460020 260788 460072 260840
rect 460204 260788 460256 260840
rect 463792 260788 463844 260840
rect 272156 260720 272208 260772
rect 327172 260720 327224 260772
rect 247224 259607 247276 259616
rect 247224 259573 247233 259607
rect 247233 259573 247267 259607
rect 247267 259573 247276 259607
rect 247224 259564 247276 259573
rect 244372 259428 244424 259480
rect 244464 259428 244516 259480
rect 250168 259471 250220 259480
rect 250168 259437 250177 259471
rect 250177 259437 250211 259471
rect 250211 259437 250220 259471
rect 250168 259428 250220 259437
rect 266728 259471 266780 259480
rect 266728 259437 266737 259471
rect 266737 259437 266771 259471
rect 266771 259437 266780 259471
rect 266728 259428 266780 259437
rect 281816 259471 281868 259480
rect 281816 259437 281825 259471
rect 281825 259437 281859 259471
rect 281859 259437 281868 259471
rect 281816 259428 281868 259437
rect 284760 259428 284812 259480
rect 284852 259428 284904 259480
rect 337108 259428 337160 259480
rect 337292 259428 337344 259480
rect 331404 259403 331456 259412
rect 331404 259369 331413 259403
rect 331413 259369 331447 259403
rect 331447 259369 331456 259403
rect 331404 259360 331456 259369
rect 288900 259088 288952 259140
rect 324596 258111 324648 258120
rect 324596 258077 324605 258111
rect 324605 258077 324639 258111
rect 324639 258077 324648 258111
rect 324596 258068 324648 258077
rect 247224 258043 247276 258052
rect 247224 258009 247233 258043
rect 247233 258009 247267 258043
rect 247267 258009 247276 258043
rect 247224 258000 247276 258009
rect 262312 258000 262364 258052
rect 262588 258000 262640 258052
rect 291476 258000 291528 258052
rect 291568 258000 291620 258052
rect 295524 258000 295576 258052
rect 295708 258000 295760 258052
rect 330116 258000 330168 258052
rect 330300 258000 330352 258052
rect 296996 257932 297048 257984
rect 310888 256071 310940 256080
rect 310888 256037 310897 256071
rect 310897 256037 310931 256071
rect 310931 256037 310940 256071
rect 310888 256028 310940 256037
rect 270684 256003 270736 256012
rect 270684 255969 270693 256003
rect 270693 255969 270727 256003
rect 270727 255969 270736 256003
rect 270684 255960 270736 255969
rect 286140 255892 286192 255944
rect 259736 254600 259788 254652
rect 323308 253920 323360 253972
rect 337108 253920 337160 253972
rect 239128 253852 239180 253904
rect 337292 253784 337344 253836
rect 239128 253716 239180 253768
rect 294420 251812 294472 251864
rect 367008 251404 367060 251456
rect 310704 251268 310756 251320
rect 366824 251268 366876 251320
rect 235080 251243 235132 251252
rect 235080 251209 235089 251243
rect 235089 251209 235123 251243
rect 235123 251209 235132 251243
rect 235080 251200 235132 251209
rect 236276 251243 236328 251252
rect 236276 251209 236285 251243
rect 236285 251209 236319 251243
rect 236319 251209 236328 251243
rect 236276 251200 236328 251209
rect 251180 251200 251232 251252
rect 251456 251200 251508 251252
rect 273536 251243 273588 251252
rect 273536 251209 273545 251243
rect 273545 251209 273579 251243
rect 273579 251209 273588 251243
rect 273536 251200 273588 251209
rect 290004 251200 290056 251252
rect 290096 251200 290148 251252
rect 366916 251200 366968 251252
rect 367008 251200 367060 251252
rect 372712 251243 372764 251252
rect 372712 251209 372721 251243
rect 372721 251209 372755 251243
rect 372755 251209 372764 251243
rect 372712 251200 372764 251209
rect 375840 251243 375892 251252
rect 375840 251209 375849 251243
rect 375849 251209 375883 251243
rect 375883 251209 375892 251243
rect 375840 251200 375892 251209
rect 377128 251243 377180 251252
rect 377128 251209 377137 251243
rect 377137 251209 377171 251243
rect 377171 251209 377180 251243
rect 377128 251200 377180 251209
rect 389180 251200 389232 251252
rect 389364 251200 389416 251252
rect 463700 251243 463752 251252
rect 463700 251209 463709 251243
rect 463709 251209 463743 251243
rect 463743 251209 463752 251243
rect 463700 251200 463752 251209
rect 250168 251175 250220 251184
rect 250168 251141 250177 251175
rect 250177 251141 250211 251175
rect 250211 251141 250220 251175
rect 250168 251132 250220 251141
rect 281816 251175 281868 251184
rect 281816 251141 281825 251175
rect 281825 251141 281859 251175
rect 281859 251141 281868 251175
rect 281816 251132 281868 251141
rect 284668 251132 284720 251184
rect 284760 251132 284812 251184
rect 310704 251175 310756 251184
rect 310704 251141 310713 251175
rect 310713 251141 310747 251175
rect 310747 251141 310756 251175
rect 310704 251132 310756 251141
rect 460112 251132 460164 251184
rect 367008 251107 367060 251116
rect 367008 251073 367017 251107
rect 367017 251073 367051 251107
rect 367051 251073 367060 251107
rect 367008 251064 367060 251073
rect 301136 249840 301188 249892
rect 330024 249840 330076 249892
rect 245844 249772 245896 249824
rect 246028 249772 246080 249824
rect 299756 249772 299808 249824
rect 299940 249772 299992 249824
rect 302516 249772 302568 249824
rect 302608 249772 302660 249824
rect 306748 249772 306800 249824
rect 306932 249772 306984 249824
rect 323400 249815 323452 249824
rect 323400 249781 323409 249815
rect 323409 249781 323443 249815
rect 323443 249781 323452 249815
rect 323400 249772 323452 249781
rect 393596 249772 393648 249824
rect 393780 249772 393832 249824
rect 247224 249747 247276 249756
rect 247224 249713 247233 249747
rect 247233 249713 247267 249747
rect 247267 249713 247276 249747
rect 247224 249704 247276 249713
rect 330024 249704 330076 249756
rect 296812 249475 296864 249484
rect 296812 249441 296821 249475
rect 296821 249441 296855 249475
rect 296855 249441 296864 249475
rect 296812 249432 296864 249441
rect 301044 248455 301096 248464
rect 301044 248421 301053 248455
rect 301053 248421 301087 248455
rect 301087 248421 301096 248455
rect 301044 248412 301096 248421
rect 284668 248387 284720 248396
rect 284668 248353 284677 248387
rect 284677 248353 284711 248387
rect 284711 248353 284720 248387
rect 284668 248344 284720 248353
rect 306748 248387 306800 248396
rect 306748 248353 306757 248387
rect 306757 248353 306791 248387
rect 306791 248353 306800 248387
rect 306748 248344 306800 248353
rect 286048 247095 286100 247104
rect 286048 247061 286057 247095
rect 286057 247061 286091 247095
rect 286091 247061 286100 247095
rect 286048 247052 286100 247061
rect 329932 244944 329984 244996
rect 330208 244944 330260 244996
rect 341248 244332 341300 244384
rect 357532 244264 357584 244316
rect 357716 244264 357768 244316
rect 431316 244264 431368 244316
rect 431500 244264 431552 244316
rect 341156 244196 341208 244248
rect 259644 241587 259696 241596
rect 259644 241553 259653 241587
rect 259653 241553 259687 241587
rect 259687 241553 259696 241587
rect 259644 241544 259696 241553
rect 250168 241519 250220 241528
rect 250168 241485 250177 241519
rect 250177 241485 250211 241519
rect 250211 241485 250220 241519
rect 250168 241476 250220 241485
rect 266636 241476 266688 241528
rect 266728 241476 266780 241528
rect 281816 241519 281868 241528
rect 281816 241485 281825 241519
rect 281825 241485 281859 241519
rect 281859 241485 281868 241519
rect 281816 241476 281868 241485
rect 288808 241519 288860 241528
rect 288808 241485 288817 241519
rect 288817 241485 288851 241519
rect 288851 241485 288860 241519
rect 288808 241476 288860 241485
rect 290004 241476 290056 241528
rect 290188 241476 290240 241528
rect 291476 241476 291528 241528
rect 291660 241476 291712 241528
rect 310888 241476 310940 241528
rect 367008 241519 367060 241528
rect 367008 241485 367017 241519
rect 367017 241485 367051 241519
rect 367051 241485 367060 241519
rect 367008 241476 367060 241485
rect 460020 241519 460072 241528
rect 460020 241485 460029 241519
rect 460029 241485 460063 241519
rect 460063 241485 460072 241519
rect 460020 241476 460072 241485
rect 270684 241408 270736 241460
rect 270868 241408 270920 241460
rect 272156 241408 272208 241460
rect 272340 241408 272392 241460
rect 299480 241451 299532 241460
rect 299480 241417 299489 241451
rect 299489 241417 299523 241451
rect 299523 241417 299532 241451
rect 375840 241451 375892 241460
rect 299480 241408 299532 241417
rect 375840 241417 375849 241451
rect 375849 241417 375883 241451
rect 375883 241417 375892 241451
rect 375840 241408 375892 241417
rect 463792 241451 463844 241460
rect 463792 241417 463801 241451
rect 463801 241417 463835 241451
rect 463835 241417 463844 241451
rect 463792 241408 463844 241417
rect 244372 240116 244424 240168
rect 244556 240116 244608 240168
rect 245936 240116 245988 240168
rect 246120 240116 246172 240168
rect 251180 240116 251232 240168
rect 251364 240116 251416 240168
rect 262496 240116 262548 240168
rect 262588 240116 262640 240168
rect 267740 240116 267792 240168
rect 267832 240116 267884 240168
rect 299756 240116 299808 240168
rect 299940 240116 299992 240168
rect 301044 240116 301096 240168
rect 301136 240116 301188 240168
rect 302516 240116 302568 240168
rect 302700 240116 302752 240168
rect 306840 240048 306892 240100
rect 284760 238756 284812 238808
rect 294420 238756 294472 238808
rect 285956 238688 286008 238740
rect 393320 238688 393372 238740
rect 393504 238688 393556 238740
rect 286140 238552 286192 238604
rect 3332 237328 3384 237380
rect 17224 237328 17276 237380
rect 331404 236691 331456 236700
rect 331404 236657 331413 236691
rect 331413 236657 331447 236691
rect 331447 236657 331456 236691
rect 331404 236648 331456 236657
rect 267740 234676 267792 234728
rect 281816 234676 281868 234728
rect 244464 234608 244516 234660
rect 250076 234608 250128 234660
rect 310888 234676 310940 234728
rect 463976 234608 464028 234660
rect 239128 234540 239180 234592
rect 244372 234540 244424 234592
rect 267740 234540 267792 234592
rect 281816 234540 281868 234592
rect 310796 234540 310848 234592
rect 239128 234404 239180 234456
rect 323400 233860 323452 233912
rect 323584 233860 323636 233912
rect 234896 231820 234948 231872
rect 235080 231820 235132 231872
rect 236276 231820 236328 231872
rect 236460 231820 236512 231872
rect 273536 231820 273588 231872
rect 273720 231820 273772 231872
rect 299480 231863 299532 231872
rect 299480 231829 299489 231863
rect 299489 231829 299523 231863
rect 299523 231829 299532 231863
rect 299480 231820 299532 231829
rect 301136 231820 301188 231872
rect 302700 231888 302752 231940
rect 306932 231888 306984 231940
rect 324688 231820 324740 231872
rect 324780 231820 324832 231872
rect 325976 231820 326028 231872
rect 326068 231820 326120 231872
rect 327264 231820 327316 231872
rect 327356 231820 327408 231872
rect 372528 231820 372580 231872
rect 372712 231820 372764 231872
rect 375840 231863 375892 231872
rect 375840 231829 375849 231863
rect 375849 231829 375883 231863
rect 375883 231829 375892 231863
rect 375840 231820 375892 231829
rect 376944 231820 376996 231872
rect 377128 231820 377180 231872
rect 301228 231752 301280 231804
rect 302608 231752 302660 231804
rect 306840 231752 306892 231804
rect 310796 231795 310848 231804
rect 310796 231761 310805 231795
rect 310805 231761 310839 231795
rect 310839 231761 310848 231795
rect 310796 231752 310848 231761
rect 367008 231795 367060 231804
rect 367008 231761 367017 231795
rect 367017 231761 367051 231795
rect 367051 231761 367060 231795
rect 367008 231752 367060 231761
rect 250168 230503 250220 230512
rect 250168 230469 250177 230503
rect 250177 230469 250211 230503
rect 250211 230469 250220 230503
rect 250168 230460 250220 230469
rect 251088 230460 251140 230512
rect 251364 230460 251416 230512
rect 259552 230460 259604 230512
rect 259644 230460 259696 230512
rect 270684 230460 270736 230512
rect 270776 230460 270828 230512
rect 288716 230460 288768 230512
rect 288808 230460 288860 230512
rect 330208 230460 330260 230512
rect 330392 230460 330444 230512
rect 341248 230460 341300 230512
rect 341432 230460 341484 230512
rect 337292 225335 337344 225344
rect 337292 225301 337301 225335
rect 337301 225301 337335 225335
rect 337335 225301 337344 225335
rect 337292 225292 337344 225301
rect 270684 224952 270736 225004
rect 288716 224952 288768 225004
rect 270684 224816 270736 224868
rect 341248 225020 341300 225072
rect 357532 224952 357584 225004
rect 357716 224952 357768 225004
rect 431316 224952 431368 225004
rect 431500 224952 431552 225004
rect 460112 225020 460164 225072
rect 341156 224884 341208 224936
rect 460020 224884 460072 224936
rect 288808 224816 288860 224868
rect 393320 224204 393372 224256
rect 393504 224204 393556 224256
rect 2780 223048 2832 223100
rect 5172 223048 5224 223100
rect 325976 222232 326028 222284
rect 327264 222232 327316 222284
rect 265164 222164 265216 222216
rect 265348 222164 265400 222216
rect 294328 222164 294380 222216
rect 294420 222164 294472 222216
rect 295524 222164 295576 222216
rect 295616 222164 295668 222216
rect 296812 222164 296864 222216
rect 296904 222164 296956 222216
rect 301044 222164 301096 222216
rect 301228 222164 301280 222216
rect 310888 222164 310940 222216
rect 325884 222164 325936 222216
rect 327172 222164 327224 222216
rect 330116 222164 330168 222216
rect 330208 222164 330260 222216
rect 331404 222207 331456 222216
rect 331404 222173 331413 222207
rect 331413 222173 331447 222207
rect 331447 222173 331456 222207
rect 331404 222164 331456 222173
rect 337292 222207 337344 222216
rect 337292 222173 337301 222207
rect 337301 222173 337335 222207
rect 337335 222173 337344 222207
rect 337292 222164 337344 222173
rect 367008 222207 367060 222216
rect 367008 222173 367017 222207
rect 367017 222173 367051 222207
rect 367051 222173 367060 222207
rect 367008 222164 367060 222173
rect 389272 222164 389324 222216
rect 389548 222164 389600 222216
rect 463792 222164 463844 222216
rect 464068 222164 464120 222216
rect 270684 222139 270736 222148
rect 270684 222105 270693 222139
rect 270693 222105 270727 222139
rect 270727 222105 270736 222139
rect 270684 222096 270736 222105
rect 272156 222096 272208 222148
rect 272248 222096 272300 222148
rect 375840 222139 375892 222148
rect 375840 222105 375849 222139
rect 375849 222105 375883 222139
rect 375883 222105 375892 222139
rect 375840 222096 375892 222105
rect 290372 220872 290424 220924
rect 291844 220940 291896 220992
rect 245844 220804 245896 220856
rect 246028 220804 246080 220856
rect 251548 220804 251600 220856
rect 251640 220804 251692 220856
rect 290188 220804 290240 220856
rect 291660 220804 291712 220856
rect 331404 220847 331456 220856
rect 331404 220813 331413 220847
rect 331413 220813 331447 220847
rect 331447 220813 331456 220847
rect 331404 220804 331456 220813
rect 244372 220779 244424 220788
rect 244372 220745 244381 220779
rect 244381 220745 244415 220779
rect 244415 220745 244424 220779
rect 244372 220736 244424 220745
rect 341156 220779 341208 220788
rect 341156 220745 341165 220779
rect 341165 220745 341199 220779
rect 341199 220745 341208 220779
rect 341156 220736 341208 220745
rect 290188 219419 290240 219428
rect 290188 219385 290197 219419
rect 290197 219385 290231 219419
rect 290231 219385 290240 219419
rect 290188 219376 290240 219385
rect 291660 219419 291712 219428
rect 291660 219385 291669 219419
rect 291669 219385 291703 219419
rect 291703 219385 291712 219419
rect 291660 219376 291712 219385
rect 317512 219376 317564 219428
rect 317696 219376 317748 219428
rect 301044 215296 301096 215348
rect 239128 215228 239180 215280
rect 310888 215364 310940 215416
rect 389548 215364 389600 215416
rect 464068 215364 464120 215416
rect 310796 215228 310848 215280
rect 341156 215271 341208 215280
rect 341156 215237 341165 215271
rect 341165 215237 341199 215271
rect 341199 215237 341208 215271
rect 341156 215228 341208 215237
rect 389456 215228 389508 215280
rect 459836 215228 459888 215280
rect 460020 215228 460072 215280
rect 463976 215228 464028 215280
rect 301136 215160 301188 215212
rect 239128 215092 239180 215144
rect 299756 213664 299808 213716
rect 299940 213664 299992 213716
rect 306748 213664 306800 213716
rect 306932 213664 306984 213716
rect 330208 212576 330260 212628
rect 234896 212508 234948 212560
rect 235080 212508 235132 212560
rect 236276 212508 236328 212560
rect 236460 212508 236512 212560
rect 245844 212508 245896 212560
rect 245936 212508 245988 212560
rect 250076 212508 250128 212560
rect 250260 212508 250312 212560
rect 270776 212508 270828 212560
rect 273536 212508 273588 212560
rect 273720 212508 273772 212560
rect 281724 212508 281776 212560
rect 281908 212508 281960 212560
rect 284668 212508 284720 212560
rect 284852 212508 284904 212560
rect 324688 212508 324740 212560
rect 324780 212508 324832 212560
rect 325884 212508 325936 212560
rect 325976 212508 326028 212560
rect 327172 212508 327224 212560
rect 327264 212508 327316 212560
rect 372528 212508 372580 212560
rect 372712 212508 372764 212560
rect 375840 212551 375892 212560
rect 375840 212517 375849 212551
rect 375849 212517 375883 212551
rect 375883 212517 375892 212551
rect 375840 212508 375892 212517
rect 376944 212508 376996 212560
rect 377128 212508 377180 212560
rect 244464 212440 244516 212492
rect 286048 212483 286100 212492
rect 286048 212449 286057 212483
rect 286057 212449 286091 212483
rect 286091 212449 286100 212483
rect 286048 212440 286100 212449
rect 310796 212483 310848 212492
rect 310796 212449 310805 212483
rect 310805 212449 310839 212483
rect 310839 212449 310848 212483
rect 310796 212440 310848 212449
rect 330208 212440 330260 212492
rect 367008 212483 367060 212492
rect 367008 212449 367017 212483
rect 367017 212449 367051 212483
rect 367051 212449 367060 212483
rect 367008 212440 367060 212449
rect 262496 212100 262548 212152
rect 262680 212100 262732 212152
rect 246948 211080 247000 211132
rect 247224 211080 247276 211132
rect 249984 211080 250036 211132
rect 250076 211080 250128 211132
rect 290188 211123 290240 211132
rect 290188 211089 290197 211123
rect 290197 211089 290231 211123
rect 290231 211089 290240 211123
rect 290188 211080 290240 211089
rect 330300 211080 330352 211132
rect 317512 209788 317564 209840
rect 317696 209788 317748 209840
rect 281724 205640 281776 205692
rect 284668 205640 284720 205692
rect 288716 205640 288768 205692
rect 357532 205640 357584 205692
rect 357716 205640 357768 205692
rect 431316 205640 431368 205692
rect 431500 205640 431552 205692
rect 281816 205504 281868 205556
rect 460112 205708 460164 205760
rect 288808 205572 288860 205624
rect 460020 205572 460072 205624
rect 284760 205504 284812 205556
rect 393504 204935 393556 204944
rect 393504 204901 393513 204935
rect 393513 204901 393547 204935
rect 393547 204901 393556 204935
rect 393504 204892 393556 204901
rect 291660 204323 291712 204332
rect 291660 204289 291669 204323
rect 291669 204289 291703 204323
rect 291703 204289 291712 204323
rect 291660 204280 291712 204289
rect 331404 202988 331456 203040
rect 325976 202920 326028 202972
rect 327264 202920 327316 202972
rect 244372 202852 244424 202904
rect 244556 202852 244608 202904
rect 245844 202852 245896 202904
rect 245936 202852 245988 202904
rect 262496 202852 262548 202904
rect 262588 202852 262640 202904
rect 270500 202852 270552 202904
rect 270684 202852 270736 202904
rect 286140 202852 286192 202904
rect 294236 202852 294288 202904
rect 294328 202852 294380 202904
rect 295524 202852 295576 202904
rect 295616 202852 295668 202904
rect 296812 202852 296864 202904
rect 296904 202852 296956 202904
rect 299756 202852 299808 202904
rect 299848 202852 299900 202904
rect 301044 202852 301096 202904
rect 301136 202852 301188 202904
rect 302516 202852 302568 202904
rect 302608 202852 302660 202904
rect 306748 202852 306800 202904
rect 306840 202852 306892 202904
rect 310888 202852 310940 202904
rect 325884 202852 325936 202904
rect 327172 202852 327224 202904
rect 331404 202852 331456 202904
rect 337200 202852 337252 202904
rect 337292 202852 337344 202904
rect 341156 202852 341208 202904
rect 341248 202852 341300 202904
rect 367008 202895 367060 202904
rect 367008 202861 367017 202895
rect 367017 202861 367051 202895
rect 367051 202861 367060 202895
rect 367008 202852 367060 202861
rect 389272 202852 389324 202904
rect 389548 202852 389600 202904
rect 463792 202852 463844 202904
rect 464068 202852 464120 202904
rect 330116 202827 330168 202836
rect 330116 202793 330125 202827
rect 330125 202793 330159 202827
rect 330159 202793 330168 202827
rect 330116 202784 330168 202793
rect 375840 202827 375892 202836
rect 375840 202793 375849 202827
rect 375849 202793 375883 202827
rect 375883 202793 375892 202827
rect 375840 202784 375892 202793
rect 250076 201424 250128 201476
rect 250168 201424 250220 201476
rect 306840 201424 306892 201476
rect 306932 201424 306984 201476
rect 324596 201467 324648 201476
rect 324596 201433 324605 201467
rect 324605 201433 324639 201467
rect 324639 201433 324648 201467
rect 324596 201424 324648 201433
rect 327172 201467 327224 201476
rect 327172 201433 327181 201467
rect 327181 201433 327215 201467
rect 327215 201433 327224 201467
rect 327172 201424 327224 201433
rect 330116 201424 330168 201476
rect 330300 201424 330352 201476
rect 250076 200064 250128 200116
rect 250260 200064 250312 200116
rect 290188 200064 290240 200116
rect 317512 200064 317564 200116
rect 317696 200064 317748 200116
rect 330300 200064 330352 200116
rect 330484 200064 330536 200116
rect 331404 200107 331456 200116
rect 331404 200073 331413 200107
rect 331413 200073 331447 200107
rect 331447 200073 331456 200107
rect 331404 200064 331456 200073
rect 266728 198092 266780 198144
rect 266728 197956 266780 198008
rect 232228 195984 232280 196036
rect 299848 196052 299900 196104
rect 301044 195984 301096 196036
rect 232320 195916 232372 195968
rect 235080 195916 235132 195968
rect 299756 195916 299808 195968
rect 302608 196052 302660 196104
rect 310888 196052 310940 196104
rect 337200 196052 337252 196104
rect 389548 196052 389600 196104
rect 460020 195984 460072 196036
rect 302516 195916 302568 195968
rect 310796 195916 310848 195968
rect 337108 195916 337160 195968
rect 389456 195916 389508 195968
rect 301136 195848 301188 195900
rect 464068 196052 464120 196104
rect 463976 195916 464028 195968
rect 460112 195848 460164 195900
rect 235080 195780 235132 195832
rect 230848 193196 230900 193248
rect 231032 193196 231084 193248
rect 236276 193196 236328 193248
rect 236460 193196 236512 193248
rect 244372 193196 244424 193248
rect 244464 193196 244516 193248
rect 247132 193196 247184 193248
rect 247224 193196 247276 193248
rect 259736 193196 259788 193248
rect 259920 193196 259972 193248
rect 265256 193196 265308 193248
rect 265348 193196 265400 193248
rect 267832 193196 267884 193248
rect 267924 193196 267976 193248
rect 270500 193196 270552 193248
rect 270776 193196 270828 193248
rect 273536 193196 273588 193248
rect 273720 193196 273772 193248
rect 281724 193196 281776 193248
rect 281908 193196 281960 193248
rect 284668 193196 284720 193248
rect 284852 193196 284904 193248
rect 288716 193196 288768 193248
rect 288900 193196 288952 193248
rect 341248 193196 341300 193248
rect 341432 193196 341484 193248
rect 372528 193196 372580 193248
rect 372712 193196 372764 193248
rect 375840 193239 375892 193248
rect 375840 193205 375849 193239
rect 375849 193205 375883 193239
rect 375883 193205 375892 193239
rect 375840 193196 375892 193205
rect 376944 193196 376996 193248
rect 377128 193196 377180 193248
rect 324688 193128 324740 193180
rect 327264 193128 327316 193180
rect 367008 193171 367060 193180
rect 367008 193137 367017 193171
rect 367017 193137 367051 193171
rect 367051 193137 367060 193171
rect 367008 193128 367060 193137
rect 393504 193103 393556 193112
rect 393504 193069 393513 193103
rect 393513 193069 393547 193103
rect 393547 193069 393556 193103
rect 393504 193060 393556 193069
rect 245844 191879 245896 191888
rect 245844 191845 245853 191879
rect 245853 191845 245887 191879
rect 245887 191845 245896 191879
rect 245844 191836 245896 191845
rect 285956 191768 286008 191820
rect 286048 191768 286100 191820
rect 331588 191768 331640 191820
rect 337108 191811 337160 191820
rect 337108 191777 337117 191811
rect 337117 191777 337151 191811
rect 337151 191777 337160 191811
rect 337108 191768 337160 191777
rect 393504 191811 393556 191820
rect 393504 191777 393513 191811
rect 393513 191777 393547 191811
rect 393547 191777 393556 191811
rect 393504 191768 393556 191777
rect 290004 190519 290056 190528
rect 290004 190485 290013 190519
rect 290013 190485 290047 190519
rect 290047 190485 290056 190519
rect 290004 190476 290056 190485
rect 317512 190476 317564 190528
rect 317696 190476 317748 190528
rect 267740 190408 267792 190460
rect 267832 190408 267884 190460
rect 331404 190408 331456 190460
rect 331680 190408 331732 190460
rect 245384 189048 245436 189100
rect 290004 188300 290056 188352
rect 290004 188164 290056 188216
rect 339776 186940 339828 186992
rect 339960 186940 340012 186992
rect 251364 186328 251416 186380
rect 266636 186328 266688 186380
rect 251364 186192 251416 186244
rect 295616 186328 295668 186380
rect 296904 186396 296956 186448
rect 357532 186328 357584 186380
rect 357716 186328 357768 186380
rect 431316 186328 431368 186380
rect 431500 186328 431552 186380
rect 460020 186328 460072 186380
rect 295524 186260 295576 186312
rect 296812 186260 296864 186312
rect 337108 186303 337160 186312
rect 337108 186269 337117 186303
rect 337117 186269 337151 186303
rect 337151 186269 337160 186303
rect 337108 186260 337160 186269
rect 460112 186260 460164 186312
rect 266728 186192 266780 186244
rect 264980 183540 265032 183592
rect 265164 183540 265216 183592
rect 270500 183540 270552 183592
rect 270684 183540 270736 183592
rect 291568 183540 291620 183592
rect 291660 183540 291712 183592
rect 299756 183540 299808 183592
rect 299848 183540 299900 183592
rect 301044 183540 301096 183592
rect 301136 183540 301188 183592
rect 302516 183540 302568 183592
rect 302608 183540 302660 183592
rect 306840 183540 306892 183592
rect 306932 183540 306984 183592
rect 310888 183540 310940 183592
rect 311072 183540 311124 183592
rect 324596 183540 324648 183592
rect 324780 183540 324832 183592
rect 327172 183540 327224 183592
rect 327356 183540 327408 183592
rect 367008 183583 367060 183592
rect 367008 183549 367017 183583
rect 367017 183549 367051 183583
rect 367051 183549 367060 183583
rect 367008 183540 367060 183549
rect 389272 183540 389324 183592
rect 389548 183540 389600 183592
rect 463792 183540 463844 183592
rect 464068 183540 464120 183592
rect 251364 183472 251416 183524
rect 251548 183472 251600 183524
rect 393504 183515 393556 183524
rect 393504 183481 393513 183515
rect 393513 183481 393547 183515
rect 393547 183481 393556 183515
rect 393504 183472 393556 183481
rect 460112 183515 460164 183524
rect 460112 183481 460121 183515
rect 460121 183481 460155 183515
rect 460155 183481 460164 183515
rect 460112 183472 460164 183481
rect 272064 182112 272116 182164
rect 272340 182112 272392 182164
rect 273720 182112 273772 182164
rect 290004 182155 290056 182164
rect 290004 182121 290013 182155
rect 290013 182121 290047 182155
rect 290047 182121 290056 182155
rect 290004 182112 290056 182121
rect 291660 182155 291712 182164
rect 291660 182121 291669 182155
rect 291669 182121 291703 182155
rect 291703 182121 291712 182155
rect 291660 182112 291712 182121
rect 341156 182112 341208 182164
rect 341248 182112 341300 182164
rect 393320 182112 393372 182164
rect 393504 182112 393556 182164
rect 329932 182044 329984 182096
rect 330116 182044 330168 182096
rect 245752 180931 245804 180940
rect 245752 180897 245761 180931
rect 245761 180897 245795 180931
rect 245795 180897 245804 180931
rect 245752 180888 245804 180897
rect 245660 180820 245712 180872
rect 267832 180752 267884 180804
rect 267924 180752 267976 180804
rect 301044 180795 301096 180804
rect 301044 180761 301053 180795
rect 301053 180761 301087 180795
rect 301087 180761 301096 180795
rect 301044 180752 301096 180761
rect 306840 180795 306892 180804
rect 306840 180761 306849 180795
rect 306849 180761 306883 180795
rect 306883 180761 306892 180795
rect 306840 180752 306892 180761
rect 317512 180752 317564 180804
rect 317696 180752 317748 180804
rect 245660 180684 245712 180736
rect 245384 180616 245436 180668
rect 245844 180616 245896 180668
rect 245752 179435 245804 179444
rect 245752 179401 245761 179435
rect 245761 179401 245795 179435
rect 245795 179401 245804 179435
rect 245752 179392 245804 179401
rect 267832 179367 267884 179376
rect 267832 179333 267841 179367
rect 267841 179333 267875 179367
rect 267875 179333 267884 179367
rect 267832 179324 267884 179333
rect 266728 178780 266780 178832
rect 294236 178712 294288 178764
rect 294420 178712 294472 178764
rect 295524 178712 295576 178764
rect 295708 178712 295760 178764
rect 296812 178712 296864 178764
rect 296996 178712 297048 178764
rect 266728 178644 266780 178696
rect 247132 176740 247184 176792
rect 232228 176672 232280 176724
rect 250260 176740 250312 176792
rect 299848 176783 299900 176792
rect 299848 176749 299857 176783
rect 299857 176749 299891 176783
rect 299891 176749 299900 176783
rect 299848 176740 299900 176749
rect 302608 176740 302660 176792
rect 247224 176672 247276 176724
rect 250076 176672 250128 176724
rect 310888 176740 310940 176792
rect 389548 176740 389600 176792
rect 232320 176604 232372 176656
rect 235080 176604 235132 176656
rect 302608 176604 302660 176656
rect 310796 176604 310848 176656
rect 389456 176604 389508 176656
rect 235080 176468 235132 176520
rect 239128 176468 239180 176520
rect 460112 176511 460164 176520
rect 460112 176477 460121 176511
rect 460121 176477 460155 176511
rect 460155 176477 460164 176511
rect 460112 176468 460164 176477
rect 372712 176400 372764 176452
rect 372804 176400 372856 176452
rect 375840 176400 375892 176452
rect 375932 176400 375984 176452
rect 239128 176332 239180 176384
rect 366824 174020 366876 174072
rect 367008 174020 367060 174072
rect 230848 173884 230900 173936
rect 231032 173884 231084 173936
rect 236276 173884 236328 173936
rect 236460 173884 236512 173936
rect 259736 173884 259788 173936
rect 259920 173884 259972 173936
rect 265256 173884 265308 173936
rect 265348 173884 265400 173936
rect 270500 173884 270552 173936
rect 270776 173884 270828 173936
rect 281724 173884 281776 173936
rect 281908 173884 281960 173936
rect 284668 173884 284720 173936
rect 284852 173884 284904 173936
rect 288716 173884 288768 173936
rect 288900 173884 288952 173936
rect 323308 173884 323360 173936
rect 323492 173884 323544 173936
rect 324596 173884 324648 173936
rect 324688 173884 324740 173936
rect 325884 173884 325936 173936
rect 325976 173884 326028 173936
rect 327172 173884 327224 173936
rect 327264 173884 327316 173936
rect 357440 173884 357492 173936
rect 357716 173884 357768 173936
rect 376944 173884 376996 173936
rect 377036 173884 377088 173936
rect 463884 173884 463936 173936
rect 464068 173884 464120 173936
rect 291660 173723 291712 173732
rect 291660 173689 291669 173723
rect 291669 173689 291703 173723
rect 291703 173689 291712 173723
rect 291660 173680 291712 173689
rect 251180 172524 251232 172576
rect 251548 172524 251600 172576
rect 273536 172567 273588 172576
rect 273536 172533 273545 172567
rect 273545 172533 273579 172567
rect 273579 172533 273588 172567
rect 273536 172524 273588 172533
rect 290004 172567 290056 172576
rect 290004 172533 290013 172567
rect 290013 172533 290047 172567
rect 290047 172533 290056 172567
rect 290004 172524 290056 172533
rect 331588 172524 331640 172576
rect 337108 172524 337160 172576
rect 329932 172456 329984 172508
rect 330208 172456 330260 172508
rect 331588 172388 331640 172440
rect 337108 172388 337160 172440
rect 299756 171096 299808 171148
rect 301044 171139 301096 171148
rect 301044 171105 301053 171139
rect 301053 171105 301087 171139
rect 301087 171105 301096 171139
rect 301044 171096 301096 171105
rect 306840 171139 306892 171148
rect 306840 171105 306849 171139
rect 306849 171105 306883 171139
rect 306883 171105 306892 171139
rect 306840 171096 306892 171105
rect 244372 171028 244424 171080
rect 247224 171028 247276 171080
rect 266636 171071 266688 171080
rect 266636 171037 266645 171071
rect 266645 171037 266679 171071
rect 266679 171037 266688 171071
rect 266636 171028 266688 171037
rect 331588 171071 331640 171080
rect 331588 171037 331597 171071
rect 331597 171037 331631 171071
rect 331631 171037 331640 171071
rect 331588 171028 331640 171037
rect 337108 171071 337160 171080
rect 337108 171037 337117 171071
rect 337117 171037 337151 171071
rect 337151 171037 337160 171071
rect 337108 171028 337160 171037
rect 244556 170960 244608 171012
rect 267832 169779 267884 169788
rect 267832 169745 267841 169779
rect 267841 169745 267875 169779
rect 267875 169745 267884 169779
rect 267832 169736 267884 169745
rect 278872 167016 278924 167068
rect 310796 167016 310848 167068
rect 357532 167016 357584 167068
rect 357716 167016 357768 167068
rect 431316 167016 431368 167068
rect 431500 167016 431552 167068
rect 278780 166880 278832 166932
rect 310888 166880 310940 166932
rect 341064 164908 341116 164960
rect 341248 164908 341300 164960
rect 251272 164296 251324 164348
rect 251180 164228 251232 164280
rect 235080 164203 235132 164212
rect 235080 164169 235089 164203
rect 235089 164169 235123 164203
rect 235123 164169 235132 164203
rect 235080 164160 235132 164169
rect 236276 164160 236328 164212
rect 236460 164160 236512 164212
rect 285956 164228 286008 164280
rect 251272 164160 251324 164212
rect 270684 164160 270736 164212
rect 251364 164092 251416 164144
rect 270776 164092 270828 164144
rect 340880 164160 340932 164212
rect 341064 164160 341116 164212
rect 367008 164203 367060 164212
rect 367008 164169 367017 164203
rect 367017 164169 367051 164203
rect 367051 164169 367060 164203
rect 367008 164160 367060 164169
rect 372528 164160 372580 164212
rect 372804 164160 372856 164212
rect 375932 164160 375984 164212
rect 286140 164092 286192 164144
rect 230664 162800 230716 162852
rect 230756 162800 230808 162852
rect 250168 162800 250220 162852
rect 250260 162800 250312 162852
rect 251364 162800 251416 162852
rect 251640 162800 251692 162852
rect 393688 162800 393740 162852
rect 330116 162732 330168 162784
rect 247132 161483 247184 161492
rect 247132 161449 247141 161483
rect 247141 161449 247175 161483
rect 247175 161449 247184 161483
rect 247132 161440 247184 161449
rect 265164 161440 265216 161492
rect 265256 161440 265308 161492
rect 266820 161440 266872 161492
rect 294328 161440 294380 161492
rect 294420 161440 294472 161492
rect 295616 161440 295668 161492
rect 295708 161440 295760 161492
rect 296904 161440 296956 161492
rect 296996 161440 297048 161492
rect 331680 161440 331732 161492
rect 337292 161440 337344 161492
rect 286140 161372 286192 161424
rect 265164 160012 265216 160064
rect 272156 160012 272208 160064
rect 378232 157700 378284 157752
rect 386328 157700 386380 157752
rect 306380 157496 306432 157548
rect 315948 157496 316000 157548
rect 336740 157496 336792 157548
rect 346308 157496 346360 157548
rect 417884 157496 417936 157548
rect 418160 157496 418212 157548
rect 437204 157496 437256 157548
rect 437480 157496 437532 157548
rect 267740 157428 267792 157480
rect 357624 157360 357676 157412
rect 267740 157292 267792 157344
rect 325976 157224 326028 157276
rect 460204 157428 460256 157480
rect 460020 157292 460072 157344
rect 357716 157224 357768 157276
rect 325976 157088 326028 157140
rect 299756 156612 299808 156664
rect 299940 156612 299992 156664
rect 245844 156544 245896 156596
rect 246028 156544 246080 156596
rect 367008 154683 367060 154692
rect 367008 154649 367017 154683
rect 367017 154649 367051 154683
rect 367051 154649 367060 154683
rect 367008 154640 367060 154649
rect 235080 154615 235132 154624
rect 235080 154581 235089 154615
rect 235089 154581 235123 154615
rect 235123 154581 235132 154615
rect 235080 154572 235132 154581
rect 375840 154615 375892 154624
rect 375840 154581 375849 154615
rect 375849 154581 375883 154615
rect 375883 154581 375892 154615
rect 375840 154572 375892 154581
rect 232412 154504 232464 154556
rect 259736 154547 259788 154556
rect 259736 154513 259745 154547
rect 259745 154513 259779 154547
rect 259779 154513 259788 154547
rect 259736 154504 259788 154513
rect 366732 154504 366784 154556
rect 367008 154504 367060 154556
rect 247132 153212 247184 153264
rect 337292 153212 337344 153264
rect 393596 153255 393648 153264
rect 393596 153221 393605 153255
rect 393605 153221 393639 153255
rect 393639 153221 393648 153255
rect 393596 153212 393648 153221
rect 247040 153144 247092 153196
rect 270776 153144 270828 153196
rect 270868 153144 270920 153196
rect 273536 153187 273588 153196
rect 273536 153153 273545 153187
rect 273545 153153 273579 153187
rect 273579 153153 273588 153187
rect 273536 153144 273588 153153
rect 290004 153144 290056 153196
rect 290096 153144 290148 153196
rect 291476 153144 291528 153196
rect 291568 153144 291620 153196
rect 294236 153144 294288 153196
rect 294328 153144 294380 153196
rect 310796 153187 310848 153196
rect 310796 153153 310805 153187
rect 310805 153153 310839 153187
rect 310839 153153 310848 153187
rect 310796 153144 310848 153153
rect 337200 153144 337252 153196
rect 266820 151784 266872 151836
rect 285956 151827 286008 151836
rect 285956 151793 285965 151827
rect 285965 151793 285999 151827
rect 285999 151793 286008 151827
rect 285956 151784 286008 151793
rect 3332 151716 3384 151768
rect 24124 151716 24176 151768
rect 266820 151648 266872 151700
rect 245752 150424 245804 150476
rect 246120 150424 246172 150476
rect 265348 150467 265400 150476
rect 265348 150433 265357 150467
rect 265357 150433 265391 150467
rect 265391 150433 265400 150467
rect 265348 150424 265400 150433
rect 296628 150356 296680 150408
rect 296904 150356 296956 150408
rect 393596 148495 393648 148504
rect 393596 148461 393605 148495
rect 393605 148461 393639 148495
rect 393639 148461 393648 148495
rect 393596 148452 393648 148461
rect 281724 148359 281776 148368
rect 281724 148325 281733 148359
rect 281733 148325 281767 148359
rect 281767 148325 281776 148359
rect 281724 148316 281776 148325
rect 272340 148291 272392 148300
rect 272340 148257 272349 148291
rect 272349 148257 272383 148291
rect 272383 148257 272392 148291
rect 272340 148248 272392 148257
rect 235080 147704 235132 147756
rect 463792 147704 463844 147756
rect 357532 147636 357584 147688
rect 357716 147636 357768 147688
rect 235080 147568 235132 147620
rect 259736 147611 259788 147620
rect 259736 147577 259745 147611
rect 259745 147577 259779 147611
rect 259779 147577 259788 147611
rect 259736 147568 259788 147577
rect 310796 147611 310848 147620
rect 310796 147577 310805 147611
rect 310805 147577 310839 147611
rect 310839 147577 310848 147611
rect 310796 147568 310848 147577
rect 331404 146047 331456 146056
rect 331404 146013 331413 146047
rect 331413 146013 331447 146047
rect 331447 146013 331456 146047
rect 331404 146004 331456 146013
rect 232320 145027 232372 145036
rect 232320 144993 232329 145027
rect 232329 144993 232363 145027
rect 232363 144993 232372 145027
rect 232320 144984 232372 144993
rect 330208 144959 330260 144968
rect 330208 144925 330217 144959
rect 330217 144925 330251 144959
rect 330251 144925 330260 144959
rect 330208 144916 330260 144925
rect 463700 144959 463752 144968
rect 463700 144925 463709 144959
rect 463709 144925 463743 144959
rect 463743 144925 463752 144959
rect 463700 144916 463752 144925
rect 267740 144848 267792 144900
rect 267924 144848 267976 144900
rect 273536 144891 273588 144900
rect 273536 144857 273545 144891
rect 273545 144857 273579 144891
rect 273579 144857 273588 144891
rect 273536 144848 273588 144857
rect 284668 144848 284720 144900
rect 284760 144848 284812 144900
rect 323400 144848 323452 144900
rect 323492 144848 323544 144900
rect 324596 144848 324648 144900
rect 324780 144848 324832 144900
rect 325884 144848 325936 144900
rect 326068 144848 326120 144900
rect 357624 144891 357676 144900
rect 357624 144857 357633 144891
rect 357633 144857 357667 144891
rect 357667 144857 357676 144891
rect 357624 144848 357676 144857
rect 367008 144891 367060 144900
rect 367008 144857 367017 144891
rect 367017 144857 367051 144891
rect 367051 144857 367060 144891
rect 367008 144848 367060 144857
rect 459928 144848 459980 144900
rect 460204 144848 460256 144900
rect 251364 143624 251416 143676
rect 251548 143624 251600 143676
rect 281724 143599 281776 143608
rect 281724 143565 281733 143599
rect 281733 143565 281767 143599
rect 281767 143565 281776 143599
rect 281724 143556 281776 143565
rect 230848 143531 230900 143540
rect 230848 143497 230857 143531
rect 230857 143497 230891 143531
rect 230891 143497 230900 143531
rect 230848 143488 230900 143497
rect 232320 143531 232372 143540
rect 232320 143497 232329 143531
rect 232329 143497 232363 143531
rect 232363 143497 232372 143531
rect 232320 143488 232372 143497
rect 245844 143531 245896 143540
rect 245844 143497 245853 143531
rect 245853 143497 245887 143531
rect 245887 143497 245896 143531
rect 245844 143488 245896 143497
rect 250168 143531 250220 143540
rect 250168 143497 250177 143531
rect 250177 143497 250211 143531
rect 250211 143497 250220 143531
rect 250168 143488 250220 143497
rect 329932 143488 329984 143540
rect 330208 143488 330260 143540
rect 393688 142128 393740 142180
rect 251364 142103 251416 142112
rect 251364 142069 251373 142103
rect 251373 142069 251407 142103
rect 251407 142069 251416 142103
rect 251364 142060 251416 142069
rect 296812 140700 296864 140752
rect 296996 140700 297048 140752
rect 324780 139927 324832 139936
rect 324780 139893 324789 139927
rect 324789 139893 324823 139927
rect 324823 139893 324832 139927
rect 324780 139884 324832 139893
rect 296996 139340 297048 139392
rect 341248 138660 341300 138712
rect 302516 138524 302568 138576
rect 302700 138524 302752 138576
rect 244372 138048 244424 138100
rect 235080 137980 235132 138032
rect 259644 137980 259696 138032
rect 259828 137980 259880 138032
rect 310888 138048 310940 138100
rect 463700 137980 463752 138032
rect 244372 137912 244424 137964
rect 245844 137955 245896 137964
rect 245844 137921 245853 137955
rect 245853 137921 245887 137955
rect 245887 137921 245896 137955
rect 245844 137912 245896 137921
rect 250168 137955 250220 137964
rect 250168 137921 250177 137955
rect 250177 137921 250211 137955
rect 250211 137921 250220 137955
rect 250168 137912 250220 137921
rect 310796 137912 310848 137964
rect 357624 137955 357676 137964
rect 357624 137921 357633 137955
rect 357633 137921 357667 137955
rect 357667 137921 357676 137955
rect 357624 137912 357676 137921
rect 463884 137912 463936 137964
rect 235080 137844 235132 137896
rect 285772 137708 285824 137760
rect 286140 137708 286192 137760
rect 326068 137751 326120 137760
rect 326068 137717 326077 137751
rect 326077 137717 326111 137751
rect 326111 137717 326120 137751
rect 326068 137708 326120 137717
rect 299756 137368 299808 137420
rect 299940 137368 299992 137420
rect 2780 136484 2832 136536
rect 5080 136484 5132 136536
rect 367008 135371 367060 135380
rect 367008 135337 367017 135371
rect 367017 135337 367051 135371
rect 367051 135337 367060 135371
rect 367008 135328 367060 135337
rect 273536 135260 273588 135312
rect 273628 135260 273680 135312
rect 337108 135192 337160 135244
rect 337200 135192 337252 135244
rect 339776 135235 339828 135244
rect 339776 135201 339785 135235
rect 339785 135201 339819 135235
rect 339819 135201 339828 135235
rect 339776 135192 339828 135201
rect 357532 135192 357584 135244
rect 357716 135192 357768 135244
rect 367008 135235 367060 135244
rect 367008 135201 367017 135235
rect 367017 135201 367051 135235
rect 367051 135201 367060 135235
rect 367008 135192 367060 135201
rect 378232 134172 378284 134224
rect 386328 134172 386380 134224
rect 456524 134104 456576 134156
rect 457444 134104 457496 134156
rect 309048 134036 309100 134088
rect 315948 134036 316000 134088
rect 437204 134036 437256 134088
rect 437572 134036 437624 134088
rect 475568 134036 475620 134088
rect 482928 134036 482980 134088
rect 417884 133968 417936 134020
rect 418160 133968 418212 134020
rect 230848 133943 230900 133952
rect 230848 133909 230857 133943
rect 230857 133909 230891 133943
rect 230891 133909 230900 133943
rect 230848 133900 230900 133909
rect 232320 133943 232372 133952
rect 232320 133909 232329 133943
rect 232329 133909 232363 133943
rect 232363 133909 232372 133943
rect 232320 133900 232372 133909
rect 324780 133943 324832 133952
rect 324780 133909 324789 133943
rect 324789 133909 324823 133943
rect 324823 133909 324832 133943
rect 324780 133900 324832 133909
rect 326068 133943 326120 133952
rect 326068 133909 326077 133943
rect 326077 133909 326111 133943
rect 326111 133909 326120 133943
rect 326068 133900 326120 133909
rect 331404 133943 331456 133952
rect 331404 133909 331413 133943
rect 331413 133909 331447 133943
rect 331447 133909 331456 133943
rect 331404 133900 331456 133909
rect 270776 133832 270828 133884
rect 271052 133832 271104 133884
rect 299756 133875 299808 133884
rect 299756 133841 299765 133875
rect 299765 133841 299799 133875
rect 299799 133841 299808 133875
rect 299756 133832 299808 133841
rect 301044 133875 301096 133884
rect 301044 133841 301053 133875
rect 301053 133841 301087 133875
rect 301087 133841 301096 133875
rect 301044 133832 301096 133841
rect 357532 133875 357584 133884
rect 357532 133841 357541 133875
rect 357541 133841 357575 133875
rect 357575 133841 357584 133875
rect 357532 133832 357584 133841
rect 251456 132472 251508 132524
rect 289912 132472 289964 132524
rect 290096 132472 290148 132524
rect 295524 132472 295576 132524
rect 295616 132472 295668 132524
rect 259736 132404 259788 132456
rect 262680 132404 262732 132456
rect 245752 131112 245804 131164
rect 245936 131112 245988 131164
rect 393596 131044 393648 131096
rect 393780 131044 393832 131096
rect 375840 130364 375892 130416
rect 376116 130364 376168 130416
rect 463884 130364 463936 130416
rect 464068 130364 464120 130416
rect 291568 129888 291620 129940
rect 291476 129616 291528 129668
rect 306748 128324 306800 128376
rect 306840 128256 306892 128308
rect 341340 128299 341392 128308
rect 341340 128265 341349 128299
rect 341349 128265 341383 128299
rect 341383 128265 341392 128299
rect 341340 128256 341392 128265
rect 310796 125783 310848 125792
rect 310796 125749 310805 125783
rect 310805 125749 310839 125783
rect 310839 125749 310848 125783
rect 310796 125740 310848 125749
rect 367008 125647 367060 125656
rect 367008 125613 367017 125647
rect 367017 125613 367051 125647
rect 367051 125613 367060 125647
rect 367008 125604 367060 125613
rect 377128 125604 377180 125656
rect 377220 125604 377272 125656
rect 235080 125579 235132 125588
rect 235080 125545 235089 125579
rect 235089 125545 235123 125579
rect 235123 125545 235132 125579
rect 235080 125536 235132 125545
rect 236276 125536 236328 125588
rect 236460 125536 236512 125588
rect 330116 125536 330168 125588
rect 330300 125536 330352 125588
rect 331404 125536 331456 125588
rect 331588 125536 331640 125588
rect 337108 125536 337160 125588
rect 337292 125536 337344 125588
rect 375840 125536 375892 125588
rect 339684 124244 339736 124296
rect 289912 124176 289964 124228
rect 290004 124176 290056 124228
rect 299848 124176 299900 124228
rect 301136 124176 301188 124228
rect 357624 124176 357676 124228
rect 232320 124151 232372 124160
rect 232320 124117 232329 124151
rect 232329 124117 232363 124151
rect 232363 124117 232372 124151
rect 232320 124108 232372 124117
rect 247316 124151 247368 124160
rect 247316 124117 247325 124151
rect 247325 124117 247359 124151
rect 247359 124117 247368 124151
rect 247316 124108 247368 124117
rect 377128 124108 377180 124160
rect 456524 123088 456576 123140
rect 457444 123088 457496 123140
rect 306012 123020 306064 123072
rect 314568 123020 314620 123072
rect 369676 123020 369728 123072
rect 376668 123020 376720 123072
rect 417884 122952 417936 123004
rect 419356 122952 419408 123004
rect 437204 122952 437256 123004
rect 437480 122952 437532 123004
rect 259644 122859 259696 122868
rect 259644 122825 259653 122859
rect 259653 122825 259687 122859
rect 259687 122825 259696 122859
rect 259644 122816 259696 122825
rect 262588 122859 262640 122868
rect 262588 122825 262597 122859
rect 262597 122825 262631 122859
rect 262631 122825 262640 122859
rect 262588 122816 262640 122825
rect 251364 122791 251416 122800
rect 251364 122757 251373 122791
rect 251373 122757 251407 122791
rect 251407 122757 251416 122791
rect 251364 122748 251416 122757
rect 270868 122748 270920 122800
rect 285956 122748 286008 122800
rect 286048 122748 286100 122800
rect 288716 122748 288768 122800
rect 288808 122748 288860 122800
rect 294420 122791 294472 122800
rect 294420 122757 294429 122791
rect 294429 122757 294463 122791
rect 294463 122757 294472 122791
rect 294420 122748 294472 122757
rect 295708 122791 295760 122800
rect 295708 122757 295717 122791
rect 295717 122757 295751 122791
rect 295751 122757 295760 122791
rect 295708 122748 295760 122757
rect 303896 122791 303948 122800
rect 303896 122757 303905 122791
rect 303905 122757 303939 122791
rect 303939 122757 303948 122791
rect 303896 122748 303948 122757
rect 324596 122791 324648 122800
rect 324596 122757 324605 122791
rect 324605 122757 324639 122791
rect 324639 122757 324648 122791
rect 324596 122748 324648 122757
rect 325884 122791 325936 122800
rect 325884 122757 325893 122791
rect 325893 122757 325927 122791
rect 325927 122757 325936 122791
rect 325884 122748 325936 122757
rect 339776 122791 339828 122800
rect 339776 122757 339785 122791
rect 339785 122757 339819 122791
rect 339819 122757 339828 122791
rect 339776 122748 339828 122757
rect 372804 122791 372856 122800
rect 372804 122757 372813 122791
rect 372813 122757 372847 122791
rect 372847 122757 372856 122791
rect 372804 122748 372856 122757
rect 296996 122680 297048 122732
rect 2780 122272 2832 122324
rect 4988 122272 5040 122324
rect 310796 121499 310848 121508
rect 310796 121465 310805 121499
rect 310805 121465 310839 121499
rect 310839 121465 310848 121499
rect 310796 121456 310848 121465
rect 389364 121431 389416 121440
rect 389364 121397 389373 121431
rect 389373 121397 389407 121431
rect 389407 121397 389416 121431
rect 389364 121388 389416 121397
rect 291476 120071 291528 120080
rect 291476 120037 291485 120071
rect 291485 120037 291519 120071
rect 291519 120037 291528 120071
rect 291476 120028 291528 120037
rect 393596 120071 393648 120080
rect 393596 120037 393605 120071
rect 393605 120037 393639 120071
rect 393639 120037 393648 120071
rect 393596 120028 393648 120037
rect 278872 118736 278924 118788
rect 341248 118668 341300 118720
rect 341432 118668 341484 118720
rect 278872 118600 278924 118652
rect 339776 118031 339828 118040
rect 339776 117997 339785 118031
rect 339785 117997 339819 118031
rect 339819 117997 339828 118031
rect 339776 117988 339828 117997
rect 295800 116560 295852 116612
rect 235080 115991 235132 116000
rect 235080 115957 235089 115991
rect 235089 115957 235123 115991
rect 235123 115957 235132 115991
rect 235080 115948 235132 115957
rect 245936 115991 245988 116000
rect 245936 115957 245945 115991
rect 245945 115957 245979 115991
rect 245979 115957 245988 115991
rect 245936 115948 245988 115957
rect 375748 115991 375800 116000
rect 375748 115957 375757 115991
rect 375757 115957 375791 115991
rect 375791 115957 375800 115991
rect 375748 115948 375800 115957
rect 341248 115880 341300 115932
rect 366732 115880 366784 115932
rect 367008 115880 367060 115932
rect 232320 114563 232372 114572
rect 232320 114529 232329 114563
rect 232329 114529 232363 114563
rect 232363 114529 232372 114563
rect 232320 114520 232372 114529
rect 244280 114520 244332 114572
rect 244464 114520 244516 114572
rect 245936 114563 245988 114572
rect 245936 114529 245945 114563
rect 245945 114529 245979 114563
rect 245979 114529 245988 114563
rect 245936 114520 245988 114529
rect 247132 114520 247184 114572
rect 265164 114520 265216 114572
rect 265256 114520 265308 114572
rect 377036 114563 377088 114572
rect 377036 114529 377045 114563
rect 377045 114529 377079 114563
rect 377079 114529 377088 114563
rect 377036 114520 377088 114529
rect 272248 114452 272300 114504
rect 272340 114452 272392 114504
rect 337200 114452 337252 114504
rect 463976 114452 464028 114504
rect 326068 114384 326120 114436
rect 301136 113228 301188 113280
rect 251456 113160 251508 113212
rect 259736 113160 259788 113212
rect 259920 113160 259972 113212
rect 270776 113203 270828 113212
rect 270776 113169 270785 113203
rect 270785 113169 270819 113203
rect 270819 113169 270828 113203
rect 270776 113160 270828 113169
rect 294420 113203 294472 113212
rect 294420 113169 294429 113203
rect 294429 113169 294463 113203
rect 294463 113169 294472 113203
rect 294420 113160 294472 113169
rect 301044 113160 301096 113212
rect 303896 113203 303948 113212
rect 303896 113169 303905 113203
rect 303905 113169 303939 113203
rect 303939 113169 303948 113203
rect 303896 113160 303948 113169
rect 324596 113203 324648 113212
rect 324596 113169 324605 113203
rect 324605 113169 324639 113203
rect 324639 113169 324648 113203
rect 324596 113160 324648 113169
rect 372804 113203 372856 113212
rect 372804 113169 372813 113203
rect 372813 113169 372847 113203
rect 372847 113169 372856 113203
rect 372804 113160 372856 113169
rect 244280 113092 244332 113144
rect 285956 113135 286008 113144
rect 285956 113101 285965 113135
rect 285965 113101 285999 113135
rect 285999 113101 286008 113135
rect 285956 113092 286008 113101
rect 296996 112820 297048 112872
rect 296996 112684 297048 112736
rect 310796 111800 310848 111852
rect 310980 111800 311032 111852
rect 290096 111732 290148 111784
rect 295708 111775 295760 111784
rect 295708 111741 295717 111775
rect 295717 111741 295751 111775
rect 295751 111741 295760 111775
rect 295708 111732 295760 111741
rect 306288 110780 306340 110832
rect 315948 110780 316000 110832
rect 248420 110712 248472 110764
rect 254124 110712 254176 110764
rect 456524 110712 456576 110764
rect 457444 110712 457496 110764
rect 259368 110576 259420 110628
rect 267648 110576 267700 110628
rect 417884 110576 417936 110628
rect 418160 110576 418212 110628
rect 437204 110576 437256 110628
rect 437480 110576 437532 110628
rect 291476 110483 291528 110492
rect 291476 110449 291485 110483
rect 291485 110449 291519 110483
rect 291519 110449 291528 110483
rect 291476 110440 291528 110449
rect 393596 110483 393648 110492
rect 393596 110449 393605 110483
rect 393605 110449 393639 110483
rect 393639 110449 393648 110483
rect 393596 110440 393648 110449
rect 262588 109692 262640 109744
rect 357716 109692 357768 109744
rect 265164 109012 265216 109064
rect 375748 109012 375800 109064
rect 377036 109012 377088 109064
rect 265256 108944 265308 108996
rect 375840 108944 375892 108996
rect 377128 108944 377180 108996
rect 323400 108035 323452 108044
rect 323400 108001 323409 108035
rect 323409 108001 323443 108035
rect 323443 108001 323452 108035
rect 323400 107992 323452 108001
rect 247132 106292 247184 106344
rect 341156 106335 341208 106344
rect 341156 106301 341165 106335
rect 341165 106301 341199 106335
rect 341199 106301 341208 106335
rect 341156 106292 341208 106301
rect 235080 106267 235132 106276
rect 235080 106233 235089 106267
rect 235089 106233 235123 106267
rect 235123 106233 235132 106267
rect 235080 106224 235132 106233
rect 236276 106224 236328 106276
rect 236460 106224 236512 106276
rect 245936 106267 245988 106276
rect 245936 106233 245945 106267
rect 245945 106233 245979 106267
rect 245979 106233 245988 106267
rect 245936 106224 245988 106233
rect 284760 106224 284812 106276
rect 284852 106224 284904 106276
rect 367008 106267 367060 106276
rect 367008 106233 367017 106267
rect 367017 106233 367051 106267
rect 367051 106233 367060 106267
rect 367008 106224 367060 106233
rect 459928 106224 459980 106276
rect 460112 106224 460164 106276
rect 247132 106156 247184 106208
rect 262496 104907 262548 104916
rect 262496 104873 262505 104907
rect 262505 104873 262539 104907
rect 262539 104873 262548 104907
rect 262496 104864 262548 104873
rect 267740 104864 267792 104916
rect 267832 104864 267884 104916
rect 270684 104864 270736 104916
rect 270776 104864 270828 104916
rect 299664 104864 299716 104916
rect 299756 104864 299808 104916
rect 325976 104864 326028 104916
rect 326068 104864 326120 104916
rect 337016 104907 337068 104916
rect 337016 104873 337025 104907
rect 337025 104873 337059 104907
rect 337059 104873 337068 104907
rect 337016 104864 337068 104873
rect 393596 104864 393648 104916
rect 463884 104907 463936 104916
rect 463884 104873 463893 104907
rect 463893 104873 463927 104907
rect 463927 104873 463936 104907
rect 463884 104864 463936 104873
rect 232320 104839 232372 104848
rect 232320 104805 232329 104839
rect 232329 104805 232363 104839
rect 232363 104805 232372 104839
rect 232320 104796 232372 104805
rect 324596 104839 324648 104848
rect 324596 104805 324605 104839
rect 324605 104805 324639 104839
rect 324639 104805 324648 104839
rect 324596 104796 324648 104805
rect 337016 104728 337068 104780
rect 393688 104728 393740 104780
rect 290004 104227 290056 104236
rect 290004 104193 290013 104227
rect 290013 104193 290047 104227
rect 290047 104193 290056 104227
rect 290004 104184 290056 104193
rect 244372 103547 244424 103556
rect 244372 103513 244381 103547
rect 244381 103513 244415 103547
rect 244415 103513 244424 103547
rect 244372 103504 244424 103513
rect 286048 103504 286100 103556
rect 291476 103504 291528 103556
rect 294420 103504 294472 103556
rect 296904 103504 296956 103556
rect 296996 103504 297048 103556
rect 389364 103547 389416 103556
rect 389364 103513 389373 103547
rect 389373 103513 389407 103547
rect 389407 103513 389416 103547
rect 389364 103504 389416 103513
rect 247132 103479 247184 103488
rect 247132 103445 247141 103479
rect 247141 103445 247175 103479
rect 247175 103445 247184 103479
rect 247132 103436 247184 103445
rect 291660 103436 291712 103488
rect 294604 103436 294656 103488
rect 327172 103479 327224 103488
rect 327172 103445 327181 103479
rect 327181 103445 327215 103479
rect 327215 103445 327224 103479
rect 327172 103436 327224 103445
rect 331404 103479 331456 103488
rect 331404 103445 331413 103479
rect 331413 103445 331447 103479
rect 331447 103445 331456 103479
rect 331404 103436 331456 103445
rect 372804 103436 372856 103488
rect 244372 103368 244424 103420
rect 244556 103368 244608 103420
rect 317696 103411 317748 103420
rect 317696 103377 317705 103411
rect 317705 103377 317739 103411
rect 317739 103377 317748 103411
rect 317696 103368 317748 103377
rect 330116 103411 330168 103420
rect 330116 103377 330125 103411
rect 330125 103377 330159 103411
rect 330159 103377 330168 103411
rect 330116 103368 330168 103377
rect 310980 102212 311032 102264
rect 295892 102144 295944 102196
rect 310888 102144 310940 102196
rect 393688 100648 393740 100700
rect 267832 99424 267884 99476
rect 377128 99424 377180 99476
rect 341156 99356 341208 99408
rect 267740 99288 267792 99340
rect 341248 99288 341300 99340
rect 357624 99331 357676 99340
rect 357624 99297 357633 99331
rect 357633 99297 357667 99331
rect 357667 99297 357676 99331
rect 357624 99288 357676 99297
rect 377128 99288 377180 99340
rect 310888 98676 310940 98728
rect 330208 98676 330260 98728
rect 389364 98676 389416 98728
rect 290004 97971 290056 97980
rect 290004 97937 290013 97971
rect 290013 97937 290047 97971
rect 290047 97937 290056 97971
rect 290004 97928 290056 97937
rect 367008 96747 367060 96756
rect 367008 96713 367017 96747
rect 367017 96713 367051 96747
rect 367051 96713 367060 96747
rect 367008 96704 367060 96713
rect 235080 96679 235132 96688
rect 235080 96645 235089 96679
rect 235089 96645 235123 96679
rect 235123 96645 235132 96679
rect 235080 96636 235132 96645
rect 245936 96679 245988 96688
rect 245936 96645 245945 96679
rect 245945 96645 245979 96679
rect 245979 96645 245988 96679
rect 245936 96636 245988 96645
rect 284852 96636 284904 96688
rect 284760 96568 284812 96620
rect 327172 96611 327224 96620
rect 327172 96577 327181 96611
rect 327181 96577 327215 96611
rect 327215 96577 327224 96611
rect 327172 96568 327224 96577
rect 265256 95319 265308 95328
rect 265256 95285 265265 95319
rect 265265 95285 265299 95319
rect 265299 95285 265308 95319
rect 265256 95276 265308 95285
rect 272340 95276 272392 95328
rect 299756 95276 299808 95328
rect 232320 95251 232372 95260
rect 232320 95217 232329 95251
rect 232329 95217 232363 95251
rect 232363 95217 232372 95251
rect 232320 95208 232372 95217
rect 262496 95208 262548 95260
rect 262588 95208 262640 95260
rect 270684 95208 270736 95260
rect 270776 95208 270828 95260
rect 272248 95208 272300 95260
rect 299848 95208 299900 95260
rect 317788 95208 317840 95260
rect 323400 95251 323452 95260
rect 323400 95217 323409 95251
rect 323409 95217 323443 95251
rect 323443 95217 323452 95251
rect 323400 95208 323452 95217
rect 324596 95251 324648 95260
rect 324596 95217 324605 95251
rect 324605 95217 324639 95251
rect 324639 95217 324648 95251
rect 324596 95208 324648 95217
rect 337200 95251 337252 95260
rect 337200 95217 337209 95251
rect 337209 95217 337243 95251
rect 337243 95217 337252 95251
rect 337200 95208 337252 95217
rect 463700 95208 463752 95260
rect 463884 95208 463936 95260
rect 259644 95140 259696 95192
rect 296904 95140 296956 95192
rect 296996 95140 297048 95192
rect 463700 94163 463752 94172
rect 463700 94129 463709 94163
rect 463709 94129 463743 94163
rect 463743 94129 463752 94163
rect 463700 94120 463752 94129
rect 247224 93848 247276 93900
rect 331404 93891 331456 93900
rect 331404 93857 331413 93891
rect 331413 93857 331447 93891
rect 331447 93857 331456 93891
rect 331404 93848 331456 93857
rect 262588 93823 262640 93832
rect 262588 93789 262597 93823
rect 262597 93789 262631 93823
rect 262631 93789 262640 93823
rect 262588 93780 262640 93789
rect 290004 93823 290056 93832
rect 290004 93789 290013 93823
rect 290013 93789 290047 93823
rect 290047 93789 290056 93823
rect 290004 93780 290056 93789
rect 330116 93780 330168 93832
rect 245752 92488 245804 92540
rect 245844 92488 245896 92540
rect 265256 92531 265308 92540
rect 265256 92497 265265 92531
rect 265265 92497 265299 92531
rect 265299 92497 265308 92531
rect 265256 92488 265308 92497
rect 270776 90380 270828 90432
rect 272248 90380 272300 90432
rect 317788 89700 317840 89752
rect 357532 89700 357584 89752
rect 357716 89700 357768 89752
rect 431316 89700 431368 89752
rect 431500 89700 431552 89752
rect 310796 89675 310848 89684
rect 310796 89641 310805 89675
rect 310805 89641 310839 89675
rect 310839 89641 310848 89675
rect 310796 89632 310848 89641
rect 389272 89675 389324 89684
rect 389272 89641 389281 89675
rect 389281 89641 389315 89675
rect 389315 89641 389324 89675
rect 389272 89632 389324 89641
rect 317880 89564 317932 89616
rect 281724 88952 281776 89004
rect 366916 87227 366968 87236
rect 366916 87193 366925 87227
rect 366925 87193 366959 87227
rect 366959 87193 366968 87227
rect 366916 87184 366968 87193
rect 417884 87116 417936 87168
rect 418620 87116 418672 87168
rect 454040 87116 454092 87168
rect 463424 87116 463476 87168
rect 463700 87116 463752 87168
rect 467932 87116 467984 87168
rect 494612 87116 494664 87168
rect 502248 87116 502300 87168
rect 336740 87048 336792 87100
rect 346308 87048 346360 87100
rect 366916 87091 366968 87100
rect 366916 87057 366925 87091
rect 366925 87057 366959 87091
rect 366959 87057 366968 87091
rect 366916 87048 366968 87057
rect 379060 87048 379112 87100
rect 386236 87048 386288 87100
rect 396080 87048 396132 87100
rect 405556 87048 405608 87100
rect 437204 87048 437256 87100
rect 437480 87048 437532 87100
rect 235080 86955 235132 86964
rect 235080 86921 235089 86955
rect 235089 86921 235123 86955
rect 235123 86921 235132 86955
rect 235080 86912 235132 86921
rect 236276 86955 236328 86964
rect 236276 86921 236285 86955
rect 236285 86921 236319 86955
rect 236319 86921 236328 86955
rect 236276 86912 236328 86921
rect 284576 86912 284628 86964
rect 284760 86912 284812 86964
rect 323308 86912 323360 86964
rect 323400 86912 323452 86964
rect 324596 86912 324648 86964
rect 327172 86912 327224 86964
rect 341156 86912 341208 86964
rect 357624 86955 357676 86964
rect 357624 86921 357633 86955
rect 357633 86921 357667 86955
rect 357667 86921 357676 86955
rect 357624 86912 357676 86921
rect 375840 86955 375892 86964
rect 375840 86921 375849 86955
rect 375849 86921 375883 86955
rect 375883 86921 375892 86955
rect 375840 86912 375892 86921
rect 377128 86955 377180 86964
rect 377128 86921 377137 86955
rect 377137 86921 377171 86955
rect 377171 86921 377180 86955
rect 377128 86912 377180 86921
rect 431316 86955 431368 86964
rect 431316 86921 431325 86955
rect 431325 86921 431359 86955
rect 431359 86921 431368 86955
rect 431316 86912 431368 86921
rect 324688 86844 324740 86896
rect 327264 86844 327316 86896
rect 393596 86887 393648 86896
rect 393596 86853 393605 86887
rect 393605 86853 393639 86887
rect 393639 86853 393648 86887
rect 393596 86844 393648 86853
rect 267740 85552 267792 85604
rect 291568 85552 291620 85604
rect 291660 85552 291712 85604
rect 294420 85552 294472 85604
rect 294604 85552 294656 85604
rect 306840 85552 306892 85604
rect 306932 85552 306984 85604
rect 331404 85552 331456 85604
rect 331680 85552 331732 85604
rect 463884 85552 463936 85604
rect 232320 85527 232372 85536
rect 232320 85493 232329 85527
rect 232329 85493 232363 85527
rect 232363 85493 232372 85527
rect 232320 85484 232372 85493
rect 310796 85527 310848 85536
rect 310796 85493 310805 85527
rect 310805 85493 310839 85527
rect 310839 85493 310848 85527
rect 310796 85484 310848 85493
rect 367008 85527 367060 85536
rect 367008 85493 367017 85527
rect 367017 85493 367051 85527
rect 367051 85493 367060 85527
rect 367008 85484 367060 85493
rect 267832 85416 267884 85468
rect 286140 84940 286192 84992
rect 262680 84192 262732 84244
rect 290096 84192 290148 84244
rect 329932 84235 329984 84244
rect 329932 84201 329941 84235
rect 329941 84201 329975 84235
rect 329975 84201 329984 84235
rect 329932 84192 329984 84201
rect 290188 84056 290240 84108
rect 295708 82832 295760 82884
rect 295892 82832 295944 82884
rect 267832 82807 267884 82816
rect 267832 82773 267841 82807
rect 267841 82773 267875 82807
rect 267875 82773 267884 82807
rect 267832 82764 267884 82773
rect 278872 80112 278924 80164
rect 339776 80112 339828 80164
rect 247224 80044 247276 80096
rect 389364 80044 389416 80096
rect 273536 80019 273588 80028
rect 273536 79985 273545 80019
rect 273545 79985 273579 80019
rect 273579 79985 273588 80019
rect 273536 79976 273588 79985
rect 278872 79976 278924 80028
rect 339776 79976 339828 80028
rect 389456 79908 389508 79960
rect 2780 79772 2832 79824
rect 4896 79772 4948 79824
rect 235080 77299 235132 77308
rect 235080 77265 235089 77299
rect 235089 77265 235123 77299
rect 235123 77265 235132 77299
rect 235080 77256 235132 77265
rect 236276 77299 236328 77308
rect 236276 77265 236285 77299
rect 236285 77265 236319 77299
rect 236319 77265 236328 77299
rect 236276 77256 236328 77265
rect 259736 77299 259788 77308
rect 259736 77265 259745 77299
rect 259745 77265 259779 77299
rect 259779 77265 259788 77299
rect 259736 77256 259788 77265
rect 266636 77256 266688 77308
rect 266728 77256 266780 77308
rect 270776 77256 270828 77308
rect 272248 77256 272300 77308
rect 296996 77324 297048 77376
rect 299848 77324 299900 77376
rect 330024 77324 330076 77376
rect 302516 77256 302568 77308
rect 302608 77256 302660 77308
rect 306748 77256 306800 77308
rect 306840 77256 306892 77308
rect 341064 77299 341116 77308
rect 341064 77265 341073 77299
rect 341073 77265 341107 77299
rect 341107 77265 341116 77299
rect 341064 77256 341116 77265
rect 357716 77256 357768 77308
rect 372712 77299 372764 77308
rect 372712 77265 372721 77299
rect 372721 77265 372755 77299
rect 372755 77265 372764 77299
rect 372712 77256 372764 77265
rect 375840 77299 375892 77308
rect 375840 77265 375849 77299
rect 375849 77265 375883 77299
rect 375883 77265 375892 77299
rect 375840 77256 375892 77265
rect 377128 77299 377180 77308
rect 377128 77265 377137 77299
rect 377137 77265 377171 77299
rect 377171 77265 377180 77299
rect 377128 77256 377180 77265
rect 431316 77299 431368 77308
rect 431316 77265 431325 77299
rect 431325 77265 431359 77299
rect 431359 77265 431368 77299
rect 431316 77256 431368 77265
rect 251456 77188 251508 77240
rect 296812 77188 296864 77240
rect 299848 77188 299900 77240
rect 330024 77188 330076 77240
rect 341064 77163 341116 77172
rect 341064 77129 341073 77163
rect 341073 77129 341107 77163
rect 341107 77129 341116 77163
rect 341064 77120 341116 77129
rect 431316 77163 431368 77172
rect 431316 77129 431325 77163
rect 431325 77129 431359 77163
rect 431359 77129 431368 77163
rect 431316 77120 431368 77129
rect 378232 76236 378284 76288
rect 386328 76236 386380 76288
rect 434720 76100 434772 76152
rect 437480 76100 437532 76152
rect 463700 76100 463752 76152
rect 467932 76100 467984 76152
rect 417884 76032 417936 76084
rect 419356 76032 419408 76084
rect 270500 75964 270552 76016
rect 275376 75964 275428 76016
rect 232320 75939 232372 75948
rect 232320 75905 232329 75939
rect 232329 75905 232363 75939
rect 232363 75905 232372 75939
rect 232320 75896 232372 75905
rect 273536 75939 273588 75948
rect 273536 75905 273545 75939
rect 273545 75905 273579 75939
rect 273579 75905 273588 75939
rect 273536 75896 273588 75905
rect 281816 75939 281868 75948
rect 281816 75905 281825 75939
rect 281825 75905 281859 75939
rect 281859 75905 281868 75939
rect 281816 75896 281868 75905
rect 286140 75896 286192 75948
rect 310796 75939 310848 75948
rect 310796 75905 310805 75939
rect 310805 75905 310839 75939
rect 310839 75905 310848 75939
rect 310796 75896 310848 75905
rect 317696 75896 317748 75948
rect 317972 75896 318024 75948
rect 331404 75896 331456 75948
rect 331680 75896 331732 75948
rect 367008 75939 367060 75948
rect 367008 75905 367017 75939
rect 367017 75905 367051 75939
rect 367051 75905 367060 75939
rect 367008 75896 367060 75905
rect 389456 75828 389508 75880
rect 303896 74672 303948 74724
rect 291384 74536 291436 74588
rect 291568 74536 291620 74588
rect 303896 74536 303948 74588
rect 294420 74468 294472 74520
rect 393688 74511 393740 74520
rect 393688 74477 393697 74511
rect 393697 74477 393731 74511
rect 393731 74477 393740 74511
rect 393688 74468 393740 74477
rect 245752 73176 245804 73228
rect 245844 73176 245896 73228
rect 247132 73219 247184 73228
rect 247132 73185 247141 73219
rect 247141 73185 247175 73219
rect 247175 73185 247184 73219
rect 247132 73176 247184 73185
rect 267924 73176 267976 73228
rect 272248 70524 272300 70576
rect 270776 70456 270828 70508
rect 327264 70456 327316 70508
rect 375840 70456 375892 70508
rect 377128 70499 377180 70508
rect 377128 70465 377137 70499
rect 377137 70465 377171 70499
rect 377171 70465 377180 70499
rect 377128 70456 377180 70465
rect 270684 70320 270736 70372
rect 327172 70320 327224 70372
rect 375840 70320 375892 70372
rect 341156 70252 341208 70304
rect 245936 67668 245988 67720
rect 235080 67575 235132 67584
rect 235080 67541 235089 67575
rect 235089 67541 235123 67575
rect 235123 67541 235132 67575
rect 235080 67532 235132 67541
rect 236276 67575 236328 67584
rect 236276 67541 236285 67575
rect 236285 67541 236319 67575
rect 236319 67541 236328 67575
rect 236276 67532 236328 67541
rect 357716 67668 357768 67720
rect 265164 67600 265216 67652
rect 265256 67600 265308 67652
rect 272156 67643 272208 67652
rect 272156 67609 272165 67643
rect 272165 67609 272199 67643
rect 272199 67609 272208 67643
rect 272156 67600 272208 67609
rect 281724 67600 281776 67652
rect 281816 67600 281868 67652
rect 291384 67600 291436 67652
rect 291476 67600 291528 67652
rect 299756 67600 299808 67652
rect 299848 67600 299900 67652
rect 301044 67600 301096 67652
rect 301228 67600 301280 67652
rect 329932 67600 329984 67652
rect 330116 67600 330168 67652
rect 357624 67600 357676 67652
rect 377128 67643 377180 67652
rect 377128 67609 377137 67643
rect 377137 67609 377171 67643
rect 377171 67609 377180 67643
rect 377128 67600 377180 67609
rect 431408 67600 431460 67652
rect 459928 67532 459980 67584
rect 460204 67532 460256 67584
rect 245936 67464 245988 67516
rect 389364 66283 389416 66292
rect 389364 66249 389373 66283
rect 389373 66249 389407 66283
rect 389407 66249 389416 66283
rect 389364 66240 389416 66249
rect 232320 66172 232372 66224
rect 244372 66215 244424 66224
rect 244372 66181 244381 66215
rect 244381 66181 244415 66215
rect 244415 66181 244424 66215
rect 244372 66172 244424 66181
rect 245936 66172 245988 66224
rect 265164 66172 265216 66224
rect 273536 66215 273588 66224
rect 273536 66181 273545 66215
rect 273545 66181 273579 66215
rect 273579 66181 273588 66215
rect 273536 66172 273588 66181
rect 302516 66172 302568 66224
rect 302700 66172 302752 66224
rect 306748 66172 306800 66224
rect 306932 66172 306984 66224
rect 310796 66215 310848 66224
rect 310796 66181 310805 66215
rect 310805 66181 310839 66215
rect 310839 66181 310848 66215
rect 310796 66172 310848 66181
rect 323400 66215 323452 66224
rect 323400 66181 323409 66215
rect 323409 66181 323443 66215
rect 323443 66181 323452 66215
rect 323400 66172 323452 66181
rect 327172 66215 327224 66224
rect 327172 66181 327181 66215
rect 327181 66181 327215 66215
rect 327215 66181 327224 66215
rect 327172 66172 327224 66181
rect 367008 66215 367060 66224
rect 367008 66181 367017 66215
rect 367017 66181 367051 66215
rect 367051 66181 367060 66215
rect 367008 66172 367060 66181
rect 246028 66104 246080 66156
rect 267924 64948 267976 65000
rect 251364 64923 251416 64932
rect 251364 64889 251373 64923
rect 251373 64889 251407 64923
rect 251407 64889 251416 64923
rect 251364 64880 251416 64889
rect 267740 64880 267792 64932
rect 294236 64923 294288 64932
rect 294236 64889 294245 64923
rect 294245 64889 294279 64923
rect 294279 64889 294288 64923
rect 294236 64880 294288 64889
rect 295616 64880 295668 64932
rect 295708 64880 295760 64932
rect 393780 64880 393832 64932
rect 3332 64812 3384 64864
rect 31024 64812 31076 64864
rect 378232 63860 378284 63912
rect 386328 63860 386380 63912
rect 417884 63656 417936 63708
rect 418160 63656 418212 63708
rect 437204 63656 437256 63708
rect 437480 63656 437532 63708
rect 456524 63656 456576 63708
rect 456892 63656 456944 63708
rect 303896 63495 303948 63504
rect 303896 63461 303905 63495
rect 303905 63461 303939 63495
rect 303939 63461 303948 63495
rect 303896 63452 303948 63461
rect 235080 62747 235132 62756
rect 235080 62713 235089 62747
rect 235089 62713 235123 62747
rect 235123 62713 235132 62747
rect 235080 62704 235132 62713
rect 259736 62636 259788 62688
rect 259920 62568 259972 62620
rect 262772 61412 262824 61464
rect 262956 61412 263008 61464
rect 281724 61455 281776 61464
rect 281724 61421 281733 61455
rect 281733 61421 281767 61455
rect 281767 61421 281776 61455
rect 281724 61412 281776 61421
rect 295616 61412 295668 61464
rect 330116 61455 330168 61464
rect 330116 61421 330125 61455
rect 330125 61421 330159 61455
rect 330159 61421 330168 61455
rect 330116 61412 330168 61421
rect 267740 60800 267792 60852
rect 324596 60800 324648 60852
rect 337200 60800 337252 60852
rect 339776 60843 339828 60852
rect 339776 60809 339785 60843
rect 339785 60809 339819 60843
rect 339819 60809 339828 60843
rect 339776 60800 339828 60809
rect 266636 60732 266688 60784
rect 230848 60596 230900 60648
rect 325884 60732 325936 60784
rect 267740 60664 267792 60716
rect 310796 60707 310848 60716
rect 310796 60673 310805 60707
rect 310805 60673 310839 60707
rect 310839 60673 310848 60707
rect 310796 60664 310848 60673
rect 324596 60664 324648 60716
rect 266728 60596 266780 60648
rect 325976 60596 326028 60648
rect 337200 60596 337252 60648
rect 270684 58012 270736 58064
rect 284760 58012 284812 58064
rect 236276 57987 236328 57996
rect 236276 57953 236285 57987
rect 236285 57953 236319 57987
rect 236319 57953 236328 57987
rect 236276 57944 236328 57953
rect 272156 57944 272208 57996
rect 272248 57944 272300 57996
rect 291476 58012 291528 58064
rect 270684 57876 270736 57928
rect 284760 57876 284812 57928
rect 291384 57876 291436 57928
rect 357716 57876 357768 57928
rect 460112 57876 460164 57928
rect 330300 57808 330352 57860
rect 389364 57536 389416 57588
rect 288716 57035 288768 57044
rect 288716 57001 288725 57035
rect 288725 57001 288759 57035
rect 288759 57001 288768 57035
rect 288716 56992 288768 57001
rect 232320 56627 232372 56636
rect 232320 56593 232329 56627
rect 232329 56593 232363 56627
rect 232363 56593 232372 56627
rect 232320 56584 232372 56593
rect 244464 56584 244516 56636
rect 250168 56627 250220 56636
rect 250168 56593 250177 56627
rect 250177 56593 250211 56627
rect 250211 56593 250220 56627
rect 250168 56584 250220 56593
rect 273536 56627 273588 56636
rect 273536 56593 273545 56627
rect 273545 56593 273579 56627
rect 273579 56593 273588 56627
rect 273536 56584 273588 56593
rect 323400 56627 323452 56636
rect 323400 56593 323409 56627
rect 323409 56593 323443 56627
rect 323443 56593 323452 56627
rect 323400 56584 323452 56593
rect 327448 56584 327500 56636
rect 339776 56627 339828 56636
rect 339776 56593 339785 56627
rect 339785 56593 339819 56627
rect 339819 56593 339828 56627
rect 339776 56584 339828 56593
rect 259920 56559 259972 56568
rect 259920 56525 259929 56559
rect 259929 56525 259963 56559
rect 259963 56525 259972 56559
rect 259920 56516 259972 56525
rect 310796 56516 310848 56568
rect 310888 56516 310940 56568
rect 341340 56559 341392 56568
rect 341340 56525 341349 56559
rect 341349 56525 341383 56559
rect 341383 56525 341392 56559
rect 341340 56516 341392 56525
rect 317512 55224 317564 55276
rect 317696 55224 317748 55276
rect 393504 55224 393556 55276
rect 393780 55224 393832 55276
rect 247224 55199 247276 55208
rect 247224 55165 247233 55199
rect 247233 55165 247267 55199
rect 247267 55165 247276 55199
rect 247224 55156 247276 55165
rect 250168 53839 250220 53848
rect 250168 53805 250177 53839
rect 250177 53805 250211 53839
rect 250211 53805 250220 53839
rect 250168 53796 250220 53805
rect 303988 53796 304040 53848
rect 278872 51187 278924 51196
rect 278872 51153 278881 51187
rect 278881 51153 278915 51187
rect 278915 51153 278924 51187
rect 278872 51144 278924 51153
rect 375840 51144 375892 51196
rect 232320 51076 232372 51128
rect 273536 51076 273588 51128
rect 337200 51076 337252 51128
rect 232228 51008 232280 51060
rect 375840 51008 375892 51060
rect 265164 50872 265216 50924
rect 273536 50872 273588 50924
rect 341340 50643 341392 50652
rect 341340 50609 341349 50643
rect 341349 50609 341383 50643
rect 341383 50609 341392 50643
rect 341340 50600 341392 50609
rect 2780 50464 2832 50516
rect 4804 50464 4856 50516
rect 367008 48399 367060 48408
rect 367008 48365 367017 48399
rect 367017 48365 367051 48399
rect 367051 48365 367060 48399
rect 367008 48356 367060 48365
rect 230756 48331 230808 48340
rect 230756 48297 230765 48331
rect 230765 48297 230799 48331
rect 230799 48297 230808 48331
rect 230756 48288 230808 48297
rect 244372 48288 244424 48340
rect 244556 48288 244608 48340
rect 278872 48331 278924 48340
rect 278872 48297 278881 48331
rect 278881 48297 278915 48331
rect 278915 48297 278924 48331
rect 278872 48288 278924 48297
rect 281724 48331 281776 48340
rect 281724 48297 281733 48331
rect 281733 48297 281767 48331
rect 281767 48297 281776 48331
rect 281724 48288 281776 48297
rect 284668 48288 284720 48340
rect 284760 48288 284812 48340
rect 288716 48331 288768 48340
rect 288716 48297 288725 48331
rect 288725 48297 288759 48331
rect 288759 48297 288768 48331
rect 288716 48288 288768 48297
rect 291384 48288 291436 48340
rect 291476 48288 291528 48340
rect 295524 48331 295576 48340
rect 295524 48297 295533 48331
rect 295533 48297 295567 48331
rect 295567 48297 295576 48331
rect 295524 48288 295576 48297
rect 299756 48288 299808 48340
rect 301044 48288 301096 48340
rect 325884 48288 325936 48340
rect 326068 48288 326120 48340
rect 327356 48331 327408 48340
rect 327356 48297 327365 48331
rect 327365 48297 327399 48331
rect 327399 48297 327408 48331
rect 327356 48288 327408 48297
rect 337108 48331 337160 48340
rect 337108 48297 337117 48331
rect 337117 48297 337151 48331
rect 337151 48297 337160 48331
rect 337108 48288 337160 48297
rect 357624 48331 357676 48340
rect 357624 48297 357633 48331
rect 357633 48297 357667 48331
rect 357667 48297 357676 48331
rect 357624 48288 357676 48297
rect 389272 48288 389324 48340
rect 460020 48331 460072 48340
rect 460020 48297 460029 48331
rect 460029 48297 460063 48331
rect 460063 48297 460072 48331
rect 460020 48288 460072 48297
rect 236276 48263 236328 48272
rect 236276 48229 236285 48263
rect 236285 48229 236319 48263
rect 236319 48229 236328 48263
rect 236276 48220 236328 48229
rect 299848 48152 299900 48204
rect 323308 48220 323360 48272
rect 323400 48220 323452 48272
rect 301136 48152 301188 48204
rect 460020 48195 460072 48204
rect 460020 48161 460029 48195
rect 460029 48161 460063 48195
rect 460063 48161 460072 48195
rect 460020 48152 460072 48161
rect 250168 46996 250220 47048
rect 327356 46971 327408 46980
rect 327356 46937 327365 46971
rect 327365 46937 327399 46971
rect 327399 46937 327408 46971
rect 327356 46928 327408 46937
rect 250076 46860 250128 46912
rect 265164 46903 265216 46912
rect 265164 46869 265173 46903
rect 265173 46869 265207 46903
rect 265207 46869 265216 46903
rect 265164 46860 265216 46869
rect 266728 46903 266780 46912
rect 266728 46869 266737 46903
rect 266737 46869 266771 46903
rect 266771 46869 266780 46903
rect 266728 46860 266780 46869
rect 284668 46860 284720 46912
rect 286048 46860 286100 46912
rect 286140 46860 286192 46912
rect 291476 46903 291528 46912
rect 291476 46869 291485 46903
rect 291485 46869 291519 46903
rect 291519 46869 291528 46903
rect 291476 46860 291528 46869
rect 323308 46903 323360 46912
rect 323308 46869 323317 46903
rect 323317 46869 323351 46903
rect 323351 46869 323360 46903
rect 323308 46860 323360 46869
rect 339776 46903 339828 46912
rect 339776 46869 339785 46903
rect 339785 46869 339819 46903
rect 339819 46869 339828 46903
rect 339776 46860 339828 46869
rect 367008 46860 367060 46912
rect 375748 46860 375800 46912
rect 375840 46860 375892 46912
rect 377036 46860 377088 46912
rect 377128 46860 377180 46912
rect 247224 45611 247276 45620
rect 247224 45577 247233 45611
rect 247233 45577 247267 45611
rect 247267 45577 247276 45611
rect 247224 45568 247276 45577
rect 259736 45568 259788 45620
rect 393412 45568 393464 45620
rect 393688 45568 393740 45620
rect 251364 45543 251416 45552
rect 251364 45509 251373 45543
rect 251373 45509 251407 45543
rect 251407 45509 251416 45543
rect 251364 45500 251416 45509
rect 299848 45500 299900 45552
rect 310888 45500 310940 45552
rect 311072 45500 311124 45552
rect 317512 45500 317564 45552
rect 317696 45500 317748 45552
rect 245752 44115 245804 44124
rect 245752 44081 245761 44115
rect 245761 44081 245795 44115
rect 245795 44081 245804 44115
rect 245752 44072 245804 44081
rect 303804 42372 303856 42424
rect 304080 42372 304132 42424
rect 339776 42075 339828 42084
rect 339776 42041 339785 42075
rect 339785 42041 339819 42075
rect 339819 42041 339828 42075
rect 339776 42032 339828 42041
rect 460204 41352 460256 41404
rect 306932 40783 306984 40792
rect 306932 40749 306941 40783
rect 306941 40749 306975 40783
rect 306975 40749 306984 40783
rect 306932 40740 306984 40749
rect 245568 40332 245620 40384
rect 245936 40332 245988 40384
rect 437204 40196 437256 40248
rect 437572 40196 437624 40248
rect 456524 40196 456576 40248
rect 456892 40196 456944 40248
rect 417884 40128 417936 40180
rect 418160 40128 418212 40180
rect 230756 38743 230808 38752
rect 230756 38709 230765 38743
rect 230765 38709 230799 38743
rect 230799 38709 230808 38743
rect 230756 38700 230808 38709
rect 244372 38700 244424 38752
rect 267924 38700 267976 38752
rect 325884 38700 325936 38752
rect 366916 38700 366968 38752
rect 236276 38675 236328 38684
rect 236276 38641 236285 38675
rect 236285 38641 236319 38675
rect 236319 38641 236328 38675
rect 236276 38632 236328 38641
rect 244464 38632 244516 38684
rect 270684 38632 270736 38684
rect 270776 38632 270828 38684
rect 272156 38632 272208 38684
rect 272248 38632 272300 38684
rect 324596 38632 324648 38684
rect 324688 38632 324740 38684
rect 327264 38632 327316 38684
rect 327356 38632 327408 38684
rect 329932 38632 329984 38684
rect 330208 38632 330260 38684
rect 331128 38632 331180 38684
rect 331496 38632 331548 38684
rect 267924 38564 267976 38616
rect 281724 38607 281776 38616
rect 281724 38573 281733 38607
rect 281733 38573 281767 38607
rect 281767 38573 281776 38607
rect 281724 38564 281776 38573
rect 325884 38564 325936 38616
rect 366916 38564 366968 38616
rect 372712 38564 372764 38616
rect 372804 38564 372856 38616
rect 460204 38564 460256 38616
rect 232320 37340 232372 37392
rect 230756 37315 230808 37324
rect 230756 37281 230765 37315
rect 230765 37281 230799 37315
rect 230799 37281 230808 37315
rect 230756 37272 230808 37281
rect 232228 37272 232280 37324
rect 265164 37315 265216 37324
rect 265164 37281 265173 37315
rect 265173 37281 265207 37315
rect 265207 37281 265216 37315
rect 265164 37272 265216 37281
rect 266728 37315 266780 37324
rect 266728 37281 266737 37315
rect 266737 37281 266771 37315
rect 266771 37281 266780 37315
rect 266728 37272 266780 37281
rect 284760 37315 284812 37324
rect 284760 37281 284769 37315
rect 284769 37281 284803 37315
rect 284803 37281 284812 37315
rect 323308 37315 323360 37324
rect 284760 37272 284812 37281
rect 323308 37281 323317 37315
rect 323317 37281 323351 37315
rect 323351 37281 323360 37315
rect 323308 37272 323360 37281
rect 366824 37315 366876 37324
rect 366824 37281 366833 37315
rect 366833 37281 366867 37315
rect 366867 37281 366876 37315
rect 366824 37272 366876 37281
rect 389180 37272 389232 37324
rect 389364 37272 389416 37324
rect 270776 37204 270828 37256
rect 270868 37204 270920 37256
rect 288808 37204 288860 37256
rect 288900 37204 288952 37256
rect 393596 37247 393648 37256
rect 393596 37213 393605 37247
rect 393605 37213 393639 37247
rect 393639 37213 393648 37247
rect 393596 37204 393648 37213
rect 232228 37179 232280 37188
rect 232228 37145 232237 37179
rect 232237 37145 232271 37179
rect 232271 37145 232280 37179
rect 232228 37136 232280 37145
rect 259644 37136 259696 37188
rect 259736 37136 259788 37188
rect 249984 35912 250036 35964
rect 250076 35912 250128 35964
rect 251456 35912 251508 35964
rect 291568 35912 291620 35964
rect 299756 35955 299808 35964
rect 299756 35921 299765 35955
rect 299765 35921 299799 35955
rect 299799 35921 299808 35955
rect 299756 35912 299808 35921
rect 306748 35912 306800 35964
rect 3148 35844 3200 35896
rect 6184 35844 6236 35896
rect 247224 35887 247276 35896
rect 247224 35853 247233 35887
rect 247233 35853 247267 35887
rect 247267 35853 247276 35887
rect 247224 35844 247276 35853
rect 259644 35844 259696 35896
rect 270868 35844 270920 35896
rect 294144 35844 294196 35896
rect 294512 35844 294564 35896
rect 250076 35819 250128 35828
rect 250076 35785 250085 35819
rect 250085 35785 250119 35819
rect 250119 35785 250128 35819
rect 250076 35776 250128 35785
rect 245752 34527 245804 34536
rect 245752 34493 245761 34527
rect 245761 34493 245795 34527
rect 245795 34493 245804 34527
rect 245752 34484 245804 34493
rect 317512 31764 317564 31816
rect 317696 31764 317748 31816
rect 339776 31764 339828 31816
rect 341156 31764 341208 31816
rect 377128 31764 377180 31816
rect 460112 31739 460164 31748
rect 460112 31705 460121 31739
rect 460121 31705 460155 31739
rect 460155 31705 460164 31739
rect 460112 31696 460164 31705
rect 341156 31628 341208 31680
rect 377128 31628 377180 31680
rect 306748 31084 306800 31136
rect 253112 29180 253164 29232
rect 257988 29180 258040 29232
rect 366824 29180 366876 29232
rect 437204 29180 437256 29232
rect 437480 29180 437532 29232
rect 465264 29180 465316 29232
rect 467932 29180 467984 29232
rect 367008 29112 367060 29164
rect 417884 29112 417936 29164
rect 418160 29112 418212 29164
rect 357716 29044 357768 29096
rect 492772 29044 492824 29096
rect 502248 29044 502300 29096
rect 262680 28976 262732 29028
rect 262772 28976 262824 29028
rect 265164 28976 265216 29028
rect 265256 28976 265308 29028
rect 267832 28976 267884 29028
rect 267924 28976 267976 29028
rect 281724 29019 281776 29028
rect 281724 28985 281733 29019
rect 281733 28985 281767 29019
rect 281767 28985 281776 29019
rect 281724 28976 281776 28985
rect 301136 28976 301188 29028
rect 301228 28976 301280 29028
rect 339684 29019 339736 29028
rect 339684 28985 339693 29019
rect 339693 28985 339727 29019
rect 339727 28985 339736 29019
rect 339684 28976 339736 28985
rect 357624 28976 357676 29028
rect 375748 28976 375800 29028
rect 375840 28976 375892 29028
rect 284576 28908 284628 28960
rect 284760 28908 284812 28960
rect 306288 28908 306340 28960
rect 314568 28908 314620 28960
rect 323308 28908 323360 28960
rect 323400 28908 323452 28960
rect 324596 28908 324648 28960
rect 324688 28908 324740 28960
rect 325884 28908 325936 28960
rect 325976 28908 326028 28960
rect 295616 27684 295668 27736
rect 389272 27684 389324 27736
rect 389364 27684 389416 27736
rect 232320 27616 232372 27668
rect 291568 27616 291620 27668
rect 291660 27616 291712 27668
rect 295524 27616 295576 27668
rect 393688 27616 393740 27668
rect 230756 27591 230808 27600
rect 230756 27557 230765 27591
rect 230765 27557 230799 27591
rect 230799 27557 230808 27591
rect 230756 27548 230808 27557
rect 265256 27591 265308 27600
rect 265256 27557 265265 27591
rect 265265 27557 265299 27591
rect 265299 27557 265308 27591
rect 265256 27548 265308 27557
rect 302516 27548 302568 27600
rect 302608 27548 302660 27600
rect 367008 27548 367060 27600
rect 375840 27591 375892 27600
rect 375840 27557 375849 27591
rect 375849 27557 375883 27591
rect 375883 27557 375892 27591
rect 375840 27548 375892 27557
rect 247224 26367 247276 26376
rect 247224 26333 247233 26367
rect 247233 26333 247267 26367
rect 247267 26333 247276 26367
rect 247224 26324 247276 26333
rect 259552 26367 259604 26376
rect 259552 26333 259561 26367
rect 259561 26333 259595 26367
rect 259595 26333 259604 26367
rect 259552 26324 259604 26333
rect 306656 26367 306708 26376
rect 306656 26333 306665 26367
rect 306665 26333 306699 26367
rect 306699 26333 306708 26367
rect 306656 26324 306708 26333
rect 250168 26256 250220 26308
rect 270776 26299 270828 26308
rect 270776 26265 270785 26299
rect 270785 26265 270819 26299
rect 270819 26265 270828 26299
rect 270776 26256 270828 26265
rect 303988 26299 304040 26308
rect 303988 26265 303997 26299
rect 303997 26265 304031 26299
rect 304031 26265 304040 26299
rect 303988 26256 304040 26265
rect 329932 26256 329984 26308
rect 330208 26256 330260 26308
rect 245936 26188 245988 26240
rect 247224 26188 247276 26240
rect 259552 26231 259604 26240
rect 259552 26197 259561 26231
rect 259561 26197 259595 26231
rect 259595 26197 259604 26231
rect 259552 26188 259604 26197
rect 272248 26188 272300 26240
rect 291660 26188 291712 26240
rect 310888 26231 310940 26240
rect 310888 26197 310897 26231
rect 310897 26197 310931 26231
rect 310931 26197 310940 26231
rect 310888 26188 310940 26197
rect 331404 26231 331456 26240
rect 331404 26197 331413 26231
rect 331413 26197 331447 26231
rect 331447 26197 331456 26231
rect 331404 26188 331456 26197
rect 389364 26231 389416 26240
rect 389364 26197 389373 26231
rect 389373 26197 389407 26231
rect 389407 26197 389416 26231
rect 389364 26188 389416 26197
rect 329932 25848 329984 25900
rect 303988 24871 304040 24880
rect 303988 24837 303997 24871
rect 303997 24837 304031 24871
rect 304031 24837 304040 24871
rect 303988 24828 304040 24837
rect 232412 22720 232464 22772
rect 267832 22584 267884 22636
rect 244464 22108 244516 22160
rect 250168 22108 250220 22160
rect 269856 22108 269908 22160
rect 270684 22108 270736 22160
rect 377128 22108 377180 22160
rect 377128 21972 377180 22024
rect 460112 21972 460164 22024
rect 460388 21972 460440 22024
rect 375840 20859 375892 20868
rect 375840 20825 375849 20859
rect 375849 20825 375883 20859
rect 375883 20825 375892 20859
rect 375840 20816 375892 20825
rect 251364 19320 251416 19372
rect 251548 19320 251600 19372
rect 266728 19388 266780 19440
rect 281724 19388 281776 19440
rect 281632 19320 281684 19372
rect 339684 19320 339736 19372
rect 339776 19320 339828 19372
rect 341248 19320 341300 19372
rect 341340 19320 341392 19372
rect 266636 19252 266688 19304
rect 295524 19295 295576 19304
rect 295524 19261 295533 19295
rect 295533 19261 295567 19295
rect 295567 19261 295576 19295
rect 295524 19252 295576 19261
rect 339776 19184 339828 19236
rect 230756 18003 230808 18012
rect 230756 17969 230765 18003
rect 230765 17969 230799 18003
rect 230799 17969 230808 18003
rect 230756 17960 230808 17969
rect 259552 17935 259604 17944
rect 259552 17901 259561 17935
rect 259561 17901 259595 17935
rect 259595 17901 259604 17935
rect 259552 17892 259604 17901
rect 264980 17892 265032 17944
rect 393688 18028 393740 18080
rect 273444 17935 273496 17944
rect 273444 17901 273453 17935
rect 273453 17901 273487 17935
rect 273487 17901 273496 17935
rect 273444 17892 273496 17901
rect 393688 17892 393740 17944
rect 299388 16940 299440 16992
rect 311164 16940 311216 16992
rect 417884 16736 417936 16788
rect 418160 16736 418212 16788
rect 437204 16736 437256 16788
rect 437480 16736 437532 16788
rect 463792 16668 463844 16720
rect 466552 16668 466604 16720
rect 244188 16643 244240 16652
rect 244188 16609 244197 16643
rect 244197 16609 244231 16643
rect 244231 16609 244240 16643
rect 244188 16600 244240 16609
rect 245844 16643 245896 16652
rect 245844 16609 245853 16643
rect 245853 16609 245887 16643
rect 245887 16609 245896 16643
rect 245844 16600 245896 16609
rect 249984 16643 250036 16652
rect 249984 16609 249993 16643
rect 249993 16609 250027 16643
rect 250027 16609 250036 16643
rect 249984 16600 250036 16609
rect 291568 16643 291620 16652
rect 291568 16609 291577 16643
rect 291577 16609 291611 16643
rect 291611 16609 291620 16643
rect 291568 16600 291620 16609
rect 310888 16643 310940 16652
rect 310888 16609 310897 16643
rect 310897 16609 310931 16643
rect 310931 16609 310940 16643
rect 310888 16600 310940 16609
rect 389364 16643 389416 16652
rect 389364 16609 389373 16643
rect 389373 16609 389407 16643
rect 389407 16609 389416 16643
rect 389364 16600 389416 16609
rect 306840 15172 306892 15224
rect 307024 15172 307076 15224
rect 110328 15104 110380 15156
rect 274732 15104 274784 15156
rect 107476 15036 107528 15088
rect 273352 15036 273404 15088
rect 103428 14968 103480 15020
rect 271972 14968 272024 15020
rect 99288 14900 99340 14952
rect 270592 14900 270644 14952
rect 96528 14832 96580 14884
rect 269212 14832 269264 14884
rect 92388 14764 92440 14816
rect 266452 14764 266504 14816
rect 89628 14696 89680 14748
rect 265072 14696 265124 14748
rect 85488 14628 85540 14680
rect 263692 14628 263744 14680
rect 82728 14560 82780 14612
rect 262588 14560 262640 14612
rect 78588 14492 78640 14544
rect 260932 14492 260984 14544
rect 74448 14424 74500 14476
rect 259552 14424 259604 14476
rect 114468 14356 114520 14408
rect 276112 14356 276164 14408
rect 117228 14288 117280 14340
rect 277676 14288 277728 14340
rect 121368 14220 121420 14272
rect 278780 14220 278832 14272
rect 125416 14152 125468 14204
rect 280252 14152 280304 14204
rect 232136 14127 232188 14136
rect 232136 14093 232145 14127
rect 232145 14093 232179 14127
rect 232179 14093 232188 14127
rect 232136 14084 232188 14093
rect 183468 13744 183520 13796
rect 303988 13744 304040 13796
rect 186228 13676 186280 13728
rect 306564 13676 306616 13728
rect 179328 13608 179380 13660
rect 302516 13608 302568 13660
rect 176568 13540 176620 13592
rect 301044 13540 301096 13592
rect 172428 13472 172480 13524
rect 299756 13472 299808 13524
rect 168288 13404 168340 13456
rect 298284 13404 298336 13456
rect 165528 13336 165580 13388
rect 296904 13336 296956 13388
rect 160008 13268 160060 13320
rect 294420 13268 294472 13320
rect 155868 13200 155920 13252
rect 292764 13200 292816 13252
rect 71688 13132 71740 13184
rect 258172 13132 258224 13184
rect 31668 13064 31720 13116
rect 241612 13064 241664 13116
rect 190368 12996 190420 13048
rect 307944 12996 307996 13048
rect 206928 12928 206980 12980
rect 314844 12928 314896 12980
rect 211068 12860 211120 12912
rect 316224 12860 316276 12912
rect 213828 12792 213880 12844
rect 317604 12792 317656 12844
rect 217968 12724 218020 12776
rect 318984 12724 319036 12776
rect 220728 12656 220780 12708
rect 320272 12656 320324 12708
rect 224868 12588 224920 12640
rect 321744 12588 321796 12640
rect 229008 12520 229060 12572
rect 323124 12520 323176 12572
rect 230756 12452 230808 12504
rect 366916 12452 366968 12504
rect 173808 12384 173860 12436
rect 300952 12384 301004 12436
rect 169668 12316 169720 12368
rect 299572 12316 299624 12368
rect 366916 12316 366968 12368
rect 166908 12248 166960 12300
rect 298192 12248 298244 12300
rect 162768 12180 162820 12232
rect 151728 12112 151780 12164
rect 291568 12112 291620 12164
rect 148968 12044 149020 12096
rect 290004 12044 290056 12096
rect 144828 11976 144880 12028
rect 288900 11976 288952 12028
rect 142068 11908 142120 11960
rect 287336 11908 287388 11960
rect 128268 11840 128320 11892
rect 281632 11840 281684 11892
rect 126888 11772 126940 11824
rect 281540 11772 281592 11824
rect 23388 11704 23440 11756
rect 238944 11704 238996 11756
rect 468852 11704 468904 11756
rect 469128 11704 469180 11756
rect 176476 11636 176528 11688
rect 302332 11636 302384 11688
rect 180708 11568 180760 11620
rect 303712 11568 303764 11620
rect 184848 11500 184900 11552
rect 305092 11500 305144 11552
rect 187608 11432 187660 11484
rect 306472 11432 306524 11484
rect 191748 11364 191800 11416
rect 308036 11364 308088 11416
rect 194508 11296 194560 11348
rect 309416 11296 309468 11348
rect 198648 11228 198700 11280
rect 310888 11228 310940 11280
rect 230664 11203 230716 11212
rect 230664 11169 230673 11203
rect 230673 11169 230707 11203
rect 230707 11169 230716 11203
rect 230664 11160 230716 11169
rect 113088 10956 113140 11008
rect 276020 10956 276072 11008
rect 108948 10888 109000 10940
rect 106188 10820 106240 10872
rect 102048 10752 102100 10804
rect 269856 10752 269908 10804
rect 99196 10684 99248 10736
rect 269304 10684 269356 10736
rect 95148 10616 95200 10668
rect 91008 10548 91060 10600
rect 266636 10548 266688 10600
rect 64788 10480 64840 10532
rect 255596 10480 255648 10532
rect 60648 10412 60700 10464
rect 254032 10412 254084 10464
rect 56508 10344 56560 10396
rect 252652 10344 252704 10396
rect 53748 10276 53800 10328
rect 251272 10276 251324 10328
rect 117136 10208 117188 10260
rect 277584 10208 277636 10260
rect 119988 10140 120040 10192
rect 278964 10140 279016 10192
rect 124128 10072 124180 10124
rect 280344 10072 280396 10124
rect 143448 10004 143500 10056
rect 288532 10004 288584 10056
rect 147588 9936 147640 9988
rect 289820 9936 289872 9988
rect 151636 9868 151688 9920
rect 291292 9868 291344 9920
rect 154488 9800 154540 9852
rect 292856 9800 292908 9852
rect 158628 9732 158680 9784
rect 294052 9732 294104 9784
rect 161388 9664 161440 9716
rect 295432 9664 295484 9716
rect 330208 9707 330260 9716
rect 330208 9673 330217 9707
rect 330217 9673 330251 9707
rect 330251 9673 330260 9707
rect 330208 9664 330260 9673
rect 331404 9707 331456 9716
rect 331404 9673 331413 9707
rect 331413 9673 331447 9707
rect 331447 9673 331456 9707
rect 331404 9664 331456 9673
rect 339684 9707 339736 9716
rect 339684 9673 339693 9707
rect 339693 9673 339727 9707
rect 339727 9673 339736 9707
rect 339684 9664 339736 9673
rect 366824 9707 366876 9716
rect 366824 9673 366833 9707
rect 366833 9673 366867 9707
rect 366867 9673 366876 9707
rect 366824 9664 366876 9673
rect 203892 9596 203944 9648
rect 313372 9596 313424 9648
rect 200396 9528 200448 9580
rect 311992 9528 312044 9580
rect 196808 9460 196860 9512
rect 310612 9460 310664 9512
rect 193220 9392 193272 9444
rect 309232 9392 309284 9444
rect 139676 9324 139728 9376
rect 287152 9324 287204 9376
rect 136088 9256 136140 9308
rect 285864 9256 285916 9308
rect 49332 9188 49384 9240
rect 249892 9188 249944 9240
rect 253848 9188 253900 9240
rect 334164 9188 334216 9240
rect 44548 9120 44600 9172
rect 250352 9120 250404 9172
rect 332784 9120 332836 9172
rect 27896 9052 27948 9104
rect 233884 9052 233936 9104
rect 243176 9052 243228 9104
rect 330024 9052 330076 9104
rect 18328 8984 18380 9036
rect 236184 8984 236236 9036
rect 239588 8984 239640 9036
rect 328644 8984 328696 9036
rect 13636 8916 13688 8968
rect 234804 8916 234856 8968
rect 236000 8916 236052 8968
rect 325976 8916 326028 8968
rect 207480 8848 207532 8900
rect 314936 8848 314988 8900
rect 210976 8780 211028 8832
rect 316132 8780 316184 8832
rect 214656 8712 214708 8764
rect 317512 8712 317564 8764
rect 218152 8644 218204 8696
rect 318892 8644 318944 8696
rect 221740 8576 221792 8628
rect 320180 8576 320232 8628
rect 225328 8508 225380 8560
rect 321652 8508 321704 8560
rect 228916 8440 228968 8492
rect 323308 8440 323360 8492
rect 232504 8372 232556 8424
rect 324596 8372 324648 8424
rect 246764 8304 246816 8356
rect 331404 8304 331456 8356
rect 87328 8236 87380 8288
rect 265164 8236 265216 8288
rect 270500 8236 270552 8288
rect 340972 8236 341024 8288
rect 445484 8236 445536 8288
rect 523868 8236 523920 8288
rect 83832 8168 83884 8220
rect 263876 8168 263928 8220
rect 267004 8168 267056 8220
rect 339592 8168 339644 8220
rect 446956 8168 447008 8220
rect 527456 8168 527508 8220
rect 80244 8100 80296 8152
rect 262404 8100 262456 8152
rect 263416 8100 263468 8152
rect 338304 8100 338356 8152
rect 448244 8100 448296 8152
rect 531044 8100 531096 8152
rect 40960 8032 41012 8084
rect 245936 8032 245988 8084
rect 259828 8032 259880 8084
rect 336924 8032 336976 8084
rect 451004 8032 451056 8084
rect 534540 8032 534592 8084
rect 37372 7964 37424 8016
rect 244280 7964 244332 8016
rect 256240 7964 256292 8016
rect 334072 7964 334124 8016
rect 452476 7964 452528 8016
rect 538128 7964 538180 8016
rect 33876 7896 33928 7948
rect 242992 7896 243044 7948
rect 252652 7896 252704 7948
rect 332692 7896 332744 7948
rect 453764 7896 453816 7948
rect 541716 7896 541768 7948
rect 30288 7828 30340 7880
rect 241796 7828 241848 7880
rect 249156 7828 249208 7880
rect 331312 7828 331364 7880
rect 455236 7828 455288 7880
rect 545304 7828 545356 7880
rect 26700 7760 26752 7812
rect 240416 7760 240468 7812
rect 245568 7760 245620 7812
rect 330208 7760 330260 7812
rect 456616 7760 456668 7812
rect 548892 7760 548944 7812
rect 21916 7692 21968 7744
rect 238852 7692 238904 7744
rect 241980 7692 242032 7744
rect 328552 7692 328604 7744
rect 457996 7692 458048 7744
rect 552388 7692 552440 7744
rect 8852 7624 8904 7676
rect 4068 7556 4120 7608
rect 230664 7624 230716 7676
rect 234804 7624 234856 7676
rect 325792 7624 325844 7676
rect 459376 7624 459428 7676
rect 555976 7624 556028 7676
rect 227720 7556 227772 7608
rect 229008 7556 229060 7608
rect 231308 7556 231360 7608
rect 324412 7556 324464 7608
rect 460756 7556 460808 7608
rect 559564 7556 559616 7608
rect 134892 7488 134944 7540
rect 284576 7488 284628 7540
rect 444196 7488 444248 7540
rect 520280 7488 520332 7540
rect 138480 7420 138532 7472
rect 285956 7420 286008 7472
rect 442816 7420 442868 7472
rect 516784 7420 516836 7472
rect 141976 7352 142028 7404
rect 287060 7352 287112 7404
rect 441436 7352 441488 7404
rect 513196 7352 513248 7404
rect 145656 7284 145708 7336
rect 288440 7284 288492 7336
rect 440056 7284 440108 7336
rect 509608 7284 509660 7336
rect 149244 7216 149296 7268
rect 291200 7216 291252 7268
rect 152740 7148 152792 7200
rect 292580 7148 292632 7200
rect 156328 7080 156380 7132
rect 293960 7080 294012 7132
rect 159916 7012 159968 7064
rect 295340 7012 295392 7064
rect 233424 6944 233476 6996
rect 238392 6944 238444 6996
rect 327264 6944 327316 6996
rect 306656 6876 306708 6928
rect 306840 6876 306892 6928
rect 389364 6876 389416 6928
rect 389548 6876 389600 6928
rect 393688 6876 393740 6928
rect 394148 6876 394200 6928
rect 516692 6876 516744 6928
rect 516876 6876 516928 6928
rect 170588 6808 170640 6860
rect 299480 6808 299532 6860
rect 431868 6808 431920 6860
rect 490564 6808 490616 6860
rect 167092 6740 167144 6792
rect 298376 6740 298428 6792
rect 433156 6740 433208 6792
rect 491760 6740 491812 6792
rect 163504 6672 163556 6724
rect 296720 6672 296772 6724
rect 297364 6672 297416 6724
rect 336832 6672 336884 6724
rect 434628 6672 434680 6724
rect 495348 6672 495400 6724
rect 131396 6604 131448 6656
rect 283012 6604 283064 6656
rect 295892 6604 295944 6656
rect 335452 6604 335504 6656
rect 433248 6604 433300 6656
rect 494152 6604 494204 6656
rect 76656 6536 76708 6588
rect 261024 6536 261076 6588
rect 298100 6536 298152 6588
rect 338396 6536 338448 6588
rect 435916 6536 435968 6588
rect 497740 6536 497792 6588
rect 73068 6468 73120 6520
rect 259460 6468 259512 6520
rect 289820 6468 289872 6520
rect 339684 6468 339736 6520
rect 436008 6468 436060 6520
rect 498936 6468 498988 6520
rect 69480 6400 69532 6452
rect 258264 6400 258316 6452
rect 288440 6400 288492 6452
rect 341248 6400 341300 6452
rect 437388 6400 437440 6452
rect 501236 6400 501288 6452
rect 65984 6332 66036 6384
rect 256792 6332 256844 6384
rect 288532 6332 288584 6384
rect 343640 6332 343692 6384
rect 437296 6332 437348 6384
rect 502432 6332 502484 6384
rect 62396 6264 62448 6316
rect 255504 6264 255556 6316
rect 294328 6264 294380 6316
rect 350632 6264 350684 6316
rect 438676 6264 438728 6316
rect 504824 6264 504876 6316
rect 58808 6196 58860 6248
rect 253940 6196 253992 6248
rect 280068 6196 280120 6248
rect 345204 6196 345256 6248
rect 438768 6196 438820 6248
rect 506020 6196 506072 6248
rect 55220 6128 55272 6180
rect 251456 6128 251508 6180
rect 274088 6128 274140 6180
rect 342352 6128 342404 6180
rect 440148 6128 440200 6180
rect 508412 6128 508464 6180
rect 174176 6060 174228 6112
rect 300860 6060 300912 6112
rect 431776 6060 431828 6112
rect 488172 6060 488224 6112
rect 177764 5992 177816 6044
rect 302240 5992 302292 6044
rect 430488 5992 430540 6044
rect 486976 5992 487028 6044
rect 181352 5924 181404 5976
rect 303620 5924 303672 5976
rect 430396 5924 430448 5976
rect 484584 5924 484636 5976
rect 184848 5856 184900 5908
rect 305000 5856 305052 5908
rect 429108 5856 429160 5908
rect 483480 5856 483532 5908
rect 188436 5788 188488 5840
rect 306656 5788 306708 5840
rect 427728 5788 427780 5840
rect 479892 5788 479944 5840
rect 192024 5720 192076 5772
rect 307760 5720 307812 5772
rect 426348 5720 426400 5772
rect 476304 5720 476356 5772
rect 195612 5652 195664 5704
rect 309140 5652 309192 5704
rect 202696 5584 202748 5636
rect 313280 5584 313332 5636
rect 199200 5516 199252 5568
rect 310520 5516 310572 5568
rect 137284 5448 137336 5500
rect 285680 5448 285732 5500
rect 297824 5448 297876 5500
rect 352104 5448 352156 5500
rect 452568 5448 452620 5500
rect 540520 5448 540572 5500
rect 133788 5380 133840 5432
rect 284300 5380 284352 5432
rect 290740 5380 290792 5432
rect 349344 5380 349396 5432
rect 408408 5380 408460 5432
rect 433524 5380 433576 5432
rect 453856 5380 453908 5432
rect 544108 5380 544160 5432
rect 130200 5312 130252 5364
rect 283196 5312 283248 5364
rect 287152 5312 287204 5364
rect 347964 5312 348016 5364
rect 412456 5312 412508 5364
rect 440608 5312 440660 5364
rect 455328 5312 455380 5364
rect 547696 5312 547748 5364
rect 67180 5244 67232 5296
rect 256976 5244 257028 5296
rect 283656 5244 283708 5296
rect 346584 5244 346636 5296
rect 413836 5244 413888 5296
rect 444196 5244 444248 5296
rect 459468 5244 459520 5296
rect 48136 5176 48188 5228
rect 248512 5176 248564 5228
rect 251456 5176 251508 5228
rect 332600 5176 332652 5228
rect 415308 5176 415360 5228
rect 447784 5176 447836 5228
rect 460848 5176 460900 5228
rect 551192 5244 551244 5296
rect 17224 5108 17276 5160
rect 236092 5108 236144 5160
rect 247960 5108 248012 5160
rect 331220 5108 331272 5160
rect 416596 5108 416648 5160
rect 451280 5108 451332 5160
rect 12440 5040 12492 5092
rect 234712 5040 234764 5092
rect 244372 5040 244424 5092
rect 321652 5040 321704 5092
rect 327080 5040 327132 5092
rect 329840 5040 329892 5092
rect 337108 5040 337160 5092
rect 368572 5040 368624 5092
rect 417976 5040 418028 5092
rect 454868 5040 454920 5092
rect 7656 4972 7708 5024
rect 232136 4972 232188 5024
rect 240784 4972 240836 5024
rect 328736 4972 328788 5024
rect 333612 4972 333664 5024
rect 367192 4972 367244 5024
rect 380164 4972 380216 5024
rect 419448 4972 419500 5024
rect 458456 4972 458508 5024
rect 463516 5108 463568 5160
rect 554780 5176 554832 5228
rect 464988 5040 465040 5092
rect 558368 5108 558420 5160
rect 465632 4972 465684 5024
rect 561956 5040 562008 5092
rect 2872 4904 2924 4956
rect 572 4836 624 4888
rect 229100 4904 229152 4956
rect 237196 4904 237248 4956
rect 321652 4904 321704 4956
rect 327080 4904 327132 4956
rect 361672 4904 361724 4956
rect 381544 4904 381596 4956
rect 420736 4904 420788 4956
rect 458088 4904 458140 4956
rect 466184 4904 466236 4956
rect 565544 4972 565596 5024
rect 230112 4836 230164 4888
rect 324320 4836 324372 4888
rect 326344 4836 326396 4888
rect 360384 4836 360436 4888
rect 422208 4836 422260 4888
rect 1676 4768 1728 4820
rect 230572 4768 230624 4820
rect 233700 4768 233752 4820
rect 325700 4768 325752 4820
rect 328460 4768 328512 4820
rect 363052 4768 363104 4820
rect 423588 4768 423640 4820
rect 469128 4836 469180 4888
rect 569040 4904 569092 4956
rect 572628 4836 572680 4888
rect 462136 4768 462188 4820
rect 468944 4768 468996 4820
rect 579804 4768 579856 4820
rect 212264 4700 212316 4752
rect 316040 4700 316092 4752
rect 318708 4700 318760 4752
rect 215852 4632 215904 4684
rect 317420 4632 317472 4684
rect 323308 4700 323360 4752
rect 359004 4700 359056 4752
rect 451096 4700 451148 4752
rect 536932 4700 536984 4752
rect 333980 4632 334032 4684
rect 365720 4632 365772 4684
rect 366916 4632 366968 4684
rect 449808 4632 449860 4684
rect 533436 4632 533488 4684
rect 219348 4564 219400 4616
rect 318800 4564 318852 4616
rect 222936 4496 222988 4548
rect 321376 4564 321428 4616
rect 322756 4564 322808 4616
rect 337200 4564 337252 4616
rect 448336 4564 448388 4616
rect 529848 4564 529900 4616
rect 320364 4496 320416 4548
rect 335360 4496 335412 4548
rect 353484 4496 353536 4548
rect 447048 4496 447100 4548
rect 526260 4496 526312 4548
rect 226524 4428 226576 4480
rect 322940 4428 322992 4480
rect 325148 4428 325200 4480
rect 338120 4428 338172 4480
rect 352564 4428 352616 4480
rect 445576 4428 445628 4480
rect 522672 4428 522724 4480
rect 201500 4360 201552 4412
rect 271144 4360 271196 4412
rect 301412 4360 301464 4412
rect 444288 4360 444340 4412
rect 519084 4360 519136 4412
rect 205088 4292 205140 4344
rect 272524 4292 272576 4344
rect 305000 4292 305052 4344
rect 354956 4292 355008 4344
rect 442908 4292 442960 4344
rect 515588 4292 515640 4344
rect 230480 4224 230532 4276
rect 308588 4224 308640 4276
rect 356152 4224 356204 4276
rect 441528 4224 441580 4276
rect 512000 4224 512052 4276
rect 124220 4156 124272 4208
rect 125416 4156 125468 4208
rect 140872 4156 140924 4208
rect 142068 4156 142120 4208
rect 150440 4156 150492 4208
rect 151636 4156 151688 4208
rect 158720 4156 158772 4208
rect 160008 4156 160060 4208
rect 175372 4156 175424 4208
rect 176568 4156 176620 4208
rect 209872 4156 209924 4208
rect 211068 4156 211120 4208
rect 57612 4088 57664 4140
rect 250444 4088 250496 4140
rect 268108 4088 268160 4140
rect 269028 4088 269080 4140
rect 284760 4088 284812 4140
rect 285588 4088 285640 4140
rect 312176 4156 312228 4208
rect 357532 4156 357584 4208
rect 424968 4156 425020 4208
rect 472716 4156 472768 4208
rect 50528 4020 50580 4072
rect 249064 4020 249116 4072
rect 295892 4088 295944 4140
rect 296720 4088 296772 4140
rect 297916 4088 297968 4140
rect 300308 4088 300360 4140
rect 332416 4088 332468 4140
rect 333244 4088 333296 4140
rect 334716 4088 334768 4140
rect 335268 4088 335320 4140
rect 338764 4088 338816 4140
rect 339500 4088 339552 4140
rect 340788 4088 340840 4140
rect 345664 4088 345716 4140
rect 347872 4088 347924 4140
rect 349068 4088 349120 4140
rect 351184 4088 351236 4140
rect 351368 4088 351420 4140
rect 351828 4088 351880 4140
rect 358912 4088 358964 4140
rect 362132 4088 362184 4140
rect 362868 4088 362920 4140
rect 363328 4088 363380 4140
rect 364248 4088 364300 4140
rect 369216 4088 369268 4140
rect 369768 4088 369820 4140
rect 370412 4088 370464 4140
rect 371148 4088 371200 4140
rect 377588 4088 377640 4140
rect 378048 4088 378100 4140
rect 378784 4088 378836 4140
rect 385316 4088 385368 4140
rect 390836 4088 390888 4140
rect 391848 4088 391900 4140
rect 393228 4088 393280 4140
rect 395436 4088 395488 4140
rect 398104 4088 398156 4140
rect 403716 4088 403768 4140
rect 409696 4088 409748 4140
rect 437020 4088 437072 4140
rect 445668 4088 445720 4140
rect 521476 4088 521528 4140
rect 529204 4088 529256 4140
rect 575020 4088 575072 4140
rect 298100 4020 298152 4072
rect 302608 4020 302660 4072
rect 309784 4020 309836 4072
rect 314568 4020 314620 4072
rect 46940 3952 46992 4004
rect 248696 3952 248748 4004
rect 257436 3952 257488 4004
rect 297364 3952 297416 4004
rect 313372 3952 313424 4004
rect 374000 4020 374052 4072
rect 383568 4020 383620 4072
rect 384304 4020 384356 4072
rect 393136 4020 393188 4072
rect 396632 4020 396684 4072
rect 411076 4020 411128 4072
rect 439412 4020 439464 4072
rect 442264 4020 442316 4072
rect 355324 3952 355376 4004
rect 359096 3952 359148 4004
rect 359740 3952 359792 4004
rect 377128 3952 377180 4004
rect 406384 3952 406436 4004
rect 414480 3952 414532 4004
rect 420184 3952 420236 4004
rect 423956 3952 424008 4004
rect 424416 3952 424468 4004
rect 446588 3952 446640 4004
rect 448428 4020 448480 4072
rect 528652 4020 528704 4072
rect 530584 4020 530636 4072
rect 582196 4020 582248 4072
rect 451188 3952 451240 4004
rect 535736 3952 535788 4004
rect 45744 3884 45796 3936
rect 247684 3884 247736 3936
rect 282460 3884 282512 3936
rect 39764 3816 39816 3868
rect 238116 3816 238168 3868
rect 264612 3816 264664 3868
rect 20720 3748 20772 3800
rect 35164 3748 35216 3800
rect 38568 3748 38620 3800
rect 245660 3748 245712 3800
rect 278872 3748 278924 3800
rect 289544 3816 289596 3868
rect 365812 3884 365864 3936
rect 371608 3884 371660 3936
rect 405004 3884 405056 3936
rect 416872 3884 416924 3936
rect 420276 3884 420328 3936
rect 450176 3884 450228 3936
rect 453948 3884 454000 3936
rect 542912 3884 542964 3936
rect 285956 3748 286008 3800
rect 335544 3748 335596 3800
rect 342904 3816 342956 3868
rect 343088 3816 343140 3868
rect 369124 3816 369176 3868
rect 372804 3816 372856 3868
rect 373908 3816 373960 3868
rect 399484 3816 399536 3868
rect 407304 3816 407356 3868
rect 412548 3816 412600 3868
rect 443000 3816 443052 3868
rect 341524 3748 341576 3800
rect 341892 3748 341944 3800
rect 370136 3748 370188 3800
rect 374000 3748 374052 3800
rect 375288 3748 375340 3800
rect 399576 3748 399628 3800
rect 408500 3748 408552 3800
rect 413284 3748 413336 3800
rect 413468 3748 413520 3800
rect 413928 3748 413980 3800
rect 445392 3748 445444 3800
rect 32680 3680 32732 3732
rect 243084 3680 243136 3732
rect 326436 3680 326488 3732
rect 328460 3680 328512 3732
rect 331220 3680 331272 3732
rect 338304 3680 338356 3732
rect 368664 3680 368716 3732
rect 375196 3680 375248 3732
rect 383844 3680 383896 3732
rect 402796 3680 402848 3732
rect 419172 3680 419224 3732
rect 421564 3680 421616 3732
rect 24308 3612 24360 3664
rect 239036 3612 239088 3664
rect 262220 3612 262272 3664
rect 11244 3544 11296 3596
rect 19984 3544 20036 3596
rect 25504 3544 25556 3596
rect 240324 3544 240376 3596
rect 265808 3544 265860 3596
rect 325148 3612 325200 3664
rect 325240 3612 325292 3664
rect 322848 3544 322900 3596
rect 327080 3544 327132 3596
rect 358084 3612 358136 3664
rect 360936 3612 360988 3664
rect 377404 3612 377456 3664
rect 400128 3612 400180 3664
rect 412088 3612 412140 3664
rect 417424 3612 417476 3664
rect 427084 3612 427136 3664
rect 431132 3612 431184 3664
rect 453672 3816 453724 3868
rect 550088 3816 550140 3868
rect 460388 3748 460440 3800
rect 463240 3748 463292 3800
rect 452476 3680 452528 3732
rect 456708 3680 456760 3732
rect 460296 3680 460348 3732
rect 449164 3612 449216 3664
rect 557172 3748 557224 3800
rect 14832 3476 14884 3528
rect 234896 3476 234948 3528
rect 258632 3476 258684 3528
rect 320364 3476 320416 3528
rect 320456 3476 320508 3528
rect 321192 3476 321244 3528
rect 321652 3476 321704 3528
rect 361856 3544 361908 3596
rect 382372 3544 382424 3596
rect 386604 3544 386656 3596
rect 402888 3544 402940 3596
rect 420368 3544 420420 3596
rect 420828 3544 420880 3596
rect 460848 3544 460900 3596
rect 462228 3544 462280 3596
rect 564348 3680 564400 3732
rect 463608 3612 463660 3664
rect 566740 3612 566792 3664
rect 466368 3544 466420 3596
rect 571432 3544 571484 3596
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 16028 3408 16080 3460
rect 236276 3408 236328 3460
rect 255044 3408 255096 3460
rect 318708 3408 318760 3460
rect 322756 3408 322808 3460
rect 324044 3408 324096 3460
rect 363144 3476 363196 3528
rect 363604 3408 363656 3460
rect 368020 3408 368072 3460
rect 379980 3476 380032 3528
rect 380808 3476 380860 3528
rect 381176 3476 381228 3528
rect 382188 3476 382240 3528
rect 388260 3476 388312 3528
rect 389088 3476 389140 3528
rect 389272 3476 389324 3528
rect 394608 3476 394660 3528
rect 399024 3476 399076 3528
rect 402244 3476 402296 3528
rect 415676 3476 415728 3528
rect 418068 3476 418120 3528
rect 457260 3476 457312 3528
rect 466276 3476 466328 3528
rect 573824 3476 573876 3528
rect 379704 3408 379756 3460
rect 404268 3408 404320 3460
rect 422760 3408 422812 3460
rect 424324 3408 424376 3460
rect 425152 3408 425204 3460
rect 467932 3408 467984 3460
rect 469036 3408 469088 3460
rect 578608 3408 578660 3460
rect 19524 3340 19576 3392
rect 28264 3340 28316 3392
rect 29092 3340 29144 3392
rect 32404 3340 32456 3392
rect 34980 3340 35032 3392
rect 57244 3340 57296 3392
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 64696 3340 64748 3392
rect 251824 3340 251876 3392
rect 289820 3340 289872 3392
rect 299112 3340 299164 3392
rect 302884 3340 302936 3392
rect 310980 3340 311032 3392
rect 353760 3340 353812 3392
rect 375656 3340 375708 3392
rect 409788 3340 409840 3392
rect 10048 3272 10100 3324
rect 13084 3272 13136 3324
rect 42156 3272 42208 3324
rect 66904 3272 66956 3324
rect 70676 3272 70728 3324
rect 71688 3272 71740 3324
rect 71872 3272 71924 3324
rect 253204 3272 253256 3324
rect 43352 3204 43404 3256
rect 61384 3204 61436 3256
rect 63592 3204 63644 3256
rect 64788 3204 64840 3256
rect 77852 3204 77904 3256
rect 78588 3204 78640 3256
rect 81440 3204 81492 3256
rect 82728 3204 82780 3256
rect 84844 3204 84896 3256
rect 84936 3204 84988 3256
rect 85488 3204 85540 3256
rect 88524 3204 88576 3256
rect 89628 3204 89680 3256
rect 52828 3136 52880 3188
rect 53748 3136 53800 3188
rect 54024 3136 54076 3188
rect 71044 3136 71096 3188
rect 79048 3136 79100 3188
rect 254584 3204 254636 3256
rect 269304 3204 269356 3256
rect 61200 3068 61252 3120
rect 77944 3068 77996 3120
rect 82636 3068 82688 3120
rect 36176 3000 36228 3052
rect 39304 3000 39356 3052
rect 68284 3000 68336 3052
rect 75460 3000 75512 3052
rect 79324 2864 79376 2916
rect 89720 3068 89772 3120
rect 255964 3136 256016 3188
rect 272892 3136 272944 3188
rect 288440 3272 288492 3324
rect 303804 3272 303856 3324
rect 344376 3272 344428 3324
rect 345756 3272 345808 3324
rect 348424 3272 348476 3324
rect 349068 3272 349120 3324
rect 365536 3272 365588 3324
rect 394516 3272 394568 3324
rect 400220 3272 400272 3324
rect 403624 3272 403676 3324
rect 410892 3272 410944 3324
rect 411168 3340 411220 3392
rect 438216 3340 438268 3392
rect 443644 3340 443696 3392
rect 276480 3204 276532 3256
rect 288532 3204 288584 3256
rect 291936 3204 291988 3256
rect 316684 3204 316736 3256
rect 318064 3204 318116 3256
rect 350264 3204 350316 3256
rect 352564 3204 352616 3256
rect 357348 3204 357400 3256
rect 376024 3204 376076 3256
rect 407028 3204 407080 3256
rect 277676 3136 277728 3188
rect 290464 3136 290516 3188
rect 309784 3136 309836 3188
rect 335912 3136 335964 3188
rect 340696 3136 340748 3188
rect 346676 3136 346728 3188
rect 370504 3136 370556 3188
rect 405648 3136 405700 3188
rect 426348 3136 426400 3188
rect 428464 3272 428516 3324
rect 434076 3272 434128 3324
rect 441804 3272 441856 3324
rect 442356 3272 442408 3324
rect 503628 3272 503680 3324
rect 514024 3340 514076 3392
rect 517888 3340 517940 3392
rect 514392 3272 514444 3324
rect 516876 3272 516928 3324
rect 525064 3340 525116 3392
rect 527824 3340 527876 3392
rect 567844 3340 567896 3392
rect 429936 3204 429988 3256
rect 430120 3204 430172 3256
rect 433984 3204 434036 3256
rect 434628 3136 434680 3188
rect 439504 3204 439556 3256
rect 496544 3204 496596 3256
rect 512644 3204 512696 3256
rect 577412 3272 577464 3324
rect 570236 3204 570288 3256
rect 489368 3136 489420 3188
rect 505744 3136 505796 3188
rect 563152 3136 563204 3188
rect 94504 3068 94556 3120
rect 95148 3068 95200 3120
rect 95700 3068 95752 3120
rect 96528 3068 96580 3120
rect 98092 3068 98144 3120
rect 99196 3068 99248 3120
rect 101588 3068 101640 3120
rect 102048 3068 102100 3120
rect 102784 3068 102836 3120
rect 103428 3068 103480 3120
rect 105176 3068 105228 3120
rect 106188 3068 106240 3120
rect 106372 3068 106424 3120
rect 107476 3068 107528 3120
rect 86132 3000 86184 3052
rect 93308 2932 93360 2984
rect 97264 3000 97316 3052
rect 95884 2796 95936 2848
rect 96896 2932 96948 2984
rect 257344 3068 257396 3120
rect 295524 3068 295576 3120
rect 319444 3068 319496 3120
rect 327724 3068 327776 3120
rect 328828 3068 328880 3120
rect 359464 3068 359516 3120
rect 372988 3068 373040 3120
rect 398196 3068 398248 3120
rect 103980 2864 104032 2916
rect 258816 3000 258868 3052
rect 293132 3000 293184 3052
rect 312544 3000 312596 3052
rect 315764 3000 315816 3052
rect 323308 3000 323360 3052
rect 327632 3000 327684 3052
rect 335912 3000 335964 3052
rect 112352 2932 112404 2984
rect 113088 2932 113140 2984
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 115940 2932 115992 2984
rect 116952 2932 117004 2984
rect 119436 2932 119488 2984
rect 119988 2932 120040 2984
rect 120632 2932 120684 2984
rect 121368 2932 121420 2984
rect 111156 2864 111208 2916
rect 258724 2932 258776 2984
rect 316960 2932 317012 2984
rect 344376 2932 344428 2984
rect 345480 2932 345532 2984
rect 102600 2796 102652 2848
rect 114744 2796 114796 2848
rect 260104 2864 260156 2916
rect 275284 2864 275336 2916
rect 275928 2864 275980 2916
rect 319260 2864 319312 2916
rect 326344 2864 326396 2916
rect 340880 2864 340932 2916
rect 344284 2864 344336 2916
rect 354956 2932 355008 2984
rect 355968 2932 356020 2984
rect 364524 3000 364576 3052
rect 365536 3000 365588 3052
rect 376392 3000 376444 3052
rect 381636 3000 381688 3052
rect 395896 3000 395948 3052
rect 401324 3000 401376 3052
rect 411904 3068 411956 3120
rect 428740 3068 428792 3120
rect 431224 3068 431276 3120
rect 404912 3000 404964 3052
rect 416688 3000 416740 3052
rect 435824 3000 435876 3052
rect 475108 3000 475160 3052
rect 475384 3000 475436 3052
rect 477500 3000 477552 3052
rect 524972 3068 525024 3120
rect 560760 3068 560812 3120
rect 482284 3000 482336 3052
rect 509884 3000 509936 3052
rect 523684 3000 523736 3052
rect 553584 3000 553636 3052
rect 121828 2796 121880 2848
rect 261484 2796 261536 2848
rect 330024 2796 330076 2848
rect 335544 2796 335596 2848
rect 362224 2864 362276 2916
rect 374092 2932 374144 2984
rect 395988 2932 396040 2984
rect 402520 2932 402572 2984
rect 413468 2932 413520 2984
rect 432328 2932 432380 2984
rect 367284 2864 367336 2916
rect 385868 2864 385920 2916
rect 387064 2864 387116 2916
rect 356704 2796 356756 2848
rect 356152 2660 356204 2712
rect 375840 2796 375892 2848
rect 388444 2796 388496 2848
rect 416044 2796 416096 2848
rect 387064 2728 387116 2780
rect 431316 2864 431368 2916
rect 459652 2932 459704 2984
rect 481088 2932 481140 2984
rect 521016 2932 521068 2984
rect 546500 2932 546552 2984
rect 448980 2864 449032 2916
rect 473912 2864 473964 2916
rect 520924 2864 520976 2916
rect 539324 2864 539376 2916
rect 438124 2796 438176 2848
rect 466828 2796 466880 2848
rect 518164 2796 518216 2848
rect 532240 2796 532292 2848
rect 462044 2728 462096 2780
rect 261024 1096 261076 1148
rect 394148 1028 394200 1080
rect 23112 552 23164 604
rect 23388 552 23440 604
rect 164700 552 164752 604
rect 165528 552 165580 604
rect 165896 552 165948 604
rect 166908 552 166960 604
rect 169392 552 169444 604
rect 169668 552 169720 604
rect 182548 552 182600 604
rect 183468 552 183520 604
rect 183744 552 183796 604
rect 184756 552 184808 604
rect 187240 552 187292 604
rect 187608 552 187660 604
rect 189632 552 189684 604
rect 190368 552 190420 604
rect 281264 552 281316 604
rect 281448 552 281500 604
rect 358544 552 358596 604
rect 358728 552 358780 604
rect 384672 552 384724 604
rect 384948 552 385000 604
rect 389456 595 389508 604
rect 389456 561 389465 595
rect 389465 561 389499 595
rect 389499 561 389508 595
rect 389456 552 389508 561
rect 394240 595 394292 604
rect 394240 561 394249 595
rect 394249 561 394283 595
rect 394283 561 394292 595
rect 394240 552 394292 561
rect 405924 552 405976 604
rect 406108 552 406160 604
rect 463700 552 463752 604
rect 464436 552 464488 604
rect 469220 552 469272 604
rect 470324 552 470376 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 105464 700602 105492 703520
rect 137848 700670 137876 703520
rect 154132 700738 154160 703520
rect 170324 700942 170352 703520
rect 202800 701010 202828 703520
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 170312 700936 170364 700942
rect 170312 700878 170364 700884
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 105452 700596 105504 700602
rect 105452 700538 105504 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 218992 700262 219020 703520
rect 218980 700256 219032 700262
rect 218980 700198 219032 700204
rect 235184 700058 235212 703520
rect 235172 700052 235224 700058
rect 235172 699994 235224 700000
rect 267660 699990 267688 703520
rect 267648 699984 267700 699990
rect 267648 699926 267700 699932
rect 283852 699922 283880 703520
rect 283840 699916 283892 699922
rect 283840 699858 283892 699864
rect 300136 699718 300164 703520
rect 328368 700868 328420 700874
rect 328368 700810 328420 700816
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 300780 584662 300808 699654
rect 321468 696992 321520 696998
rect 321468 696934 321520 696940
rect 320088 673532 320140 673538
rect 320088 673474 320140 673480
rect 315948 650072 316000 650078
rect 315948 650014 316000 650020
rect 313188 626612 313240 626618
rect 313188 626554 313240 626560
rect 309048 603152 309100 603158
rect 309048 603094 309100 603100
rect 300768 584656 300820 584662
rect 300768 584598 300820 584604
rect 304540 583704 304592 583710
rect 304540 583646 304592 583652
rect 298192 583636 298244 583642
rect 298192 583578 298244 583584
rect 262404 583568 262456 583574
rect 262404 583510 262456 583516
rect 256056 583500 256108 583506
rect 256056 583442 256108 583448
rect 251824 583432 251876 583438
rect 4802 583400 4858 583409
rect 251824 583374 251876 583380
rect 4802 583335 4858 583344
rect 6644 583364 6696 583370
rect 4712 583228 4764 583234
rect 4712 583170 4764 583176
rect 3240 583092 3292 583098
rect 3240 583034 3292 583040
rect 3148 568336 3200 568342
rect 3148 568278 3200 568284
rect 3160 567361 3188 568278
rect 3146 567352 3202 567361
rect 3146 567287 3202 567296
rect 3148 553376 3200 553382
rect 3148 553318 3200 553324
rect 3160 553081 3188 553318
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3056 539096 3108 539102
rect 3056 539038 3108 539044
rect 3068 538665 3096 539038
rect 3054 538656 3110 538665
rect 3054 538591 3110 538600
rect 3148 510264 3200 510270
rect 3148 510206 3200 510212
rect 3160 509969 3188 510206
rect 3146 509960 3202 509969
rect 3146 509895 3202 509904
rect 2780 495780 2832 495786
rect 2780 495722 2832 495728
rect 2792 495553 2820 495722
rect 2778 495544 2834 495553
rect 2778 495479 2834 495488
rect 3148 481296 3200 481302
rect 3148 481238 3200 481244
rect 3160 481137 3188 481238
rect 3146 481128 3202 481137
rect 3146 481063 3202 481072
rect 3252 452441 3280 583034
rect 4068 582752 4120 582758
rect 4068 582694 4120 582700
rect 3700 582480 3752 582486
rect 3700 582422 3752 582428
rect 3332 578536 3384 578542
rect 3332 578478 3384 578484
rect 3238 452432 3294 452441
rect 3238 452367 3294 452376
rect 2780 438592 2832 438598
rect 2780 438534 2832 438540
rect 2792 438025 2820 438534
rect 2778 438016 2834 438025
rect 2778 437951 2834 437960
rect 2780 424856 2832 424862
rect 2780 424798 2832 424804
rect 2792 423745 2820 424798
rect 2778 423736 2834 423745
rect 2778 423671 2834 423680
rect 3240 395888 3292 395894
rect 3240 395830 3292 395836
rect 3252 395049 3280 395830
rect 3238 395040 3294 395049
rect 3238 394975 3294 394984
rect 2780 380792 2832 380798
rect 2780 380734 2832 380740
rect 2792 380633 2820 380734
rect 2778 380624 2834 380633
rect 2778 380559 2834 380568
rect 3344 366217 3372 578478
rect 3608 578400 3660 578406
rect 3608 578342 3660 578348
rect 3424 578332 3476 578338
rect 3424 578274 3476 578280
rect 3330 366208 3386 366217
rect 3330 366143 3386 366152
rect 3332 324284 3384 324290
rect 3332 324226 3384 324232
rect 3344 323105 3372 324226
rect 3330 323096 3386 323105
rect 3330 323031 3386 323040
rect 3332 280152 3384 280158
rect 3330 280120 3332 280129
rect 3384 280120 3386 280129
rect 3330 280055 3386 280064
rect 3146 252512 3202 252521
rect 3146 252447 3202 252456
rect 3160 251297 3188 252447
rect 3146 251288 3202 251297
rect 3146 251223 3202 251232
rect 3332 237380 3384 237386
rect 3332 237322 3384 237328
rect 3344 237017 3372 237322
rect 3330 237008 3386 237017
rect 3330 236943 3386 236952
rect 2780 223100 2832 223106
rect 2780 223042 2832 223048
rect 2792 222601 2820 223042
rect 2778 222592 2834 222601
rect 2778 222527 2834 222536
rect 3332 151768 3384 151774
rect 3332 151710 3384 151716
rect 3344 150793 3372 151710
rect 3330 150784 3386 150793
rect 3330 150719 3386 150728
rect 2780 136536 2832 136542
rect 2780 136478 2832 136484
rect 2792 136377 2820 136478
rect 2778 136368 2834 136377
rect 2778 136303 2834 136312
rect 2780 122324 2832 122330
rect 2780 122266 2832 122272
rect 2792 122097 2820 122266
rect 2778 122088 2834 122097
rect 2778 122023 2834 122032
rect 3436 93265 3464 578274
rect 3516 578264 3568 578270
rect 3516 578206 3568 578212
rect 3528 107681 3556 578206
rect 3620 179489 3648 578342
rect 3712 193905 3740 582422
rect 3976 579964 4028 579970
rect 3976 579906 4028 579912
rect 3792 579896 3844 579902
rect 3792 579838 3844 579844
rect 3804 208185 3832 579838
rect 3884 578468 3936 578474
rect 3884 578410 3936 578416
rect 3896 265713 3924 578410
rect 3988 294409 4016 579906
rect 4080 308825 4108 582694
rect 4724 495786 4752 583170
rect 4712 495780 4764 495786
rect 4712 495722 4764 495728
rect 4066 308816 4122 308825
rect 4066 308751 4122 308760
rect 3974 294400 4030 294409
rect 3974 294335 4030 294344
rect 3882 265704 3938 265713
rect 3882 265639 3938 265648
rect 3790 208176 3846 208185
rect 3790 208111 3846 208120
rect 3698 193896 3754 193905
rect 3698 193831 3754 193840
rect 3606 179480 3662 179489
rect 3606 179415 3662 179424
rect 3514 107672 3570 107681
rect 3514 107607 3570 107616
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 2780 79824 2832 79830
rect 2780 79766 2832 79772
rect 2792 78985 2820 79766
rect 2778 78976 2834 78985
rect 2778 78911 2834 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 4816 50522 4844 583335
rect 6644 583306 6696 583312
rect 6368 583296 6420 583302
rect 6368 583238 6420 583244
rect 5356 583160 5408 583166
rect 5356 583102 5408 583108
rect 5264 582888 5316 582894
rect 5264 582830 5316 582836
rect 5172 582548 5224 582554
rect 5172 582490 5224 582496
rect 5080 582412 5132 582418
rect 5080 582354 5132 582360
rect 4988 579828 5040 579834
rect 4988 579770 5040 579776
rect 4896 579760 4948 579766
rect 4896 579702 4948 579708
rect 4908 79830 4936 579702
rect 5000 122330 5028 579770
rect 5092 136542 5120 582354
rect 5184 223106 5212 582490
rect 5276 380798 5304 582830
rect 5368 424862 5396 583102
rect 5448 583024 5500 583030
rect 5448 582966 5500 582972
rect 5460 438598 5488 582966
rect 6276 580032 6328 580038
rect 6276 579974 6328 579980
rect 6184 579692 6236 579698
rect 6184 579634 6236 579640
rect 5448 438592 5500 438598
rect 5448 438534 5500 438540
rect 5356 424856 5408 424862
rect 5356 424798 5408 424804
rect 5264 380792 5316 380798
rect 5264 380734 5316 380740
rect 5172 223100 5224 223106
rect 5172 223042 5224 223048
rect 5080 136536 5132 136542
rect 5080 136478 5132 136484
rect 4988 122324 5040 122330
rect 4988 122266 5040 122272
rect 4896 79824 4948 79830
rect 4896 79766 4948 79772
rect 2780 50516 2832 50522
rect 2780 50458 2832 50464
rect 4804 50516 4856 50522
rect 4804 50458 4856 50464
rect 2792 50153 2820 50458
rect 2778 50144 2834 50153
rect 2778 50079 2834 50088
rect 6196 35902 6224 579634
rect 6288 395894 6316 579974
rect 6380 481302 6408 583238
rect 6460 580100 6512 580106
rect 6460 580042 6512 580048
rect 6472 510270 6500 580042
rect 6552 578604 6604 578610
rect 6552 578546 6604 578552
rect 6564 539102 6592 578546
rect 6656 553382 6684 583306
rect 14464 582956 14516 582962
rect 14464 582898 14516 582904
rect 6736 580168 6788 580174
rect 6736 580110 6788 580116
rect 6748 568342 6776 580110
rect 6736 568336 6788 568342
rect 6736 568278 6788 568284
rect 6644 553376 6696 553382
rect 6644 553318 6696 553324
rect 6552 539096 6604 539102
rect 6552 539038 6604 539044
rect 6460 510264 6512 510270
rect 6460 510206 6512 510212
rect 6368 481296 6420 481302
rect 6368 481238 6420 481244
rect 6276 395888 6328 395894
rect 6276 395830 6328 395836
rect 13084 337408 13136 337414
rect 10322 337376 10378 337385
rect 13084 337350 13136 337356
rect 10322 337311 10378 337320
rect 3148 35896 3200 35902
rect 3146 35864 3148 35873
rect 6184 35896 6236 35902
rect 3200 35864 3202 35873
rect 6184 35838 6236 35844
rect 3146 35799 3202 35808
rect 3146 11656 3202 11665
rect 3146 11591 3202 11600
rect 3160 7177 3188 11591
rect 8852 7676 8904 7682
rect 8852 7618 8904 7624
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 3146 7168 3202 7177
rect 3146 7103 3202 7112
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4898
rect 4080 480 4108 7550
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8864 480 8892 7618
rect 10336 3466 10364 337311
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10048 3324 10100 3330
rect 10048 3266 10100 3272
rect 10060 480 10088 3266
rect 11256 480 11284 3538
rect 12452 480 12480 5034
rect 13096 3330 13124 337350
rect 14476 324290 14504 582898
rect 15844 582820 15896 582826
rect 15844 582762 15896 582768
rect 14464 324284 14516 324290
rect 14464 324226 14516 324232
rect 15856 280158 15884 582762
rect 17224 582684 17276 582690
rect 17224 582626 17276 582632
rect 15844 280152 15896 280158
rect 15844 280094 15896 280100
rect 17236 237386 17264 582626
rect 24124 582616 24176 582622
rect 24124 582558 24176 582564
rect 31022 582584 31078 582593
rect 19984 337476 20036 337482
rect 19984 337418 20036 337424
rect 17224 237380 17276 237386
rect 17224 237322 17276 237328
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13084 3324 13136 3330
rect 13084 3266 13136 3272
rect 13648 480 13676 8910
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14844 480 14872 3470
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 16040 480 16068 3402
rect 17236 480 17264 5102
rect 18340 480 18368 8978
rect 19996 3602 20024 337418
rect 24136 151774 24164 582558
rect 31022 582519 31078 582528
rect 28264 337544 28316 337550
rect 28264 337486 28316 337492
rect 24124 151768 24176 151774
rect 24124 151710 24176 151716
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 20720 3800 20772 3806
rect 20720 3742 20772 3748
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19536 480 19564 3334
rect 20732 480 20760 3742
rect 21928 480 21956 7686
rect 23400 610 23428 11698
rect 27896 9104 27948 9110
rect 27896 9046 27948 9052
rect 26700 7812 26752 7818
rect 26700 7754 26752 7760
rect 24308 3664 24360 3670
rect 24308 3606 24360 3612
rect 23112 604 23164 610
rect 23112 546 23164 552
rect 23388 604 23440 610
rect 23388 546 23440 552
rect 23124 480 23152 546
rect 24320 480 24348 3606
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25516 480 25544 3538
rect 26712 480 26740 7754
rect 27908 480 27936 9046
rect 28276 3398 28304 337486
rect 31036 64870 31064 582519
rect 251836 579972 251864 583374
rect 256068 579972 256096 583442
rect 258172 581052 258224 581058
rect 258172 580994 258224 581000
rect 258184 579972 258212 580994
rect 262416 579972 262444 583510
rect 293958 583128 294014 583137
rect 293958 583063 294014 583072
rect 289728 581460 289780 581466
rect 289728 581402 289780 581408
rect 287612 581392 287664 581398
rect 287612 581334 287664 581340
rect 283472 581324 283524 581330
rect 283472 581266 283524 581272
rect 281356 581256 281408 581262
rect 281356 581198 281408 581204
rect 275008 581188 275060 581194
rect 275008 581130 275060 581136
rect 264520 581120 264572 581126
rect 264520 581062 264572 581068
rect 264532 579972 264560 581062
rect 268660 580304 268712 580310
rect 268660 580246 268712 580252
rect 268672 579972 268700 580246
rect 275020 579972 275048 581130
rect 281368 579972 281396 581198
rect 283484 579972 283512 581266
rect 287624 579972 287652 581334
rect 289740 579972 289768 581402
rect 293972 579972 294000 583063
rect 296076 581528 296128 581534
rect 296076 581470 296128 581476
rect 296088 579972 296116 581470
rect 298204 579972 298232 583578
rect 300306 583264 300362 583273
rect 300306 583199 300362 583208
rect 300320 579972 300348 583199
rect 302424 581596 302476 581602
rect 302424 581538 302476 581544
rect 302436 579972 302464 581538
rect 304552 579972 304580 583646
rect 306564 580236 306616 580242
rect 306564 580178 306616 580184
rect 306576 579972 306604 580178
rect 309060 579986 309088 603094
rect 311808 592068 311860 592074
rect 311808 592010 311860 592016
rect 311820 580122 311848 592010
rect 308706 579958 309088 579986
rect 311268 580094 311848 580122
rect 311268 579850 311296 580094
rect 313200 579986 313228 626554
rect 312938 579958 313228 579986
rect 315960 579850 315988 650014
rect 317328 638988 317380 638994
rect 317328 638930 317380 638936
rect 317340 579986 317368 638930
rect 320100 580122 320128 673474
rect 317170 579958 317368 579986
rect 319732 580094 320128 580122
rect 319732 579850 319760 580094
rect 321480 579986 321508 696934
rect 324228 685908 324280 685914
rect 324228 685850 324280 685856
rect 321402 579958 321508 579986
rect 324240 579850 324268 685850
rect 325516 584452 325568 584458
rect 325516 584394 325568 584400
rect 325528 579972 325556 584394
rect 328380 579850 328408 700810
rect 329748 700800 329800 700806
rect 329748 700742 329800 700748
rect 329760 579972 329788 700742
rect 332520 699718 332548 703520
rect 336648 700188 336700 700194
rect 336648 700130 336700 700136
rect 335268 700120 335320 700126
rect 335268 700062 335320 700068
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 331864 584520 331916 584526
rect 331864 584462 331916 584468
rect 331876 579972 331904 584462
rect 335280 580122 335308 700062
rect 334452 580094 335308 580122
rect 334452 579850 334480 580094
rect 336660 579850 336688 700130
rect 343548 699848 343600 699854
rect 343548 699790 343600 699796
rect 340788 699780 340840 699786
rect 340788 699722 340840 699728
rect 338212 584588 338264 584594
rect 338212 584530 338264 584536
rect 338224 579972 338252 584530
rect 340800 579986 340828 699722
rect 340354 579958 340828 579986
rect 343560 579850 343588 699790
rect 348804 699718 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365208 703474
rect 358820 701004 358872 701010
rect 358820 700946 358872 700952
rect 356060 700052 356112 700058
rect 356060 699994 356112 700000
rect 351920 699984 351972 699990
rect 351920 699926 351972 699932
rect 346400 699712 346452 699718
rect 346400 699654 346452 699660
rect 347780 699712 347832 699718
rect 347780 699654 347832 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 344468 584724 344520 584730
rect 344468 584666 344520 584672
rect 344480 579972 344508 584666
rect 346412 579986 346440 699654
rect 346412 579958 346610 579986
rect 310822 579822 311296 579850
rect 315054 579822 315988 579850
rect 319286 579822 319760 579850
rect 323426 579822 324268 579850
rect 327658 579822 328408 579850
rect 334006 579822 334480 579850
rect 336122 579822 336688 579850
rect 342378 579822 343588 579850
rect 347792 579850 347820 699654
rect 350816 584656 350868 584662
rect 350816 584598 350868 584604
rect 350828 579972 350856 584598
rect 351932 579850 351960 699926
rect 354680 699916 354732 699922
rect 354680 699858 354732 699864
rect 354692 579986 354720 699858
rect 354692 579958 355074 579986
rect 356072 579850 356100 699994
rect 358832 579850 358860 700946
rect 362960 700936 363012 700942
rect 362960 700878 363012 700884
rect 360200 700256 360252 700262
rect 360200 700198 360252 700204
rect 360212 580122 360240 700198
rect 360212 580094 360884 580122
rect 360856 579850 360884 580094
rect 362972 579986 363000 700878
rect 364340 700664 364392 700670
rect 364340 700606 364392 700612
rect 364352 580122 364380 700606
rect 365180 687818 365208 703446
rect 367100 700732 367152 700738
rect 367100 700674 367152 700680
rect 364616 687812 364668 687818
rect 364616 687754 364668 687760
rect 365168 687812 365220 687818
rect 365168 687754 365220 687760
rect 364628 685846 364656 687754
rect 364616 685840 364668 685846
rect 364616 685782 364668 685788
rect 364524 676252 364576 676258
rect 364524 676194 364576 676200
rect 364536 669338 364564 676194
rect 364536 669310 364748 669338
rect 364720 650026 364748 669310
rect 364536 649998 364748 650026
rect 364536 630714 364564 649998
rect 364536 630686 364656 630714
rect 364628 618254 364656 630686
rect 364616 618248 364668 618254
rect 364616 618190 364668 618196
rect 364524 608660 364576 608666
rect 364524 608602 364576 608608
rect 364536 601746 364564 608602
rect 364536 601718 364656 601746
rect 364628 598942 364656 601718
rect 364616 598936 364668 598942
rect 364616 598878 364668 598884
rect 364708 589348 364760 589354
rect 364708 589290 364760 589296
rect 364720 584730 364748 589290
rect 364708 584724 364760 584730
rect 364708 584666 364760 584672
rect 364352 580094 365208 580122
rect 365180 579986 365208 580094
rect 362972 579958 363446 579986
rect 365180 579958 365562 579986
rect 367112 579850 367140 700674
rect 368480 700596 368532 700602
rect 368480 700538 368532 700544
rect 368492 580122 368520 700538
rect 374000 700528 374052 700534
rect 374000 700470 374052 700476
rect 371240 700460 371292 700466
rect 371240 700402 371292 700408
rect 368492 580094 369348 580122
rect 369320 579850 369348 580094
rect 371252 579850 371280 700402
rect 374012 579972 374040 700470
rect 375380 700392 375432 700398
rect 375380 700334 375432 700340
rect 378138 700360 378194 700369
rect 375392 579850 375420 700334
rect 378138 700295 378194 700304
rect 379520 700324 379572 700330
rect 378152 579986 378180 700295
rect 379520 700266 379572 700272
rect 378152 579958 378258 579986
rect 379532 579850 379560 700266
rect 397472 699786 397500 703520
rect 413664 699854 413692 703520
rect 413652 699848 413704 699854
rect 413652 699790 413704 699796
rect 397460 699780 397512 699786
rect 397460 699722 397512 699728
rect 429856 688634 429884 703520
rect 462332 700126 462360 703520
rect 478524 700194 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700188 478564 700194
rect 478512 700130 478564 700136
rect 462320 700120 462372 700126
rect 462320 700062 462372 700068
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 429396 685930 429424 688570
rect 494900 686089 494928 703446
rect 527192 700874 527220 703520
rect 527180 700868 527232 700874
rect 527180 700810 527232 700816
rect 543476 700806 543504 703520
rect 543464 700800 543516 700806
rect 543464 700742 543516 700748
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 429304 685902 429424 685930
rect 494242 685944 494298 685953
rect 429304 684486 429332 685902
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 382280 681760 382332 681766
rect 382280 681702 382332 681708
rect 382292 579986 382320 681702
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 386420 667956 386472 667962
rect 386420 667898 386472 667904
rect 383660 652792 383712 652798
rect 383660 652734 383712 652740
rect 382292 579958 382398 579986
rect 383672 579850 383700 652734
rect 386432 579986 386460 667898
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 429672 659682 429700 666538
rect 429488 659654 429700 659682
rect 494164 659682 494192 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 429488 647290 429516 659654
rect 494256 654158 494284 659654
rect 559208 659654 559420 659682
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 429396 640422 429424 647226
rect 494072 644450 494100 654094
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 494072 644422 494284 644450
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 429488 630698 429516 640358
rect 494256 634846 494284 644422
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 429304 630578 429332 630634
rect 429304 630550 429424 630578
rect 387800 623824 387852 623830
rect 387800 623766 387852 623772
rect 386432 579958 386630 579986
rect 387812 579850 387840 623766
rect 429396 621058 429424 630550
rect 494072 625138 494100 634782
rect 559208 630698 559236 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 494072 625110 494284 625138
rect 429396 621030 429516 621058
rect 429488 611386 429516 621030
rect 494256 615534 494284 625110
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 559116 621030 559236 621058
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 429304 611266 429332 611322
rect 429304 611238 429424 611266
rect 391940 610020 391992 610026
rect 391940 609962 391992 609968
rect 390560 594856 390612 594862
rect 390560 594798 390612 594804
rect 390572 579986 390600 594798
rect 391952 580122 391980 609962
rect 429396 608598 429424 611238
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 494072 605826 494100 615470
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 494072 605798 494284 605826
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 429580 598942 429608 601666
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 494256 596222 494284 605798
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 429672 584594 429700 589290
rect 429660 584588 429712 584594
rect 429660 584530 429712 584536
rect 494256 584526 494284 596006
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 494244 584520 494296 584526
rect 494244 584462 494296 584468
rect 559392 584458 559420 589290
rect 559380 584452 559432 584458
rect 559380 584394 559432 584400
rect 471244 583704 471296 583710
rect 471244 583646 471296 583652
rect 469772 583636 469824 583642
rect 469772 583578 469824 583584
rect 460294 583400 460350 583409
rect 399208 583364 399260 583370
rect 460294 583335 460350 583344
rect 399208 583306 399260 583312
rect 395068 580168 395120 580174
rect 391952 580094 392532 580122
rect 395068 580110 395120 580116
rect 390572 579958 390862 579986
rect 392504 579850 392532 580094
rect 395080 579972 395108 580110
rect 399220 579972 399248 583306
rect 403440 583296 403492 583302
rect 403440 583238 403492 583244
rect 401324 580100 401376 580106
rect 401324 580042 401376 580048
rect 401336 579972 401364 580042
rect 403452 579972 403480 583238
rect 405556 583228 405608 583234
rect 405556 583170 405608 583176
rect 405568 579972 405596 583170
rect 409788 583160 409840 583166
rect 409788 583102 409840 583108
rect 407672 583092 407724 583098
rect 407672 583034 407724 583040
rect 407684 579972 407712 583034
rect 409800 579972 409828 583102
rect 411904 583024 411956 583030
rect 411904 582966 411956 582972
rect 420274 582992 420330 583001
rect 411916 579972 411944 582966
rect 420274 582927 420330 582936
rect 424508 582956 424560 582962
rect 418160 582888 418212 582894
rect 418160 582830 418212 582836
rect 414112 580032 414164 580038
rect 414046 579980 414112 579986
rect 414046 579974 414164 579980
rect 414046 579958 414152 579974
rect 418172 579972 418200 582830
rect 420288 579972 420316 582927
rect 424508 582898 424560 582904
rect 422392 582752 422444 582758
rect 422392 582694 422444 582700
rect 422404 579972 422432 582694
rect 424520 579972 424548 582898
rect 432970 582856 433026 582865
rect 430856 582820 430908 582826
rect 432970 582791 433026 582800
rect 430856 582762 430908 582768
rect 426452 579970 426650 579986
rect 430868 579972 430896 582762
rect 432984 579972 433012 582791
rect 445574 582720 445630 582729
rect 437112 582684 437164 582690
rect 445574 582655 445630 582664
rect 437112 582626 437164 582632
rect 434996 582548 435048 582554
rect 434996 582490 435048 582496
rect 435008 579972 435036 582490
rect 437124 579972 437152 582626
rect 443460 582480 443512 582486
rect 443460 582422 443512 582428
rect 443472 579972 443500 582422
rect 445588 579972 445616 582655
rect 449808 582616 449860 582622
rect 449808 582558 449860 582564
rect 447692 582412 447744 582418
rect 447692 582354 447744 582360
rect 447704 579972 447732 582354
rect 449820 579972 449848 582558
rect 460308 579972 460336 583335
rect 462410 582584 462466 582593
rect 462410 582519 462466 582528
rect 462424 579972 462452 582519
rect 469588 581596 469640 581602
rect 469588 581538 469640 581544
rect 426440 579964 426650 579970
rect 426492 579958 426650 579964
rect 426440 579906 426492 579912
rect 438860 579896 438912 579902
rect 347792 579822 348726 579850
rect 351932 579822 352958 579850
rect 356072 579822 357190 579850
rect 358832 579822 359306 579850
rect 360856 579822 361330 579850
rect 367112 579822 367678 579850
rect 369320 579822 369794 579850
rect 371252 579822 371910 579850
rect 375392 579822 376142 579850
rect 379532 579822 380282 579850
rect 383672 579822 384514 579850
rect 387812 579822 388746 579850
rect 392504 579822 392978 579850
rect 438912 579844 439254 579850
rect 438860 579838 439254 579844
rect 438872 579822 439254 579838
rect 451568 579834 451950 579850
rect 451556 579828 451950 579834
rect 451608 579822 451950 579828
rect 451556 579770 451608 579776
rect 458272 579760 458324 579766
rect 458206 579708 458272 579714
rect 458206 579702 458324 579708
rect 458206 579686 458312 579702
rect 464264 579698 464554 579714
rect 464252 579692 464554 579698
rect 464304 579686 464554 579692
rect 464252 579634 464304 579640
rect 270802 579426 271184 579442
rect 270802 579420 271196 579426
rect 270802 579414 271144 579420
rect 271144 579362 271196 579368
rect 254124 579352 254176 579358
rect 231122 579320 231178 579329
rect 230874 579278 231122 579306
rect 232962 579320 233018 579329
rect 232898 579278 232962 579306
rect 231122 579255 231178 579264
rect 235262 579320 235318 579329
rect 235014 579278 235262 579306
rect 232962 579255 233018 579264
rect 237194 579320 237250 579329
rect 237130 579278 237194 579306
rect 235262 579255 235318 579264
rect 239402 579320 239458 579329
rect 239246 579278 239402 579306
rect 237194 579255 237250 579264
rect 241426 579320 241482 579329
rect 241362 579278 241426 579306
rect 239402 579255 239458 579264
rect 243634 579320 243690 579329
rect 243478 579278 243634 579306
rect 241426 579255 241482 579264
rect 243634 579255 243690 579264
rect 245382 579320 245438 579329
rect 247866 579320 247922 579329
rect 245438 579278 245594 579306
rect 247710 579278 247866 579306
rect 245382 579255 245438 579264
rect 247866 579255 247922 579264
rect 249522 579320 249578 579329
rect 249578 579278 249734 579306
rect 253966 579300 254124 579306
rect 260656 579352 260708 579358
rect 253966 579294 254176 579300
rect 260314 579300 260656 579306
rect 266820 579352 266872 579358
rect 260314 579294 260708 579300
rect 266662 579300 266820 579306
rect 273168 579352 273220 579358
rect 266662 579294 266872 579300
rect 272918 579300 273168 579306
rect 277308 579352 277360 579358
rect 272918 579294 273220 579300
rect 277150 579300 277308 579306
rect 279608 579352 279660 579358
rect 277150 579294 277360 579300
rect 279266 579300 279608 579306
rect 285772 579352 285824 579358
rect 279266 579294 279660 579300
rect 285614 579300 285772 579306
rect 292120 579352 292172 579358
rect 285614 579294 285824 579300
rect 291870 579300 292120 579306
rect 291870 579294 292172 579300
rect 396724 579352 396776 579358
rect 415676 579352 415728 579358
rect 396776 579300 397118 579306
rect 396724 579294 397118 579300
rect 428372 579352 428424 579358
rect 415728 579300 416070 579306
rect 415676 579294 416070 579300
rect 441068 579352 441120 579358
rect 428424 579300 428766 579306
rect 428372 579294 428766 579300
rect 453580 579352 453632 579358
rect 441120 579300 441370 579306
rect 441068 579294 441370 579300
rect 455788 579352 455840 579358
rect 453632 579300 453974 579306
rect 453580 579294 453974 579300
rect 466458 579320 466514 579329
rect 455840 579300 456090 579306
rect 455788 579294 456090 579300
rect 253966 579278 254164 579294
rect 260314 579278 260696 579294
rect 266662 579278 266860 579294
rect 272918 579278 273208 579294
rect 277150 579278 277348 579294
rect 279266 579278 279648 579294
rect 285614 579278 285812 579294
rect 291870 579278 292160 579294
rect 396736 579278 397118 579294
rect 415688 579278 416070 579294
rect 428384 579278 428766 579294
rect 441080 579278 441370 579294
rect 453592 579278 453974 579294
rect 455800 579278 456090 579294
rect 249522 579255 249578 579264
rect 468574 579320 468630 579329
rect 466514 579278 466670 579306
rect 466458 579255 466514 579264
rect 468630 579278 468786 579306
rect 468574 579255 468630 579264
rect 469600 557530 469628 581538
rect 469680 581528 469732 581534
rect 469680 581470 469732 581476
rect 469588 557524 469640 557530
rect 469588 557466 469640 557472
rect 469692 510610 469720 581470
rect 469680 510604 469732 510610
rect 469680 510546 469732 510552
rect 469784 499526 469812 583578
rect 470508 581460 470560 581466
rect 470508 581402 470560 581408
rect 470416 581392 470468 581398
rect 470416 581334 470468 581340
rect 470324 581324 470376 581330
rect 470324 581266 470376 581272
rect 470140 581256 470192 581262
rect 470140 581198 470192 581204
rect 470048 581188 470100 581194
rect 470048 581130 470100 581136
rect 469864 580304 469916 580310
rect 469864 580246 469916 580252
rect 469772 499520 469824 499526
rect 469772 499462 469824 499468
rect 231044 340190 231426 340218
rect 232516 340190 232898 340218
rect 244752 340190 245226 340218
rect 246224 340190 246698 340218
rect 282012 340190 282394 340218
rect 290292 340190 290766 340218
rect 291764 340190 292238 340218
rect 294708 340190 295182 340218
rect 325068 340190 325542 340218
rect 337396 340190 337778 340218
rect 340340 340190 340722 340218
rect 357912 340190 358386 340218
rect 373092 340190 373566 340218
rect 374564 340190 375038 340218
rect 386800 340190 387274 340218
rect 389744 340190 390218 340218
rect 422970 340190 423444 340218
rect 424442 340190 424916 340218
rect 229112 340054 230046 340082
rect 79324 338088 79376 338094
rect 79324 338030 79376 338036
rect 71044 338020 71096 338026
rect 71044 337962 71096 337968
rect 66904 337952 66956 337958
rect 66904 337894 66956 337900
rect 61384 337884 61436 337890
rect 61384 337826 61436 337832
rect 57244 337816 57296 337822
rect 57244 337758 57296 337764
rect 35164 337748 35216 337754
rect 35164 337690 35216 337696
rect 32404 337612 32456 337618
rect 32404 337554 32456 337560
rect 31024 64864 31076 64870
rect 31024 64806 31076 64812
rect 31668 13116 31720 13122
rect 31668 13058 31720 13064
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29104 480 29132 3334
rect 30300 480 30328 7822
rect 31680 626 31708 13058
rect 32416 3398 32444 337554
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 31496 598 31708 626
rect 31496 480 31524 598
rect 32692 480 32720 3674
rect 33888 480 33916 7890
rect 35176 3806 35204 337690
rect 39304 337680 39356 337686
rect 39304 337622 39356 337628
rect 37372 8016 37424 8022
rect 37372 7958 37424 7964
rect 35164 3800 35216 3806
rect 35164 3742 35216 3748
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 34992 480 35020 3334
rect 36176 3052 36228 3058
rect 36176 2994 36228 3000
rect 36188 480 36216 2994
rect 37384 480 37412 7958
rect 38568 3800 38620 3806
rect 38568 3742 38620 3748
rect 38580 480 38608 3742
rect 39316 3058 39344 337622
rect 56508 10396 56560 10402
rect 56508 10338 56560 10344
rect 53748 10328 53800 10334
rect 53748 10270 53800 10276
rect 49332 9240 49384 9246
rect 49332 9182 49384 9188
rect 44548 9172 44600 9178
rect 44548 9114 44600 9120
rect 40960 8084 41012 8090
rect 40960 8026 41012 8032
rect 39764 3868 39816 3874
rect 39764 3810 39816 3816
rect 39304 3052 39356 3058
rect 39304 2994 39356 3000
rect 39776 480 39804 3810
rect 40972 480 41000 8026
rect 42156 3324 42208 3330
rect 42156 3266 42208 3272
rect 42168 480 42196 3266
rect 43352 3256 43404 3262
rect 43352 3198 43404 3204
rect 43364 480 43392 3198
rect 44560 480 44588 9114
rect 48136 5228 48188 5234
rect 48136 5170 48188 5176
rect 46940 4004 46992 4010
rect 46940 3946 46992 3952
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45756 480 45784 3878
rect 46952 480 46980 3946
rect 48148 480 48176 5170
rect 49344 480 49372 9182
rect 51630 6216 51686 6225
rect 51630 6151 51686 6160
rect 50528 4072 50580 4078
rect 50528 4014 50580 4020
rect 50540 480 50568 4014
rect 51644 480 51672 6151
rect 53760 3194 53788 10270
rect 55220 6180 55272 6186
rect 55220 6122 55272 6128
rect 52828 3188 52880 3194
rect 52828 3130 52880 3136
rect 53748 3188 53800 3194
rect 53748 3130 53800 3136
rect 54024 3188 54076 3194
rect 54024 3130 54076 3136
rect 52840 480 52868 3130
rect 54036 480 54064 3130
rect 55232 480 55260 6122
rect 56520 3482 56548 10338
rect 56428 3454 56548 3482
rect 56428 480 56456 3454
rect 57256 3398 57284 337758
rect 60648 10464 60700 10470
rect 60648 10406 60700 10412
rect 58808 6248 58860 6254
rect 58808 6190 58860 6196
rect 57612 4140 57664 4146
rect 57612 4082 57664 4088
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 57624 480 57652 4082
rect 58820 480 58848 6190
rect 60660 3398 60688 10406
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60016 480 60044 3334
rect 61396 3262 61424 337826
rect 64788 10532 64840 10538
rect 64788 10474 64840 10480
rect 62396 6316 62448 6322
rect 62396 6258 62448 6264
rect 61384 3256 61436 3262
rect 61384 3198 61436 3204
rect 61200 3120 61252 3126
rect 61200 3062 61252 3068
rect 61212 480 61240 3062
rect 62408 480 62436 6258
rect 64696 3392 64748 3398
rect 64696 3334 64748 3340
rect 63592 3256 63644 3262
rect 63592 3198 63644 3204
rect 63604 480 63632 3198
rect 64708 1714 64736 3334
rect 64800 3262 64828 10474
rect 65984 6384 66036 6390
rect 65984 6326 66036 6332
rect 64788 3256 64840 3262
rect 64788 3198 64840 3204
rect 64708 1686 64828 1714
rect 64800 480 64828 1686
rect 65996 480 66024 6326
rect 66916 3330 66944 337894
rect 69480 6452 69532 6458
rect 69480 6394 69532 6400
rect 67180 5296 67232 5302
rect 67180 5238 67232 5244
rect 66904 3324 66956 3330
rect 66904 3266 66956 3272
rect 67192 480 67220 5238
rect 68284 3052 68336 3058
rect 68284 2994 68336 3000
rect 68296 480 68324 2994
rect 69492 480 69520 6394
rect 70676 3324 70728 3330
rect 70676 3266 70728 3272
rect 70688 480 70716 3266
rect 71056 3194 71084 337962
rect 77944 337340 77996 337346
rect 77944 337282 77996 337288
rect 74448 14476 74500 14482
rect 74448 14418 74500 14424
rect 71688 13184 71740 13190
rect 71688 13126 71740 13132
rect 71700 3330 71728 13126
rect 73068 6520 73120 6526
rect 73068 6462 73120 6468
rect 71688 3324 71740 3330
rect 71688 3266 71740 3272
rect 71872 3324 71924 3330
rect 71872 3266 71924 3272
rect 71044 3188 71096 3194
rect 71044 3130 71096 3136
rect 71884 480 71912 3266
rect 73080 480 73108 6462
rect 74460 3380 74488 14418
rect 76656 6588 76708 6594
rect 76656 6530 76708 6536
rect 74276 3352 74488 3380
rect 74276 480 74304 3352
rect 75460 3052 75512 3058
rect 75460 2994 75512 3000
rect 75472 480 75500 2994
rect 76668 480 76696 6530
rect 77852 3256 77904 3262
rect 77852 3198 77904 3204
rect 77864 480 77892 3198
rect 77956 3126 77984 337282
rect 78588 14544 78640 14550
rect 78588 14486 78640 14492
rect 78600 3262 78628 14486
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 79048 3188 79100 3194
rect 79048 3130 79100 3136
rect 77944 3120 77996 3126
rect 77944 3062 77996 3068
rect 79060 480 79088 3130
rect 79336 2922 79364 338030
rect 84844 337340 84896 337346
rect 84844 337282 84896 337288
rect 82728 14612 82780 14618
rect 82728 14554 82780 14560
rect 80244 8152 80296 8158
rect 80244 8094 80296 8100
rect 79324 2916 79376 2922
rect 79324 2858 79376 2864
rect 80256 480 80284 8094
rect 82740 3262 82768 14554
rect 83832 8220 83884 8226
rect 83832 8162 83884 8168
rect 81440 3256 81492 3262
rect 81440 3198 81492 3204
rect 82728 3256 82780 3262
rect 82728 3198 82780 3204
rect 81452 480 81480 3198
rect 82636 3120 82688 3126
rect 82636 3062 82688 3068
rect 82648 480 82676 3062
rect 83844 480 83872 8162
rect 84856 3262 84884 337282
rect 132500 337272 132552 337278
rect 132498 337240 132500 337249
rect 142068 337272 142120 337278
rect 132552 337240 132554 337249
rect 97264 337204 97316 337210
rect 132498 337175 132554 337184
rect 142066 337240 142068 337249
rect 151820 337272 151872 337278
rect 142120 337240 142122 337249
rect 142066 337175 142122 337184
rect 151818 337240 151820 337249
rect 161388 337272 161440 337278
rect 151872 337240 151874 337249
rect 151818 337175 151874 337184
rect 161386 337240 161388 337249
rect 171140 337272 171192 337278
rect 161440 337240 161442 337249
rect 161386 337175 161442 337184
rect 171138 337240 171140 337249
rect 180708 337272 180760 337278
rect 171192 337240 171194 337249
rect 171138 337175 171194 337184
rect 180706 337240 180708 337249
rect 190460 337272 190512 337278
rect 180760 337240 180762 337249
rect 180706 337175 180762 337184
rect 190458 337240 190460 337249
rect 200028 337272 200080 337278
rect 190512 337240 190514 337249
rect 190458 337175 190514 337184
rect 200026 337240 200028 337249
rect 209780 337272 209832 337278
rect 200080 337240 200082 337249
rect 200026 337175 200082 337184
rect 209778 337240 209780 337249
rect 219348 337272 219400 337278
rect 209832 337240 209834 337249
rect 209778 337175 209834 337184
rect 219346 337240 219348 337249
rect 219400 337240 219402 337249
rect 219346 337175 219402 337184
rect 97264 337146 97316 337152
rect 95884 337068 95936 337074
rect 95884 337010 95936 337016
rect 92388 14816 92440 14822
rect 92388 14758 92440 14764
rect 89628 14748 89680 14754
rect 89628 14690 89680 14696
rect 85488 14680 85540 14686
rect 85488 14622 85540 14628
rect 85500 3262 85528 14622
rect 87328 8288 87380 8294
rect 87328 8230 87380 8236
rect 84844 3256 84896 3262
rect 84844 3198 84896 3204
rect 84936 3256 84988 3262
rect 84936 3198 84988 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 84948 480 84976 3198
rect 86132 3052 86184 3058
rect 86132 2994 86184 3000
rect 86144 480 86172 2994
rect 87340 480 87368 8230
rect 89640 3262 89668 14690
rect 91008 10600 91060 10606
rect 91008 10542 91060 10548
rect 91020 3482 91048 10542
rect 90928 3454 91048 3482
rect 88524 3256 88576 3262
rect 88524 3198 88576 3204
rect 89628 3256 89680 3262
rect 89628 3198 89680 3204
rect 88536 480 88564 3198
rect 89720 3120 89772 3126
rect 89720 3062 89772 3068
rect 89732 480 89760 3062
rect 90928 480 90956 3454
rect 92400 3346 92428 14758
rect 95148 10668 95200 10674
rect 95148 10610 95200 10616
rect 92124 3318 92428 3346
rect 92124 480 92152 3318
rect 95160 3126 95188 10610
rect 94504 3120 94556 3126
rect 94504 3062 94556 3068
rect 95148 3120 95200 3126
rect 95148 3062 95200 3068
rect 95700 3120 95752 3126
rect 95700 3062 95752 3068
rect 93308 2984 93360 2990
rect 93308 2926 93360 2932
rect 93320 480 93348 2926
rect 94516 480 94544 3062
rect 95712 480 95740 3062
rect 95896 2854 95924 337010
rect 96528 14884 96580 14890
rect 96528 14826 96580 14832
rect 96540 3126 96568 14826
rect 96528 3120 96580 3126
rect 96528 3062 96580 3068
rect 97276 3058 97304 337146
rect 100668 337136 100720 337142
rect 100668 337078 100720 337084
rect 99288 14952 99340 14958
rect 99288 14894 99340 14900
rect 99196 10736 99248 10742
rect 99196 10678 99248 10684
rect 99208 3126 99236 10678
rect 98092 3120 98144 3126
rect 98092 3062 98144 3068
rect 99196 3120 99248 3126
rect 99196 3062 99248 3068
rect 97264 3052 97316 3058
rect 97264 2994 97316 3000
rect 96896 2984 96948 2990
rect 96896 2926 96948 2932
rect 95884 2848 95936 2854
rect 95884 2790 95936 2796
rect 96908 480 96936 2926
rect 98104 480 98132 3062
rect 99300 480 99328 14894
rect 100680 3346 100708 337078
rect 107568 337000 107620 337006
rect 107568 336942 107620 336948
rect 102784 336932 102836 336938
rect 102784 336874 102836 336880
rect 102048 10804 102100 10810
rect 102048 10746 102100 10752
rect 100496 3318 100708 3346
rect 100496 480 100524 3318
rect 102060 3126 102088 10746
rect 102796 3210 102824 336874
rect 107476 15088 107528 15094
rect 107476 15030 107528 15036
rect 103428 15020 103480 15026
rect 103428 14962 103480 14968
rect 102612 3182 102824 3210
rect 101588 3120 101640 3126
rect 101588 3062 101640 3068
rect 102048 3120 102100 3126
rect 102048 3062 102100 3068
rect 101600 480 101628 3062
rect 102612 2854 102640 3182
rect 103440 3126 103468 14962
rect 106188 10872 106240 10878
rect 106188 10814 106240 10820
rect 106200 3126 106228 10814
rect 107488 3126 107516 15030
rect 102784 3120 102836 3126
rect 102784 3062 102836 3068
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 105176 3120 105228 3126
rect 105176 3062 105228 3068
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 106372 3120 106424 3126
rect 106372 3062 106424 3068
rect 107476 3120 107528 3126
rect 107476 3062 107528 3068
rect 102600 2848 102652 2854
rect 102600 2790 102652 2796
rect 102796 480 102824 3062
rect 103980 2916 104032 2922
rect 103980 2858 104032 2864
rect 103992 480 104020 2858
rect 105188 480 105216 3062
rect 106384 480 106412 3062
rect 107580 480 107608 336942
rect 118608 336864 118660 336870
rect 118608 336806 118660 336812
rect 110328 15156 110380 15162
rect 110328 15098 110380 15104
rect 108948 10940 109000 10946
rect 108948 10882 109000 10888
rect 108960 3482 108988 10882
rect 110340 3482 110368 15098
rect 114468 14408 114520 14414
rect 114468 14350 114520 14356
rect 113088 11008 113140 11014
rect 113088 10950 113140 10956
rect 108776 3454 108988 3482
rect 109972 3454 110368 3482
rect 108776 480 108804 3454
rect 109972 480 110000 3454
rect 113100 2990 113128 10950
rect 114480 2990 114508 14350
rect 117228 14340 117280 14346
rect 117228 14282 117280 14288
rect 117136 10260 117188 10266
rect 117136 10202 117188 10208
rect 117148 3618 117176 10202
rect 116964 3590 117176 3618
rect 116964 2990 116992 3590
rect 117240 3482 117268 14282
rect 117148 3454 117268 3482
rect 112352 2984 112404 2990
rect 112352 2926 112404 2932
rect 113088 2984 113140 2990
rect 113088 2926 113140 2932
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 115940 2984 115992 2990
rect 115940 2926 115992 2932
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 111156 2916 111208 2922
rect 111156 2858 111208 2864
rect 111168 480 111196 2858
rect 112364 480 112392 2926
rect 113560 480 113588 2926
rect 114744 2848 114796 2854
rect 114744 2790 114796 2796
rect 114756 480 114784 2790
rect 115952 480 115980 2926
rect 117148 480 117176 3454
rect 118620 3346 118648 336806
rect 125508 336796 125560 336802
rect 125508 336738 125560 336744
rect 121368 14272 121420 14278
rect 121368 14214 121420 14220
rect 119988 10192 120040 10198
rect 119988 10134 120040 10140
rect 118252 3318 118648 3346
rect 118252 480 118280 3318
rect 120000 2990 120028 10134
rect 121380 2990 121408 14214
rect 125416 14204 125468 14210
rect 125416 14146 125468 14152
rect 124128 10124 124180 10130
rect 124128 10066 124180 10072
rect 124140 3482 124168 10066
rect 125428 4214 125456 14146
rect 124220 4208 124272 4214
rect 124220 4150 124272 4156
rect 125416 4208 125468 4214
rect 125416 4150 125468 4156
rect 123036 3454 124168 3482
rect 119436 2984 119488 2990
rect 119436 2926 119488 2932
rect 119988 2984 120040 2990
rect 119988 2926 120040 2932
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 121368 2984 121420 2990
rect 121368 2926 121420 2932
rect 119448 480 119476 2926
rect 120644 480 120672 2926
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 121840 480 121868 2790
rect 123036 480 123064 3454
rect 124232 480 124260 4150
rect 125520 3482 125548 336738
rect 183468 13796 183520 13802
rect 183468 13738 183520 13744
rect 179328 13660 179380 13666
rect 179328 13602 179380 13608
rect 176568 13592 176620 13598
rect 176568 13534 176620 13540
rect 172428 13524 172480 13530
rect 172428 13466 172480 13472
rect 168288 13456 168340 13462
rect 168288 13398 168340 13404
rect 165528 13388 165580 13394
rect 165528 13330 165580 13336
rect 160008 13320 160060 13326
rect 160008 13262 160060 13268
rect 155868 13252 155920 13258
rect 155868 13194 155920 13200
rect 151728 12164 151780 12170
rect 151728 12106 151780 12112
rect 148968 12096 149020 12102
rect 148968 12038 149020 12044
rect 144828 12028 144880 12034
rect 144828 11970 144880 11976
rect 142068 11960 142120 11966
rect 142068 11902 142120 11908
rect 128268 11892 128320 11898
rect 128268 11834 128320 11840
rect 126888 11824 126940 11830
rect 126888 11766 126940 11772
rect 126900 3482 126928 11766
rect 128280 3482 128308 11834
rect 139676 9376 139728 9382
rect 139676 9318 139728 9324
rect 136088 9308 136140 9314
rect 136088 9250 136140 9256
rect 132590 8936 132646 8945
rect 132590 8871 132646 8880
rect 129002 7576 129058 7585
rect 129002 7511 129058 7520
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 127820 3454 128308 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3454
rect 129016 480 129044 7511
rect 131396 6656 131448 6662
rect 131396 6598 131448 6604
rect 130200 5364 130252 5370
rect 130200 5306 130252 5312
rect 130212 480 130240 5306
rect 131408 480 131436 6598
rect 132604 480 132632 8871
rect 134892 7540 134944 7546
rect 134892 7482 134944 7488
rect 133788 5432 133840 5438
rect 133788 5374 133840 5380
rect 133800 480 133828 5374
rect 134904 480 134932 7482
rect 136100 480 136128 9250
rect 138480 7472 138532 7478
rect 138480 7414 138532 7420
rect 137284 5500 137336 5506
rect 137284 5442 137336 5448
rect 137296 480 137324 5442
rect 138492 480 138520 7414
rect 139688 480 139716 9318
rect 141976 7404 142028 7410
rect 141976 7346 142028 7352
rect 140872 4208 140924 4214
rect 140872 4150 140924 4156
rect 140884 480 140912 4150
rect 141988 3482 142016 7346
rect 142080 4214 142108 11902
rect 143448 10056 143500 10062
rect 143448 9998 143500 10004
rect 142068 4208 142120 4214
rect 142068 4150 142120 4156
rect 143460 3482 143488 9998
rect 144840 3482 144868 11970
rect 147588 9988 147640 9994
rect 147588 9930 147640 9936
rect 145656 7336 145708 7342
rect 145656 7278 145708 7284
rect 141988 3454 142108 3482
rect 142080 480 142108 3454
rect 143276 3454 143488 3482
rect 144472 3454 144868 3482
rect 143276 480 143304 3454
rect 144472 480 144500 3454
rect 145668 480 145696 7278
rect 147600 3482 147628 9930
rect 148980 3482 149008 12038
rect 151636 9920 151688 9926
rect 151636 9862 151688 9868
rect 149244 7268 149296 7274
rect 149244 7210 149296 7216
rect 146864 3454 147628 3482
rect 148060 3454 149008 3482
rect 146864 480 146892 3454
rect 148060 480 148088 3454
rect 149256 480 149284 7210
rect 151648 4214 151676 9862
rect 150440 4208 150492 4214
rect 150440 4150 150492 4156
rect 151636 4208 151688 4214
rect 151636 4150 151688 4156
rect 150452 480 150480 4150
rect 151740 3482 151768 12106
rect 154488 9852 154540 9858
rect 154488 9794 154540 9800
rect 152740 7200 152792 7206
rect 152740 7142 152792 7148
rect 151556 3454 151768 3482
rect 151556 480 151584 3454
rect 152752 480 152780 7142
rect 154500 3482 154528 9794
rect 155880 3482 155908 13194
rect 158628 9784 158680 9790
rect 158628 9726 158680 9732
rect 156328 7132 156380 7138
rect 156328 7074 156380 7080
rect 153948 3454 154528 3482
rect 155144 3454 155908 3482
rect 153948 480 153976 3454
rect 155144 480 155172 3454
rect 156340 480 156368 7074
rect 158640 3482 158668 9726
rect 159916 7064 159968 7070
rect 159916 7006 159968 7012
rect 158720 4208 158772 4214
rect 158720 4150 158772 4156
rect 157536 3454 158668 3482
rect 157536 480 157564 3454
rect 158732 480 158760 4150
rect 159928 480 159956 7006
rect 160020 4214 160048 13262
rect 162768 12232 162820 12238
rect 162768 12174 162820 12180
rect 161388 9716 161440 9722
rect 161388 9658 161440 9664
rect 160008 4208 160060 4214
rect 160008 4150 160060 4156
rect 161400 3482 161428 9658
rect 161124 3454 161428 3482
rect 161124 480 161152 3454
rect 162780 626 162808 12174
rect 163504 6724 163556 6730
rect 163504 6666 163556 6672
rect 162320 598 162808 626
rect 162320 480 162348 598
rect 163516 480 163544 6666
rect 165540 610 165568 13330
rect 166908 12300 166960 12306
rect 166908 12242 166960 12248
rect 166920 610 166948 12242
rect 167092 6792 167144 6798
rect 167092 6734 167144 6740
rect 164700 604 164752 610
rect 164700 546 164752 552
rect 165528 604 165580 610
rect 165528 546 165580 552
rect 165896 604 165948 610
rect 165896 546 165948 552
rect 166908 604 166960 610
rect 166908 546 166960 552
rect 164712 480 164740 546
rect 165908 480 165936 546
rect 167104 480 167132 6734
rect 168300 626 168328 13398
rect 169668 12368 169720 12374
rect 169668 12310 169720 12316
rect 168208 598 168328 626
rect 169680 610 169708 12310
rect 170588 6860 170640 6866
rect 170588 6802 170640 6808
rect 169392 604 169444 610
rect 168208 480 168236 598
rect 169392 546 169444 552
rect 169668 604 169720 610
rect 169668 546 169720 552
rect 169404 480 169432 546
rect 170600 480 170628 6802
rect 172440 3346 172468 13466
rect 173808 12436 173860 12442
rect 173808 12378 173860 12384
rect 173820 3346 173848 12378
rect 176476 11688 176528 11694
rect 176476 11630 176528 11636
rect 174176 6112 174228 6118
rect 174176 6054 174228 6060
rect 171796 3318 172468 3346
rect 172992 3318 173848 3346
rect 171796 480 171824 3318
rect 172992 480 173020 3318
rect 174188 480 174216 6054
rect 175372 4208 175424 4214
rect 175372 4150 175424 4156
rect 175384 480 175412 4150
rect 176488 3482 176516 11630
rect 176580 4214 176608 13534
rect 177764 6044 177816 6050
rect 177764 5986 177816 5992
rect 176568 4208 176620 4214
rect 176568 4150 176620 4156
rect 176488 3454 176608 3482
rect 176580 480 176608 3454
rect 177776 480 177804 5986
rect 179340 3346 179368 13602
rect 180708 11620 180760 11626
rect 180708 11562 180760 11568
rect 180720 3346 180748 11562
rect 181352 5976 181404 5982
rect 181352 5918 181404 5924
rect 178972 3318 179368 3346
rect 180168 3318 180748 3346
rect 178972 480 179000 3318
rect 180168 480 180196 3318
rect 181364 480 181392 5918
rect 183480 610 183508 13738
rect 186228 13728 186280 13734
rect 186228 13670 186280 13676
rect 184848 11552 184900 11558
rect 184848 11494 184900 11500
rect 184860 6066 184888 11494
rect 184768 6038 184888 6066
rect 184768 610 184796 6038
rect 184848 5908 184900 5914
rect 184848 5850 184900 5856
rect 182548 604 182600 610
rect 182548 546 182600 552
rect 183468 604 183520 610
rect 183468 546 183520 552
rect 183744 604 183796 610
rect 183744 546 183796 552
rect 184756 604 184808 610
rect 184756 546 184808 552
rect 182560 480 182588 546
rect 183756 480 183784 546
rect 184860 480 184888 5850
rect 186240 626 186268 13670
rect 190368 13048 190420 13054
rect 190368 12990 190420 12996
rect 187608 11484 187660 11490
rect 187608 11426 187660 11432
rect 186056 598 186268 626
rect 187620 610 187648 11426
rect 188436 5840 188488 5846
rect 188436 5782 188488 5788
rect 187240 604 187292 610
rect 186056 480 186084 598
rect 187240 546 187292 552
rect 187608 604 187660 610
rect 187608 546 187660 552
rect 187252 480 187280 546
rect 188448 480 188476 5782
rect 190380 610 190408 12990
rect 206928 12980 206980 12986
rect 206928 12922 206980 12928
rect 191748 11416 191800 11422
rect 191748 11358 191800 11364
rect 191760 3346 191788 11358
rect 194508 11348 194560 11354
rect 194508 11290 194560 11296
rect 193220 9444 193272 9450
rect 193220 9386 193272 9392
rect 192024 5772 192076 5778
rect 192024 5714 192076 5720
rect 190840 3318 191788 3346
rect 189632 604 189684 610
rect 189632 546 189684 552
rect 190368 604 190420 610
rect 190368 546 190420 552
rect 189644 480 189672 546
rect 190840 480 190868 3318
rect 192036 480 192064 5714
rect 193232 480 193260 9386
rect 194520 3482 194548 11290
rect 198648 11280 198700 11286
rect 198648 11222 198700 11228
rect 196808 9512 196860 9518
rect 196808 9454 196860 9460
rect 195612 5704 195664 5710
rect 195612 5646 195664 5652
rect 194428 3454 194548 3482
rect 194428 480 194456 3454
rect 195624 480 195652 5646
rect 196820 480 196848 9454
rect 198660 3346 198688 11222
rect 203892 9648 203944 9654
rect 203892 9590 203944 9596
rect 200396 9580 200448 9586
rect 200396 9522 200448 9528
rect 199200 5568 199252 5574
rect 199200 5510 199252 5516
rect 198016 3318 198688 3346
rect 198016 480 198044 3318
rect 199212 480 199240 5510
rect 200408 480 200436 9522
rect 202696 5636 202748 5642
rect 202696 5578 202748 5584
rect 201500 4412 201552 4418
rect 201500 4354 201552 4360
rect 201512 480 201540 4354
rect 202708 480 202736 5578
rect 203904 480 203932 9590
rect 205088 4344 205140 4350
rect 205088 4286 205140 4292
rect 205100 480 205128 4286
rect 206940 3346 206968 12922
rect 211068 12912 211120 12918
rect 211068 12854 211120 12860
rect 207480 8900 207532 8906
rect 207480 8842 207532 8848
rect 206296 3318 206968 3346
rect 206296 480 206324 3318
rect 207492 480 207520 8842
rect 210976 8832 211028 8838
rect 210976 8774 211028 8780
rect 208674 4856 208730 4865
rect 208674 4791 208730 4800
rect 208688 480 208716 4791
rect 209872 4208 209924 4214
rect 209872 4150 209924 4156
rect 209884 480 209912 4150
rect 210988 3482 211016 8774
rect 211080 4214 211108 12854
rect 213828 12844 213880 12850
rect 213828 12786 213880 12792
rect 212264 4752 212316 4758
rect 212264 4694 212316 4700
rect 211068 4208 211120 4214
rect 211068 4150 211120 4156
rect 210988 3454 211108 3482
rect 211080 480 211108 3454
rect 212276 480 212304 4694
rect 213840 3346 213868 12786
rect 217968 12776 218020 12782
rect 217968 12718 218020 12724
rect 214656 8764 214708 8770
rect 214656 8706 214708 8712
rect 213472 3318 213868 3346
rect 213472 480 213500 3318
rect 214668 480 214696 8706
rect 215852 4684 215904 4690
rect 215852 4626 215904 4632
rect 215864 480 215892 4626
rect 217980 3346 218008 12718
rect 220728 12708 220780 12714
rect 220728 12650 220780 12656
rect 218152 8696 218204 8702
rect 218152 8638 218204 8644
rect 217060 3318 218008 3346
rect 217060 480 217088 3318
rect 218164 480 218192 8638
rect 219348 4616 219400 4622
rect 219348 4558 219400 4564
rect 219360 480 219388 4558
rect 220740 3346 220768 12650
rect 224868 12640 224920 12646
rect 224868 12582 224920 12588
rect 221740 8628 221792 8634
rect 221740 8570 221792 8576
rect 220556 3318 220768 3346
rect 220556 480 220584 3318
rect 221752 480 221780 8570
rect 222936 4548 222988 4554
rect 222936 4490 222988 4496
rect 222948 480 222976 4490
rect 224880 3346 224908 12582
rect 229008 12572 229060 12578
rect 229008 12514 229060 12520
rect 225328 8560 225380 8566
rect 225328 8502 225380 8508
rect 224144 3318 224908 3346
rect 224144 480 224172 3318
rect 225340 480 225368 8502
rect 228916 8492 228968 8498
rect 228916 8434 228968 8440
rect 227720 7608 227772 7614
rect 227720 7550 227772 7556
rect 226524 4480 226576 4486
rect 226524 4422 226576 4428
rect 226536 480 226564 4422
rect 227732 480 227760 7550
rect 228928 480 228956 8434
rect 229020 7614 229048 12514
rect 229008 7608 229060 7614
rect 229008 7550 229060 7556
rect 229112 4962 229140 340054
rect 229192 337272 229244 337278
rect 229190 337240 229192 337249
rect 229244 337240 229246 337249
rect 229190 337175 229246 337184
rect 229100 4956 229152 4962
rect 229100 4898 229152 4904
rect 230112 4888 230164 4894
rect 230112 4830 230164 4836
rect 230124 480 230152 4830
rect 230492 4282 230520 340068
rect 230584 340054 230966 340082
rect 230584 4826 230612 340054
rect 231044 337770 231072 340190
rect 230768 337742 231072 337770
rect 230768 321570 230796 337742
rect 231964 337385 231992 340068
rect 232056 340054 232438 340082
rect 231950 337376 232006 337385
rect 231950 337311 232006 337320
rect 230756 321564 230808 321570
rect 230756 321506 230808 321512
rect 230940 321564 230992 321570
rect 230940 321506 230992 321512
rect 230952 318782 230980 321506
rect 230940 318776 230992 318782
rect 230940 318718 230992 318724
rect 230848 309188 230900 309194
rect 230848 309130 230900 309136
rect 230860 205578 230888 309130
rect 230768 205550 230888 205578
rect 230768 202881 230796 205550
rect 230754 202872 230810 202881
rect 230754 202807 230810 202816
rect 231030 202872 231086 202881
rect 231030 202807 231086 202816
rect 231044 193254 231072 202807
rect 230848 193248 230900 193254
rect 230848 193190 230900 193196
rect 231032 193248 231084 193254
rect 231032 193190 231084 193196
rect 230860 186266 230888 193190
rect 230768 186238 230888 186266
rect 230768 183569 230796 186238
rect 230754 183560 230810 183569
rect 230754 183495 230810 183504
rect 231030 183560 231086 183569
rect 231030 183495 231086 183504
rect 231044 173942 231072 183495
rect 230848 173936 230900 173942
rect 230848 173878 230900 173884
rect 231032 173936 231084 173942
rect 231032 173878 231084 173884
rect 230860 166954 230888 173878
rect 230768 166926 230888 166954
rect 230768 162858 230796 166926
rect 230664 162852 230716 162858
rect 230664 162794 230716 162800
rect 230756 162852 230808 162858
rect 230756 162794 230808 162800
rect 230676 153241 230704 162794
rect 230662 153232 230718 153241
rect 230662 153167 230718 153176
rect 230846 153232 230902 153241
rect 230846 153167 230902 153176
rect 230860 143546 230888 153167
rect 230848 143540 230900 143546
rect 230848 143482 230900 143488
rect 230848 133952 230900 133958
rect 230848 133894 230900 133900
rect 230860 60654 230888 133894
rect 230848 60648 230900 60654
rect 230848 60590 230900 60596
rect 230756 48340 230808 48346
rect 230756 48282 230808 48288
rect 230768 38758 230796 48282
rect 230756 38752 230808 38758
rect 230756 38694 230808 38700
rect 230756 37324 230808 37330
rect 230756 37266 230808 37272
rect 230768 27606 230796 37266
rect 230756 27600 230808 27606
rect 230756 27542 230808 27548
rect 230756 18012 230808 18018
rect 230756 17954 230808 17960
rect 230768 12510 230796 17954
rect 230756 12504 230808 12510
rect 230756 12446 230808 12452
rect 230664 11212 230716 11218
rect 230664 11154 230716 11160
rect 230676 7682 230704 11154
rect 230664 7676 230716 7682
rect 230664 7618 230716 7624
rect 231308 7608 231360 7614
rect 231308 7550 231360 7556
rect 230572 4820 230624 4826
rect 230572 4762 230624 4768
rect 230480 4276 230532 4282
rect 230480 4218 230532 4224
rect 231320 480 231348 7550
rect 232056 3369 232084 340054
rect 232516 337770 232544 340190
rect 232240 337742 232544 337770
rect 232240 321570 232268 337742
rect 232228 321564 232280 321570
rect 232228 321506 232280 321512
rect 232412 321564 232464 321570
rect 232412 321506 232464 321512
rect 232424 311982 232452 321506
rect 232412 311976 232464 311982
rect 232412 311918 232464 311924
rect 232320 311840 232372 311846
rect 232320 311782 232372 311788
rect 232332 205578 232360 311782
rect 232240 205550 232360 205578
rect 232240 196042 232268 205550
rect 232228 196036 232280 196042
rect 232228 195978 232280 195984
rect 232320 195968 232372 195974
rect 232320 195910 232372 195916
rect 232332 186266 232360 195910
rect 232240 186238 232360 186266
rect 232240 176730 232268 186238
rect 232228 176724 232280 176730
rect 232228 176666 232280 176672
rect 232320 176656 232372 176662
rect 232320 176598 232372 176604
rect 232332 166954 232360 176598
rect 232240 166926 232360 166954
rect 232240 159338 232268 166926
rect 232240 159310 232452 159338
rect 232424 154562 232452 159310
rect 232412 154556 232464 154562
rect 232412 154498 232464 154504
rect 232320 145036 232372 145042
rect 232320 144978 232372 144984
rect 232332 143546 232360 144978
rect 232320 143540 232372 143546
rect 232320 143482 232372 143488
rect 232320 133952 232372 133958
rect 232320 133894 232372 133900
rect 232332 124166 232360 133894
rect 232320 124160 232372 124166
rect 232320 124102 232372 124108
rect 232320 114572 232372 114578
rect 232320 114514 232372 114520
rect 232332 104854 232360 114514
rect 232320 104848 232372 104854
rect 232320 104790 232372 104796
rect 232320 95260 232372 95266
rect 232320 95202 232372 95208
rect 232332 85542 232360 95202
rect 232320 85536 232372 85542
rect 232320 85478 232372 85484
rect 232320 75948 232372 75954
rect 232320 75890 232372 75896
rect 232332 66230 232360 75890
rect 232320 66224 232372 66230
rect 232320 66166 232372 66172
rect 232320 56636 232372 56642
rect 232320 56578 232372 56584
rect 232332 51134 232360 56578
rect 232320 51128 232372 51134
rect 232320 51070 232372 51076
rect 232228 51060 232280 51066
rect 232228 51002 232280 51008
rect 232240 48226 232268 51002
rect 232240 48198 232360 48226
rect 232332 37398 232360 48198
rect 232320 37392 232372 37398
rect 232320 37334 232372 37340
rect 232228 37324 232280 37330
rect 232228 37266 232280 37272
rect 232240 37194 232268 37266
rect 232228 37188 232280 37194
rect 232228 37130 232280 37136
rect 232320 27668 232372 27674
rect 232320 27610 232372 27616
rect 232332 27554 232360 27610
rect 232332 27526 232452 27554
rect 232424 22778 232452 27526
rect 232412 22772 232464 22778
rect 232412 22714 232464 22720
rect 232136 14136 232188 14142
rect 232136 14078 232188 14084
rect 232148 5030 232176 14078
rect 232504 8424 232556 8430
rect 232504 8366 232556 8372
rect 232136 5024 232188 5030
rect 232136 4966 232188 4972
rect 232042 3360 232098 3369
rect 232042 3295 232098 3304
rect 232516 480 232544 8366
rect 233436 7002 233464 340068
rect 233528 340054 233910 340082
rect 233528 337414 233556 340054
rect 234356 337482 234384 340068
rect 234724 340054 234922 340082
rect 235092 340054 235382 340082
rect 235460 340054 235842 340082
rect 236394 340054 236500 340082
rect 234344 337476 234396 337482
rect 234344 337418 234396 337424
rect 233516 337408 233568 337414
rect 233516 337350 233568 337356
rect 233884 337408 233936 337414
rect 233884 337350 233936 337356
rect 233896 9110 233924 337350
rect 234620 337272 234672 337278
rect 234618 337240 234620 337249
rect 234672 337240 234674 337249
rect 234618 337175 234674 337184
rect 233884 9104 233936 9110
rect 233884 9046 233936 9052
rect 233424 6996 233476 7002
rect 233424 6938 233476 6944
rect 234724 5098 234752 340054
rect 235092 335730 235120 340054
rect 234816 335702 235120 335730
rect 234816 8974 234844 335702
rect 235460 335594 235488 340054
rect 236184 335708 236236 335714
rect 236184 335650 236236 335656
rect 235092 335566 235488 335594
rect 236092 335640 236144 335646
rect 236092 335582 236144 335588
rect 235092 318782 235120 335566
rect 235080 318776 235132 318782
rect 235080 318718 235132 318724
rect 235080 311840 235132 311846
rect 235080 311782 235132 311788
rect 235092 299470 235120 311782
rect 235080 299464 235132 299470
rect 235080 299406 235132 299412
rect 235080 289876 235132 289882
rect 235080 289818 235132 289824
rect 235092 280158 235120 289818
rect 235080 280152 235132 280158
rect 235080 280094 235132 280100
rect 235080 270564 235132 270570
rect 235080 270506 235132 270512
rect 235092 260846 235120 270506
rect 235080 260840 235132 260846
rect 235080 260782 235132 260788
rect 235080 251252 235132 251258
rect 235080 251194 235132 251200
rect 235092 241505 235120 251194
rect 234894 241496 234950 241505
rect 234894 241431 234950 241440
rect 235078 241496 235134 241505
rect 235078 241431 235134 241440
rect 234908 231878 234936 241431
rect 234896 231872 234948 231878
rect 234896 231814 234948 231820
rect 235080 231872 235132 231878
rect 235080 231814 235132 231820
rect 235092 222193 235120 231814
rect 234894 222184 234950 222193
rect 234894 222119 234950 222128
rect 235078 222184 235134 222193
rect 235078 222119 235134 222128
rect 234908 212566 234936 222119
rect 234896 212560 234948 212566
rect 234896 212502 234948 212508
rect 235080 212560 235132 212566
rect 235080 212502 235132 212508
rect 235092 195974 235120 212502
rect 235080 195968 235132 195974
rect 235080 195910 235132 195916
rect 235080 195832 235132 195838
rect 235080 195774 235132 195780
rect 235092 176662 235120 195774
rect 235080 176656 235132 176662
rect 235080 176598 235132 176604
rect 235080 176520 235132 176526
rect 235080 176462 235132 176468
rect 235092 164218 235120 176462
rect 235080 164212 235132 164218
rect 235080 164154 235132 164160
rect 235080 154624 235132 154630
rect 235080 154566 235132 154572
rect 235092 147762 235120 154566
rect 235080 147756 235132 147762
rect 235080 147698 235132 147704
rect 235080 147620 235132 147626
rect 235080 147562 235132 147568
rect 235092 138038 235120 147562
rect 235080 138032 235132 138038
rect 235080 137974 235132 137980
rect 235080 137896 235132 137902
rect 235080 137838 235132 137844
rect 235092 125594 235120 137838
rect 235080 125588 235132 125594
rect 235080 125530 235132 125536
rect 235080 116000 235132 116006
rect 235080 115942 235132 115948
rect 235092 106282 235120 115942
rect 235080 106276 235132 106282
rect 235080 106218 235132 106224
rect 235080 96688 235132 96694
rect 235080 96630 235132 96636
rect 235092 86970 235120 96630
rect 235080 86964 235132 86970
rect 235080 86906 235132 86912
rect 235080 77308 235132 77314
rect 235080 77250 235132 77256
rect 235092 67590 235120 77250
rect 235080 67584 235132 67590
rect 235080 67526 235132 67532
rect 235080 62756 235132 62762
rect 235080 62698 235132 62704
rect 235092 41426 235120 62698
rect 235000 41398 235120 41426
rect 235000 41290 235028 41398
rect 235000 41262 235120 41290
rect 235092 22114 235120 41262
rect 235000 22086 235120 22114
rect 235000 12322 235028 22086
rect 234908 12294 235028 12322
rect 234804 8968 234856 8974
rect 234804 8910 234856 8916
rect 234804 7676 234856 7682
rect 234804 7618 234856 7624
rect 234712 5092 234764 5098
rect 234712 5034 234764 5040
rect 233700 4820 233752 4826
rect 233700 4762 233752 4768
rect 233712 480 233740 4762
rect 234816 480 234844 7618
rect 234908 3534 234936 12294
rect 236000 8968 236052 8974
rect 236000 8910 236052 8916
rect 234896 3528 234948 3534
rect 234896 3470 234948 3476
rect 236012 480 236040 8910
rect 236104 5166 236132 335582
rect 236196 9042 236224 335650
rect 236472 321586 236500 340054
rect 236564 340054 236854 340082
rect 237024 340054 237314 340082
rect 236564 335646 236592 340054
rect 237024 335714 237052 340054
rect 237852 337482 237880 340068
rect 238312 337754 238340 340068
rect 238786 340054 238892 340082
rect 238300 337748 238352 337754
rect 238300 337690 238352 337696
rect 237840 337476 237892 337482
rect 237840 337418 237892 337424
rect 237012 335708 237064 335714
rect 237012 335650 237064 335656
rect 236552 335640 236604 335646
rect 236552 335582 236604 335588
rect 236288 321558 236500 321586
rect 236288 318782 236316 321558
rect 236276 318776 236328 318782
rect 236276 318718 236328 318724
rect 236276 309188 236328 309194
rect 236276 309130 236328 309136
rect 236288 299470 236316 309130
rect 236276 299464 236328 299470
rect 236276 299406 236328 299412
rect 236276 289876 236328 289882
rect 236276 289818 236328 289824
rect 236288 280158 236316 289818
rect 236276 280152 236328 280158
rect 236276 280094 236328 280100
rect 236276 270564 236328 270570
rect 236276 270506 236328 270512
rect 236288 260846 236316 270506
rect 236276 260840 236328 260846
rect 236276 260782 236328 260788
rect 236276 251252 236328 251258
rect 236276 251194 236328 251200
rect 236288 241505 236316 251194
rect 236274 241496 236330 241505
rect 236274 241431 236330 241440
rect 236458 241496 236514 241505
rect 236458 241431 236514 241440
rect 236472 231878 236500 241431
rect 236276 231872 236328 231878
rect 236276 231814 236328 231820
rect 236460 231872 236512 231878
rect 236460 231814 236512 231820
rect 236288 222193 236316 231814
rect 236274 222184 236330 222193
rect 236274 222119 236330 222128
rect 236458 222184 236514 222193
rect 236458 222119 236514 222128
rect 236472 212566 236500 222119
rect 236276 212560 236328 212566
rect 236276 212502 236328 212508
rect 236460 212560 236512 212566
rect 236460 212502 236512 212508
rect 236288 202881 236316 212502
rect 236274 202872 236330 202881
rect 236274 202807 236330 202816
rect 236458 202872 236514 202881
rect 236458 202807 236514 202816
rect 236472 193254 236500 202807
rect 236276 193248 236328 193254
rect 236276 193190 236328 193196
rect 236460 193248 236512 193254
rect 236460 193190 236512 193196
rect 236288 183569 236316 193190
rect 236274 183560 236330 183569
rect 236274 183495 236330 183504
rect 236458 183560 236514 183569
rect 236458 183495 236514 183504
rect 236472 173942 236500 183495
rect 236276 173936 236328 173942
rect 236276 173878 236328 173884
rect 236460 173936 236512 173942
rect 236460 173878 236512 173884
rect 236288 164218 236316 173878
rect 236276 164212 236328 164218
rect 236276 164154 236328 164160
rect 236460 164212 236512 164218
rect 236460 164154 236512 164160
rect 236472 154601 236500 164154
rect 236274 154592 236330 154601
rect 236274 154527 236330 154536
rect 236458 154592 236514 154601
rect 236458 154527 236514 154536
rect 236288 147642 236316 154527
rect 236288 147614 236500 147642
rect 236472 135289 236500 147614
rect 236274 135280 236330 135289
rect 236274 135215 236330 135224
rect 236458 135280 236514 135289
rect 236458 135215 236514 135224
rect 236288 125594 236316 135215
rect 236276 125588 236328 125594
rect 236276 125530 236328 125536
rect 236460 125588 236512 125594
rect 236460 125530 236512 125536
rect 236472 115977 236500 125530
rect 236274 115968 236330 115977
rect 236274 115903 236330 115912
rect 236458 115968 236514 115977
rect 236458 115903 236514 115912
rect 236288 106282 236316 115903
rect 236276 106276 236328 106282
rect 236276 106218 236328 106224
rect 236460 106276 236512 106282
rect 236460 106218 236512 106224
rect 236472 96665 236500 106218
rect 236274 96656 236330 96665
rect 236274 96591 236330 96600
rect 236458 96656 236514 96665
rect 236458 96591 236514 96600
rect 236288 86970 236316 96591
rect 236276 86964 236328 86970
rect 236276 86906 236328 86912
rect 236276 77308 236328 77314
rect 236276 77250 236328 77256
rect 236288 67590 236316 77250
rect 236276 67584 236328 67590
rect 236276 67526 236328 67532
rect 236276 57996 236328 58002
rect 236276 57938 236328 57944
rect 236288 48278 236316 57938
rect 236276 48272 236328 48278
rect 236276 48214 236328 48220
rect 236276 38684 236328 38690
rect 236276 38626 236328 38632
rect 236288 31634 236316 38626
rect 236288 31606 236408 31634
rect 236380 12458 236408 31606
rect 236380 12430 236500 12458
rect 236472 12322 236500 12430
rect 236288 12294 236500 12322
rect 236184 9036 236236 9042
rect 236184 8978 236236 8984
rect 236092 5160 236144 5166
rect 236092 5102 236144 5108
rect 236288 3466 236316 12294
rect 238864 7750 238892 340054
rect 238956 340054 239338 340082
rect 239508 340054 239798 340082
rect 240258 340054 240364 340082
rect 238956 11762 238984 340054
rect 239508 331242 239536 340054
rect 239140 331214 239536 331242
rect 239140 311710 239168 331214
rect 239128 311704 239180 311710
rect 239128 311646 239180 311652
rect 239128 311568 239180 311574
rect 239128 311510 239180 311516
rect 239140 292534 239168 311510
rect 239128 292528 239180 292534
rect 239128 292470 239180 292476
rect 239128 292392 239180 292398
rect 239128 292334 239180 292340
rect 239140 273222 239168 292334
rect 239128 273216 239180 273222
rect 239128 273158 239180 273164
rect 239128 273080 239180 273086
rect 239128 273022 239180 273028
rect 239140 253910 239168 273022
rect 239128 253904 239180 253910
rect 239128 253846 239180 253852
rect 239128 253768 239180 253774
rect 239128 253710 239180 253716
rect 239140 234598 239168 253710
rect 239128 234592 239180 234598
rect 239128 234534 239180 234540
rect 239128 234456 239180 234462
rect 239128 234398 239180 234404
rect 239140 215286 239168 234398
rect 239128 215280 239180 215286
rect 239128 215222 239180 215228
rect 239128 215144 239180 215150
rect 239128 215086 239180 215092
rect 239140 176526 239168 215086
rect 239128 176520 239180 176526
rect 239128 176462 239180 176468
rect 239128 176384 239180 176390
rect 239128 176326 239180 176332
rect 239140 128466 239168 176326
rect 239048 128438 239168 128466
rect 239048 128330 239076 128438
rect 239048 128302 239168 128330
rect 239140 99498 239168 128302
rect 239048 99470 239168 99498
rect 239048 99362 239076 99470
rect 239048 99334 239168 99362
rect 239140 60738 239168 99334
rect 239048 60710 239168 60738
rect 239048 60602 239076 60710
rect 239048 60574 239168 60602
rect 239140 41426 239168 60574
rect 239048 41398 239168 41426
rect 239048 41290 239076 41398
rect 239048 41262 239168 41290
rect 239140 12458 239168 41262
rect 239140 12430 239260 12458
rect 239232 12322 239260 12430
rect 239048 12294 239260 12322
rect 238944 11756 238996 11762
rect 238944 11698 238996 11704
rect 238852 7744 238904 7750
rect 238852 7686 238904 7692
rect 238392 6996 238444 7002
rect 238392 6938 238444 6944
rect 238114 5400 238170 5409
rect 238114 5335 238170 5344
rect 237196 4956 237248 4962
rect 237196 4898 237248 4904
rect 236276 3460 236328 3466
rect 236276 3402 236328 3408
rect 237208 480 237236 4898
rect 238128 3874 238156 5335
rect 238116 3868 238168 3874
rect 238116 3810 238168 3816
rect 238404 480 238432 6938
rect 239048 3670 239076 12294
rect 239588 9036 239640 9042
rect 239588 8978 239640 8984
rect 239036 3664 239088 3670
rect 239036 3606 239088 3612
rect 239600 480 239628 8978
rect 240336 3602 240364 340054
rect 240428 340054 240810 340082
rect 240428 7818 240456 340054
rect 241256 337414 241284 340068
rect 241716 337618 241744 340068
rect 241808 340054 242282 340082
rect 242360 340054 242742 340082
rect 243096 340054 243202 340082
rect 243464 340054 243754 340082
rect 241704 337612 241756 337618
rect 241704 337554 241756 337560
rect 241244 337408 241296 337414
rect 241244 337350 241296 337356
rect 241612 335640 241664 335646
rect 241612 335582 241664 335588
rect 241624 13122 241652 335582
rect 241612 13116 241664 13122
rect 241612 13058 241664 13064
rect 241808 7886 241836 340054
rect 242360 335646 242388 340054
rect 242348 335640 242400 335646
rect 242348 335582 242400 335588
rect 242992 332104 243044 332110
rect 242992 332046 243044 332052
rect 243004 7954 243032 332046
rect 242992 7948 243044 7954
rect 242992 7890 243044 7896
rect 241796 7880 241848 7886
rect 241796 7822 241848 7828
rect 240416 7812 240468 7818
rect 240416 7754 240468 7760
rect 241980 7744 242032 7750
rect 241980 7686 242032 7692
rect 240784 5024 240836 5030
rect 240784 4966 240836 4972
rect 240324 3596 240376 3602
rect 240324 3538 240376 3544
rect 240796 480 240824 4966
rect 241992 480 242020 7686
rect 243096 3738 243124 340054
rect 243464 332110 243492 340054
rect 244200 337822 244228 340068
rect 244188 337816 244240 337822
rect 244188 337758 244240 337764
rect 244660 337686 244688 340068
rect 244648 337680 244700 337686
rect 244648 337622 244700 337628
rect 243452 332104 243504 332110
rect 243452 332046 243504 332052
rect 244752 331242 244780 340190
rect 244476 331214 244780 331242
rect 244476 317506 244504 331214
rect 244384 317478 244504 317506
rect 244384 311982 244412 317478
rect 244372 311976 244424 311982
rect 244372 311918 244424 311924
rect 244464 311772 244516 311778
rect 244464 311714 244516 311720
rect 244476 288454 244504 311714
rect 244464 288448 244516 288454
rect 244464 288390 244516 288396
rect 244556 288448 244608 288454
rect 244556 288390 244608 288396
rect 244568 270552 244596 288390
rect 244476 270524 244596 270552
rect 244476 259486 244504 270524
rect 244372 259480 244424 259486
rect 244372 259422 244424 259428
rect 244464 259480 244516 259486
rect 244464 259422 244516 259428
rect 244384 249801 244412 259422
rect 244370 249792 244426 249801
rect 244370 249727 244426 249736
rect 244554 249792 244610 249801
rect 244554 249727 244610 249736
rect 244384 240174 244412 240205
rect 244568 240174 244596 249727
rect 244372 240168 244424 240174
rect 244556 240168 244608 240174
rect 244424 240116 244504 240122
rect 244372 240110 244504 240116
rect 244556 240110 244608 240116
rect 244384 240094 244504 240110
rect 244476 234666 244504 240094
rect 244464 234660 244516 234666
rect 244464 234602 244516 234608
rect 244372 234592 244424 234598
rect 244372 234534 244424 234540
rect 244384 220794 244412 234534
rect 244372 220788 244424 220794
rect 244372 220730 244424 220736
rect 244464 212492 244516 212498
rect 244464 212434 244516 212440
rect 244476 211154 244504 212434
rect 244476 211126 244596 211154
rect 244568 202910 244596 211126
rect 244372 202904 244424 202910
rect 244372 202846 244424 202852
rect 244556 202904 244608 202910
rect 244556 202846 244608 202852
rect 244384 193254 244412 202846
rect 244372 193248 244424 193254
rect 244372 193190 244424 193196
rect 244464 193248 244516 193254
rect 244464 193190 244516 193196
rect 244476 185586 244504 193190
rect 245384 189100 245436 189106
rect 245384 189042 245436 189048
rect 244476 185558 244596 185586
rect 244568 182050 244596 185558
rect 244384 182022 244596 182050
rect 244384 171086 244412 182022
rect 245396 180674 245424 189042
rect 245672 180878 245700 340068
rect 245764 340054 246146 340082
rect 245764 180946 245792 340054
rect 246224 334642 246252 340190
rect 247144 337958 247172 340068
rect 247132 337952 247184 337958
rect 247132 337894 247184 337900
rect 247604 337890 247632 340068
rect 247788 340054 248170 340082
rect 247592 337884 247644 337890
rect 247592 337826 247644 337832
rect 247788 337498 247816 340054
rect 245948 334614 246252 334642
rect 247144 337470 247816 337498
rect 245948 317506 245976 334614
rect 247144 331106 247172 337470
rect 248616 337414 248644 340068
rect 248708 340054 249090 340082
rect 249168 340054 249550 340082
rect 249904 340054 250102 340082
rect 247684 337408 247736 337414
rect 247684 337350 247736 337356
rect 248604 337408 248656 337414
rect 248604 337350 248656 337356
rect 247144 331078 247264 331106
rect 245856 317478 245976 317506
rect 245856 311982 245884 317478
rect 247236 315874 247264 331078
rect 247236 315846 247356 315874
rect 245844 311976 245896 311982
rect 245844 311918 245896 311924
rect 245936 311772 245988 311778
rect 245936 311714 245988 311720
rect 245948 278769 245976 311714
rect 247328 298178 247356 315846
rect 247040 298172 247092 298178
rect 247040 298114 247092 298120
rect 247316 298172 247368 298178
rect 247316 298114 247368 298120
rect 247052 289882 247080 298114
rect 247040 289876 247092 289882
rect 247040 289818 247092 289824
rect 247224 289876 247276 289882
rect 247224 289818 247276 289824
rect 247236 282962 247264 289818
rect 247236 282934 247356 282962
rect 247328 282826 247356 282934
rect 247144 282798 247356 282826
rect 247144 280106 247172 282798
rect 247052 280078 247172 280106
rect 245934 278760 245990 278769
rect 245934 278695 245990 278704
rect 246118 278760 246174 278769
rect 246118 278695 246174 278704
rect 246132 269142 246160 278695
rect 247052 270570 247080 280078
rect 247040 270564 247092 270570
rect 247040 270506 247092 270512
rect 247224 270564 247276 270570
rect 247224 270506 247276 270512
rect 245936 269136 245988 269142
rect 245936 269078 245988 269084
rect 246120 269136 246172 269142
rect 247236 269090 247264 270506
rect 246120 269078 246172 269084
rect 245948 265690 245976 269078
rect 247144 269062 247264 269090
rect 245948 265662 246068 265690
rect 246040 263514 246068 265662
rect 245856 263486 246068 263514
rect 245856 259457 245884 263486
rect 247144 260914 247172 269062
rect 247132 260908 247184 260914
rect 247132 260850 247184 260856
rect 247224 259616 247276 259622
rect 247224 259558 247276 259564
rect 245842 259448 245898 259457
rect 245842 259383 245898 259392
rect 246026 259448 246082 259457
rect 246026 259383 246082 259392
rect 246040 249830 246068 259383
rect 247236 258058 247264 259558
rect 247224 258052 247276 258058
rect 247224 257994 247276 258000
rect 245844 249824 245896 249830
rect 245842 249792 245844 249801
rect 246028 249824 246080 249830
rect 245896 249792 245898 249801
rect 246028 249766 246080 249772
rect 246118 249792 246174 249801
rect 245842 249727 245898 249736
rect 246118 249727 246174 249736
rect 247224 249756 247276 249762
rect 246132 240174 246160 249727
rect 247224 249698 247276 249704
rect 245936 240168 245988 240174
rect 245936 240110 245988 240116
rect 246120 240168 246172 240174
rect 246120 240110 246172 240116
rect 245948 227338 245976 240110
rect 247236 239986 247264 249698
rect 247236 239958 247356 239986
rect 245948 227310 246068 227338
rect 246040 220862 246068 227310
rect 245844 220856 245896 220862
rect 245844 220798 245896 220804
rect 246028 220856 246080 220862
rect 247328 220833 247356 239958
rect 246028 220798 246080 220804
rect 247314 220824 247370 220833
rect 245856 212566 245884 220798
rect 247314 220759 247370 220768
rect 245844 212560 245896 212566
rect 245844 212502 245896 212508
rect 245936 212560 245988 212566
rect 245936 212502 245988 212508
rect 245948 202910 245976 212502
rect 247222 211168 247278 211177
rect 246948 211132 247000 211138
rect 247222 211103 247224 211112
rect 246948 211074 247000 211080
rect 247276 211103 247278 211112
rect 247224 211074 247276 211080
rect 245844 202904 245896 202910
rect 245844 202846 245896 202852
rect 245936 202904 245988 202910
rect 245936 202846 245988 202852
rect 245856 191894 245884 202846
rect 246960 201521 246988 211074
rect 246946 201512 247002 201521
rect 246946 201447 247002 201456
rect 247130 201512 247186 201521
rect 247130 201447 247186 201456
rect 247144 193254 247172 201447
rect 247132 193248 247184 193254
rect 247132 193190 247184 193196
rect 247224 193248 247276 193254
rect 247224 193190 247276 193196
rect 245844 191888 245896 191894
rect 245844 191830 245896 191836
rect 247236 182186 247264 193190
rect 247144 182158 247264 182186
rect 245752 180940 245804 180946
rect 245752 180882 245804 180888
rect 245660 180872 245712 180878
rect 245660 180814 245712 180820
rect 245660 180736 245712 180742
rect 245660 180678 245712 180684
rect 245384 180668 245436 180674
rect 245384 180610 245436 180616
rect 244372 171080 244424 171086
rect 244372 171022 244424 171028
rect 244556 171012 244608 171018
rect 244556 170954 244608 170960
rect 244568 144945 244596 170954
rect 244370 144936 244426 144945
rect 244370 144871 244426 144880
rect 244554 144936 244610 144945
rect 244554 144871 244610 144880
rect 244384 138106 244412 144871
rect 244372 138100 244424 138106
rect 244372 138042 244424 138048
rect 244372 137964 244424 137970
rect 244372 137906 244424 137912
rect 244384 130370 244412 137906
rect 244384 130342 244504 130370
rect 244476 114578 244504 130342
rect 244280 114572 244332 114578
rect 244280 114514 244332 114520
rect 244464 114572 244516 114578
rect 244464 114514 244516 114520
rect 244292 113150 244320 114514
rect 244280 113144 244332 113150
rect 244280 113086 244332 113092
rect 244372 103556 244424 103562
rect 244372 103498 244424 103504
rect 244384 103426 244412 103498
rect 244372 103420 244424 103426
rect 244372 103362 244424 103368
rect 244556 103420 244608 103426
rect 244556 103362 244608 103368
rect 244568 96506 244596 103362
rect 244476 96478 244596 96506
rect 244476 71210 244504 96478
rect 244476 71182 244596 71210
rect 244568 66473 244596 71182
rect 244554 66464 244610 66473
rect 244554 66399 244610 66408
rect 244370 66328 244426 66337
rect 244370 66263 244426 66272
rect 244384 66230 244412 66263
rect 244372 66224 244424 66230
rect 244372 66166 244424 66172
rect 244464 56636 244516 56642
rect 244464 56578 244516 56584
rect 244476 53258 244504 56578
rect 244476 53230 244596 53258
rect 244568 48346 244596 53230
rect 244372 48340 244424 48346
rect 244372 48282 244424 48288
rect 244556 48340 244608 48346
rect 244556 48282 244608 48288
rect 244384 38758 244412 48282
rect 245566 48240 245622 48249
rect 245566 48175 245622 48184
rect 245580 40390 245608 48175
rect 245568 40384 245620 40390
rect 245568 40326 245620 40332
rect 244372 38752 244424 38758
rect 244372 38694 244424 38700
rect 244464 38684 244516 38690
rect 244464 38626 244516 38632
rect 244476 22166 244504 38626
rect 244464 22160 244516 22166
rect 244464 22102 244516 22108
rect 244188 16652 244240 16658
rect 244188 16594 244240 16600
rect 244200 11098 244228 16594
rect 244200 11070 244320 11098
rect 243176 9104 243228 9110
rect 243176 9046 243228 9052
rect 243084 3732 243136 3738
rect 243084 3674 243136 3680
rect 243188 480 243216 9046
rect 244292 8022 244320 11070
rect 244280 8016 244332 8022
rect 244280 7958 244332 7964
rect 245568 7812 245620 7818
rect 245568 7754 245620 7760
rect 244372 5092 244424 5098
rect 244372 5034 244424 5040
rect 244384 480 244412 5034
rect 245580 480 245608 7754
rect 245672 3806 245700 180678
rect 245844 180668 245896 180674
rect 245844 180610 245896 180616
rect 245752 179444 245804 179450
rect 245752 179386 245804 179392
rect 245764 160041 245792 179386
rect 245750 160032 245806 160041
rect 245750 159967 245806 159976
rect 245856 156602 245884 180610
rect 247144 176798 247172 182158
rect 247132 176792 247184 176798
rect 247132 176734 247184 176740
rect 247224 176724 247276 176730
rect 247224 176666 247276 176672
rect 247236 171086 247264 176666
rect 247224 171080 247276 171086
rect 247224 171022 247276 171028
rect 247132 161492 247184 161498
rect 247132 161434 247184 161440
rect 246118 160032 246174 160041
rect 246118 159967 246174 159976
rect 245844 156596 245896 156602
rect 245844 156538 245896 156544
rect 246028 156596 246080 156602
rect 246028 156538 246080 156544
rect 245752 150476 245804 150482
rect 245752 150418 245804 150424
rect 245764 140729 245792 150418
rect 246040 143585 246068 156538
rect 246132 150482 246160 159967
rect 247144 153270 247172 161434
rect 247132 153264 247184 153270
rect 247132 153206 247184 153212
rect 247040 153196 247092 153202
rect 247040 153138 247092 153144
rect 246120 150476 246172 150482
rect 246120 150418 246172 150424
rect 245842 143576 245898 143585
rect 245842 143511 245844 143520
rect 245896 143511 245898 143520
rect 246026 143576 246082 143585
rect 246026 143511 246082 143520
rect 245844 143482 245896 143488
rect 245750 140720 245806 140729
rect 245750 140655 245806 140664
rect 245934 140720 245990 140729
rect 245934 140655 245990 140664
rect 245844 137964 245896 137970
rect 245844 137906 245896 137912
rect 245752 131164 245804 131170
rect 245752 131106 245804 131112
rect 245764 102082 245792 131106
rect 245856 130370 245884 137906
rect 245948 131170 245976 140655
rect 247052 133929 247080 153138
rect 247038 133920 247094 133929
rect 247038 133855 247094 133864
rect 247314 133784 247370 133793
rect 247314 133719 247370 133728
rect 245936 131164 245988 131170
rect 245936 131106 245988 131112
rect 245856 130342 245976 130370
rect 245948 116006 245976 130342
rect 247328 124166 247356 133719
rect 247316 124160 247368 124166
rect 247316 124102 247368 124108
rect 245936 116000 245988 116006
rect 245936 115942 245988 115948
rect 245936 114572 245988 114578
rect 245936 114514 245988 114520
rect 247132 114572 247184 114578
rect 247132 114514 247184 114520
rect 245948 106282 245976 114514
rect 247144 106350 247172 114514
rect 247132 106344 247184 106350
rect 247132 106286 247184 106292
rect 245936 106276 245988 106282
rect 245936 106218 245988 106224
rect 247132 106208 247184 106214
rect 247132 106150 247184 106156
rect 247144 103494 247172 106150
rect 247132 103488 247184 103494
rect 247132 103430 247184 103436
rect 245764 102054 245884 102082
rect 245856 92546 245884 102054
rect 245936 96688 245988 96694
rect 245936 96630 245988 96636
rect 245752 92540 245804 92546
rect 245752 92482 245804 92488
rect 245844 92540 245896 92546
rect 245844 92482 245896 92488
rect 245764 82770 245792 92482
rect 245764 82742 245884 82770
rect 245856 73234 245884 82742
rect 245752 73228 245804 73234
rect 245752 73170 245804 73176
rect 245844 73228 245896 73234
rect 245844 73170 245896 73176
rect 245764 44130 245792 73170
rect 245948 67726 245976 96630
rect 247224 93900 247276 93906
rect 247224 93842 247276 93848
rect 247236 80102 247264 93842
rect 247224 80096 247276 80102
rect 247224 80038 247276 80044
rect 247132 73228 247184 73234
rect 247132 73170 247184 73176
rect 247144 69578 247172 73170
rect 247144 69550 247264 69578
rect 245936 67720 245988 67726
rect 245936 67662 245988 67668
rect 245936 67516 245988 67522
rect 245936 67458 245988 67464
rect 245948 66230 245976 67458
rect 245936 66224 245988 66230
rect 245936 66166 245988 66172
rect 246028 66156 246080 66162
rect 246028 66098 246080 66104
rect 246040 60602 246068 66098
rect 245948 60574 246068 60602
rect 245948 48385 245976 60574
rect 247236 55214 247264 69550
rect 247224 55208 247276 55214
rect 247224 55150 247276 55156
rect 245934 48376 245990 48385
rect 245934 48311 245990 48320
rect 247224 45620 247276 45626
rect 247224 45562 247276 45568
rect 245752 44124 245804 44130
rect 245752 44066 245804 44072
rect 245936 40384 245988 40390
rect 245936 40326 245988 40332
rect 245752 34536 245804 34542
rect 245752 34478 245804 34484
rect 245764 5545 245792 34478
rect 245948 26246 245976 40326
rect 247236 35902 247264 45562
rect 247224 35896 247276 35902
rect 247224 35838 247276 35844
rect 247224 26376 247276 26382
rect 247224 26318 247276 26324
rect 247236 26246 247264 26318
rect 245936 26240 245988 26246
rect 245936 26182 245988 26188
rect 247224 26240 247276 26246
rect 247224 26182 247276 26188
rect 245844 16652 245896 16658
rect 245844 16594 245896 16600
rect 245856 13138 245884 16594
rect 245856 13110 245976 13138
rect 245948 8090 245976 13110
rect 246764 8356 246816 8362
rect 246764 8298 246816 8304
rect 245936 8084 245988 8090
rect 245936 8026 245988 8032
rect 245750 5536 245806 5545
rect 245750 5471 245806 5480
rect 245660 3800 245712 3806
rect 245660 3742 245712 3748
rect 246776 480 246804 8298
rect 247696 3942 247724 337350
rect 248512 335504 248564 335510
rect 248512 335446 248564 335452
rect 248418 110800 248474 110809
rect 248418 110735 248420 110744
rect 248472 110735 248474 110744
rect 248420 110706 248472 110712
rect 248524 5234 248552 335446
rect 248512 5228 248564 5234
rect 248512 5170 248564 5176
rect 247960 5160 248012 5166
rect 247960 5102 248012 5108
rect 247684 3936 247736 3942
rect 247684 3878 247736 3884
rect 247972 480 248000 5102
rect 248708 4010 248736 340054
rect 249064 337408 249116 337414
rect 249064 337350 249116 337356
rect 249076 4078 249104 337350
rect 249168 335510 249196 340054
rect 249156 335504 249208 335510
rect 249156 335446 249208 335452
rect 249904 9246 249932 340054
rect 250548 337414 250576 340068
rect 250640 340054 251022 340082
rect 251284 340054 251574 340082
rect 250536 337408 250588 337414
rect 250536 337350 250588 337356
rect 250640 335578 250668 340054
rect 250720 337408 250772 337414
rect 250720 337350 250772 337356
rect 250628 335572 250680 335578
rect 250628 335514 250680 335520
rect 250732 335458 250760 337350
rect 250456 335430 250760 335458
rect 250168 327140 250220 327146
rect 250168 327082 250220 327088
rect 250180 317422 250208 327082
rect 250168 317416 250220 317422
rect 250168 317358 250220 317364
rect 250168 312588 250220 312594
rect 250168 312530 250220 312536
rect 250180 280158 250208 312530
rect 250076 280152 250128 280158
rect 250076 280094 250128 280100
rect 250168 280152 250220 280158
rect 250168 280094 250220 280100
rect 250088 273970 250116 280094
rect 250076 273964 250128 273970
rect 250076 273906 250128 273912
rect 250260 273964 250312 273970
rect 250260 273906 250312 273912
rect 250272 269090 250300 273906
rect 250180 269062 250300 269090
rect 250180 264314 250208 269062
rect 250168 264308 250220 264314
rect 250168 264250 250220 264256
rect 250168 259480 250220 259486
rect 250168 259422 250220 259428
rect 250180 251190 250208 259422
rect 250168 251184 250220 251190
rect 250168 251126 250220 251132
rect 250168 241528 250220 241534
rect 250168 241470 250220 241476
rect 250180 240122 250208 241470
rect 250088 240094 250208 240122
rect 250088 234666 250116 240094
rect 250076 234660 250128 234666
rect 250076 234602 250128 234608
rect 250168 230512 250220 230518
rect 250168 230454 250220 230460
rect 250180 217410 250208 230454
rect 250180 217382 250300 217410
rect 250272 212566 250300 217382
rect 250076 212560 250128 212566
rect 250076 212502 250128 212508
rect 250260 212560 250312 212566
rect 250260 212502 250312 212508
rect 250088 211138 250116 212502
rect 249984 211132 250036 211138
rect 249984 211074 250036 211080
rect 250076 211132 250128 211138
rect 250076 211074 250128 211080
rect 249996 201521 250024 211074
rect 249982 201512 250038 201521
rect 250166 201512 250222 201521
rect 249982 201447 250038 201456
rect 250076 201476 250128 201482
rect 250166 201447 250168 201456
rect 250076 201418 250128 201424
rect 250220 201447 250222 201456
rect 250168 201418 250220 201424
rect 250088 200122 250116 201418
rect 250076 200116 250128 200122
rect 250076 200058 250128 200064
rect 250260 200116 250312 200122
rect 250260 200058 250312 200064
rect 250272 176798 250300 200058
rect 250260 176792 250312 176798
rect 250260 176734 250312 176740
rect 250076 176724 250128 176730
rect 250076 176666 250128 176672
rect 250088 164234 250116 176666
rect 250088 164206 250208 164234
rect 250180 162858 250208 164206
rect 250168 162852 250220 162858
rect 250168 162794 250220 162800
rect 250260 162852 250312 162858
rect 250260 162794 250312 162800
rect 250272 149546 250300 162794
rect 250180 149518 250300 149546
rect 250180 143546 250208 149518
rect 250168 143540 250220 143546
rect 250168 143482 250220 143488
rect 250168 137964 250220 137970
rect 250168 137906 250220 137912
rect 250180 116113 250208 137906
rect 250166 116104 250222 116113
rect 250166 116039 250222 116048
rect 250074 115968 250130 115977
rect 250074 115903 250130 115912
rect 250088 111058 250116 115903
rect 250088 111030 250208 111058
rect 250180 101402 250208 111030
rect 250088 101374 250208 101402
rect 250088 72434 250116 101374
rect 250088 72406 250208 72434
rect 250180 56642 250208 72406
rect 250168 56636 250220 56642
rect 250168 56578 250220 56584
rect 250168 53848 250220 53854
rect 250168 53790 250220 53796
rect 250180 47054 250208 53790
rect 250168 47048 250220 47054
rect 250168 46990 250220 46996
rect 250076 46912 250128 46918
rect 250076 46854 250128 46860
rect 250088 45506 250116 46854
rect 249996 45478 250116 45506
rect 249996 35970 250024 45478
rect 249984 35964 250036 35970
rect 249984 35906 250036 35912
rect 250076 35964 250128 35970
rect 250076 35906 250128 35912
rect 250088 35834 250116 35906
rect 250076 35828 250128 35834
rect 250076 35770 250128 35776
rect 250168 26308 250220 26314
rect 250168 26250 250220 26256
rect 250180 22166 250208 26250
rect 250168 22160 250220 22166
rect 250168 22102 250220 22108
rect 249984 16652 250036 16658
rect 249984 16594 250036 16600
rect 249892 9240 249944 9246
rect 249892 9182 249944 9188
rect 249156 7880 249208 7886
rect 249156 7822 249208 7828
rect 249064 4072 249116 4078
rect 249064 4014 249116 4020
rect 248696 4004 248748 4010
rect 248696 3946 248748 3952
rect 249168 480 249196 7822
rect 249996 6225 250024 16594
rect 250352 9172 250404 9178
rect 250352 9114 250404 9120
rect 249982 6216 250038 6225
rect 249982 6151 250038 6160
rect 250364 480 250392 9114
rect 250456 4146 250484 335430
rect 251178 280120 251234 280129
rect 251178 280055 251234 280064
rect 251192 270570 251220 280055
rect 251180 270564 251232 270570
rect 251180 270506 251232 270512
rect 251178 260808 251234 260817
rect 251178 260743 251234 260752
rect 251192 251258 251220 260743
rect 251180 251252 251232 251258
rect 251180 251194 251232 251200
rect 251178 249792 251234 249801
rect 251178 249727 251234 249736
rect 251192 240174 251220 249727
rect 251180 240168 251232 240174
rect 251086 240136 251142 240145
rect 251180 240110 251232 240116
rect 251086 240071 251142 240080
rect 251100 230518 251128 240071
rect 251088 230512 251140 230518
rect 251088 230454 251140 230460
rect 251180 172576 251232 172582
rect 251180 172518 251232 172524
rect 251192 164286 251220 172518
rect 251284 164354 251312 340054
rect 252020 338026 252048 340068
rect 252112 340054 252494 340082
rect 252664 340054 253046 340082
rect 252008 338020 252060 338026
rect 252008 337962 252060 337968
rect 252112 335730 252140 340054
rect 252192 337612 252244 337618
rect 252192 337554 252244 337560
rect 251468 335702 252140 335730
rect 251468 323626 251496 335702
rect 252204 334370 252232 337554
rect 251836 334342 252232 334370
rect 251468 323598 251588 323626
rect 251560 317422 251588 323598
rect 251548 317416 251600 317422
rect 251548 317358 251600 317364
rect 251548 307828 251600 307834
rect 251548 307770 251600 307776
rect 251560 307737 251588 307770
rect 251546 307728 251602 307737
rect 251546 307663 251602 307672
rect 251546 298208 251602 298217
rect 251546 298143 251602 298152
rect 251560 298110 251588 298143
rect 251548 298104 251600 298110
rect 251548 298046 251600 298052
rect 251364 288448 251416 288454
rect 251364 288390 251416 288396
rect 251376 280129 251404 288390
rect 251362 280120 251418 280129
rect 251362 280055 251418 280064
rect 251456 270564 251508 270570
rect 251456 270506 251508 270512
rect 251468 265690 251496 270506
rect 251468 265662 251588 265690
rect 251560 263514 251588 265662
rect 251376 263486 251588 263514
rect 251376 260817 251404 263486
rect 251362 260808 251418 260817
rect 251362 260743 251418 260752
rect 251456 251252 251508 251258
rect 251456 251194 251508 251200
rect 251468 249801 251496 251194
rect 251454 249792 251510 249801
rect 251454 249727 251510 249736
rect 251364 240168 251416 240174
rect 251362 240136 251364 240145
rect 251416 240136 251418 240145
rect 251362 240071 251418 240080
rect 251364 230512 251416 230518
rect 251362 230480 251364 230489
rect 251416 230480 251418 230489
rect 251362 230415 251418 230424
rect 251546 230480 251602 230489
rect 251546 230415 251602 230424
rect 251560 220862 251588 230415
rect 251548 220856 251600 220862
rect 251548 220798 251600 220804
rect 251640 220856 251692 220862
rect 251640 220798 251692 220804
rect 251652 212514 251680 220798
rect 251560 212486 251680 212514
rect 251560 205578 251588 212486
rect 251468 205550 251588 205578
rect 251468 202722 251496 205550
rect 251468 202694 251588 202722
rect 251560 193225 251588 202694
rect 251362 193216 251418 193225
rect 251362 193151 251418 193160
rect 251546 193216 251602 193225
rect 251546 193151 251602 193160
rect 251376 186386 251404 193151
rect 251364 186380 251416 186386
rect 251364 186322 251416 186328
rect 251364 186244 251416 186250
rect 251364 186186 251416 186192
rect 251376 183530 251404 186186
rect 251364 183524 251416 183530
rect 251364 183466 251416 183472
rect 251548 183524 251600 183530
rect 251548 183466 251600 183472
rect 251560 172582 251588 183466
rect 251548 172576 251600 172582
rect 251548 172518 251600 172524
rect 251272 164348 251324 164354
rect 251272 164290 251324 164296
rect 251180 164280 251232 164286
rect 251180 164222 251232 164228
rect 251272 164212 251324 164218
rect 251272 164154 251324 164160
rect 251178 76120 251234 76129
rect 251178 76055 251234 76064
rect 251192 75721 251220 76055
rect 251178 75712 251234 75721
rect 251178 75647 251234 75656
rect 251284 10334 251312 164154
rect 251364 164144 251416 164150
rect 251364 164086 251416 164092
rect 251376 162858 251404 164086
rect 251364 162852 251416 162858
rect 251364 162794 251416 162800
rect 251640 162852 251692 162858
rect 251640 162794 251692 162800
rect 251652 154442 251680 162794
rect 251560 154414 251680 154442
rect 251560 143682 251588 154414
rect 251364 143676 251416 143682
rect 251364 143618 251416 143624
rect 251548 143676 251600 143682
rect 251548 143618 251600 143624
rect 251376 142118 251404 143618
rect 251364 142112 251416 142118
rect 251364 142054 251416 142060
rect 251456 132524 251508 132530
rect 251456 132466 251508 132472
rect 251468 124250 251496 132466
rect 251376 124222 251496 124250
rect 251376 122806 251404 124222
rect 251364 122800 251416 122806
rect 251364 122742 251416 122748
rect 251456 113212 251508 113218
rect 251456 113154 251508 113160
rect 251468 77602 251496 113154
rect 251468 77574 251680 77602
rect 251652 77353 251680 77574
rect 251454 77344 251510 77353
rect 251454 77279 251510 77288
rect 251638 77344 251694 77353
rect 251638 77279 251694 77288
rect 251468 77246 251496 77279
rect 251456 77240 251508 77246
rect 251456 77182 251508 77188
rect 251364 64932 251416 64938
rect 251364 64874 251416 64880
rect 251376 45558 251404 64874
rect 251364 45552 251416 45558
rect 251364 45494 251416 45500
rect 251456 35964 251508 35970
rect 251456 35906 251508 35912
rect 251468 28914 251496 35906
rect 251468 28886 251588 28914
rect 251560 19378 251588 28886
rect 251364 19372 251416 19378
rect 251364 19314 251416 19320
rect 251548 19372 251600 19378
rect 251548 19314 251600 19320
rect 251376 19281 251404 19314
rect 251362 19272 251418 19281
rect 251362 19207 251418 19216
rect 251638 19136 251694 19145
rect 251638 19071 251694 19080
rect 251272 10328 251324 10334
rect 251272 10270 251324 10276
rect 251652 9761 251680 19071
rect 251454 9752 251510 9761
rect 251454 9687 251510 9696
rect 251638 9752 251694 9761
rect 251638 9687 251694 9696
rect 251468 6186 251496 9687
rect 251456 6180 251508 6186
rect 251456 6122 251508 6128
rect 251456 5228 251508 5234
rect 251456 5170 251508 5176
rect 250444 4140 250496 4146
rect 250444 4082 250496 4088
rect 251468 480 251496 5170
rect 251836 3398 251864 334342
rect 252664 10402 252692 340054
rect 253204 337544 253256 337550
rect 253204 337486 253256 337492
rect 253110 29336 253166 29345
rect 253110 29271 253166 29280
rect 253124 29238 253152 29271
rect 253112 29232 253164 29238
rect 253112 29174 253164 29180
rect 252652 10396 252704 10402
rect 252652 10338 252704 10344
rect 252652 7948 252704 7954
rect 252652 7890 252704 7896
rect 251824 3392 251876 3398
rect 251824 3334 251876 3340
rect 252664 480 252692 7890
rect 253216 3330 253244 337486
rect 253492 337414 253520 340068
rect 253480 337408 253532 337414
rect 253480 337350 253532 337356
rect 253848 9240 253900 9246
rect 253848 9182 253900 9188
rect 253204 3324 253256 3330
rect 253204 3266 253256 3272
rect 253860 480 253888 9182
rect 253952 6254 253980 340068
rect 254044 340054 254518 340082
rect 254044 10470 254072 340054
rect 254584 337748 254636 337754
rect 254584 337690 254636 337696
rect 254124 110764 254176 110770
rect 254124 110706 254176 110712
rect 254136 110673 254164 110706
rect 254122 110664 254178 110673
rect 254122 110599 254178 110608
rect 254032 10464 254084 10470
rect 254032 10406 254084 10412
rect 253940 6248 253992 6254
rect 253940 6190 253992 6196
rect 254596 3262 254624 337690
rect 254964 337278 254992 340068
rect 255438 340054 255544 340082
rect 254952 337272 255004 337278
rect 254952 337214 255004 337220
rect 255516 6322 255544 340054
rect 255608 340054 255990 340082
rect 255608 10538 255636 340054
rect 256436 337618 256464 340068
rect 256804 340054 256910 340082
rect 256988 340054 257462 340082
rect 256424 337612 256476 337618
rect 256424 337554 256476 337560
rect 255964 337272 256016 337278
rect 255964 337214 256016 337220
rect 255596 10532 255648 10538
rect 255596 10474 255648 10480
rect 255504 6316 255556 6322
rect 255504 6258 255556 6264
rect 255044 3460 255096 3466
rect 255044 3402 255096 3408
rect 254584 3256 254636 3262
rect 254584 3198 254636 3204
rect 255056 480 255084 3402
rect 255976 3194 256004 337214
rect 256240 8016 256292 8022
rect 256240 7958 256292 7964
rect 255964 3188 256016 3194
rect 255964 3130 256016 3136
rect 256252 480 256280 7958
rect 256804 6390 256832 340054
rect 256792 6384 256844 6390
rect 256792 6326 256844 6332
rect 256988 5302 257016 340054
rect 257908 338094 257936 340068
rect 258276 340054 258382 340082
rect 258552 340054 258934 340082
rect 257896 338088 257948 338094
rect 257896 338030 257948 338036
rect 257344 337408 257396 337414
rect 257344 337350 257396 337356
rect 256976 5296 257028 5302
rect 256976 5238 257028 5244
rect 257356 3126 257384 337350
rect 258172 334620 258224 334626
rect 258172 334562 258224 334568
rect 257988 29232 258040 29238
rect 257986 29200 257988 29209
rect 258040 29200 258042 29209
rect 257986 29135 258042 29144
rect 258184 13190 258212 334562
rect 258172 13184 258224 13190
rect 258172 13126 258224 13132
rect 258276 6458 258304 340054
rect 258552 334626 258580 340054
rect 258816 337884 258868 337890
rect 258816 337826 258868 337832
rect 258724 337476 258776 337482
rect 258724 337418 258776 337424
rect 258540 334620 258592 334626
rect 258540 334562 258592 334568
rect 258264 6452 258316 6458
rect 258264 6394 258316 6400
rect 257436 4004 257488 4010
rect 257436 3946 257488 3952
rect 257344 3120 257396 3126
rect 257344 3062 257396 3068
rect 257448 480 257476 3946
rect 258632 3528 258684 3534
rect 258632 3470 258684 3476
rect 258644 480 258672 3470
rect 258736 2990 258764 337418
rect 258828 3058 258856 337826
rect 259380 337550 259408 340068
rect 259472 340054 259854 340082
rect 260116 340054 260406 340082
rect 259368 337544 259420 337550
rect 259368 337486 259420 337492
rect 259366 110664 259422 110673
rect 259366 110599 259368 110608
rect 259420 110599 259422 110608
rect 259368 110570 259420 110576
rect 259472 6526 259500 340054
rect 260116 337822 260144 340054
rect 259644 337816 259696 337822
rect 259644 337758 259696 337764
rect 260104 337816 260156 337822
rect 260104 337758 260156 337764
rect 259656 331226 259684 337758
rect 260104 337680 260156 337686
rect 260104 337622 260156 337628
rect 259644 331220 259696 331226
rect 259644 331162 259696 331168
rect 259828 331220 259880 331226
rect 259828 331162 259880 331168
rect 259840 328438 259868 331162
rect 259828 328432 259880 328438
rect 259828 328374 259880 328380
rect 259920 318844 259972 318850
rect 259920 318786 259972 318792
rect 259932 311914 259960 318786
rect 259736 311908 259788 311914
rect 259736 311850 259788 311856
rect 259920 311908 259972 311914
rect 259920 311850 259972 311856
rect 259748 302326 259776 311850
rect 259736 302320 259788 302326
rect 259736 302262 259788 302268
rect 259644 296744 259696 296750
rect 259644 296686 259696 296692
rect 259656 269142 259684 296686
rect 259644 269136 259696 269142
rect 259644 269078 259696 269084
rect 259736 269136 259788 269142
rect 259736 269078 259788 269084
rect 259748 265690 259776 269078
rect 259564 265662 259776 265690
rect 259564 263514 259592 265662
rect 259564 263486 259684 263514
rect 259656 260794 259684 263486
rect 259656 260766 259776 260794
rect 259748 254658 259776 260766
rect 259736 254652 259788 254658
rect 259736 254594 259788 254600
rect 259644 241596 259696 241602
rect 259644 241538 259696 241544
rect 259656 230518 259684 241538
rect 259552 230512 259604 230518
rect 259552 230454 259604 230460
rect 259644 230512 259696 230518
rect 259644 230454 259696 230460
rect 259564 227066 259592 230454
rect 259564 227038 259684 227066
rect 259656 222193 259684 227038
rect 259642 222184 259698 222193
rect 259642 222119 259698 222128
rect 259734 221912 259790 221921
rect 259734 221847 259790 221856
rect 259748 205578 259776 221847
rect 259656 205550 259776 205578
rect 259656 202881 259684 205550
rect 259642 202872 259698 202881
rect 259642 202807 259698 202816
rect 259918 202872 259974 202881
rect 259918 202807 259974 202816
rect 259932 193254 259960 202807
rect 259736 193248 259788 193254
rect 259736 193190 259788 193196
rect 259920 193248 259972 193254
rect 259920 193190 259972 193196
rect 259748 186266 259776 193190
rect 259656 186238 259776 186266
rect 259656 183569 259684 186238
rect 259642 183560 259698 183569
rect 259642 183495 259698 183504
rect 259918 183560 259974 183569
rect 259918 183495 259974 183504
rect 259932 173942 259960 183495
rect 259736 173936 259788 173942
rect 259736 173878 259788 173884
rect 259920 173936 259972 173942
rect 259920 173878 259972 173884
rect 259748 157434 259776 173878
rect 259656 157406 259776 157434
rect 259656 157298 259684 157406
rect 259656 157270 259776 157298
rect 259748 154562 259776 157270
rect 259736 154556 259788 154562
rect 259736 154498 259788 154504
rect 259736 147620 259788 147626
rect 259736 147562 259788 147568
rect 259748 144922 259776 147562
rect 259748 144894 259868 144922
rect 259656 138038 259684 138069
rect 259840 138038 259868 144894
rect 259644 138032 259696 138038
rect 259828 138032 259880 138038
rect 259696 137980 259776 137986
rect 259644 137974 259776 137980
rect 259828 137974 259880 137980
rect 259656 137958 259776 137974
rect 259748 132462 259776 137958
rect 259736 132456 259788 132462
rect 259736 132398 259788 132404
rect 259644 122868 259696 122874
rect 259644 122810 259696 122816
rect 259656 122754 259684 122810
rect 259734 122768 259790 122777
rect 259656 122726 259734 122754
rect 259734 122703 259790 122712
rect 259918 122768 259974 122777
rect 259918 122703 259974 122712
rect 259932 113218 259960 122703
rect 259736 113212 259788 113218
rect 259736 113154 259788 113160
rect 259920 113212 259972 113218
rect 259920 113154 259972 113160
rect 259748 104802 259776 113154
rect 259656 104774 259776 104802
rect 259656 95198 259684 104774
rect 259644 95192 259696 95198
rect 259644 95134 259696 95140
rect 259736 77308 259788 77314
rect 259736 77250 259788 77256
rect 259748 62694 259776 77250
rect 259736 62688 259788 62694
rect 259736 62630 259788 62636
rect 259920 62620 259972 62626
rect 259920 62562 259972 62568
rect 259932 56574 259960 62562
rect 259920 56568 259972 56574
rect 259920 56510 259972 56516
rect 259736 45620 259788 45626
rect 259736 45562 259788 45568
rect 259748 37194 259776 45562
rect 259644 37188 259696 37194
rect 259644 37130 259696 37136
rect 259736 37188 259788 37194
rect 259736 37130 259788 37136
rect 259656 35902 259684 37130
rect 259644 35896 259696 35902
rect 259644 35838 259696 35844
rect 259552 26376 259604 26382
rect 259552 26318 259604 26324
rect 259564 26246 259592 26318
rect 259552 26240 259604 26246
rect 259552 26182 259604 26188
rect 259552 17944 259604 17950
rect 259552 17886 259604 17892
rect 259564 14482 259592 17886
rect 259552 14476 259604 14482
rect 259552 14418 259604 14424
rect 259828 8084 259880 8090
rect 259828 8026 259880 8032
rect 259460 6520 259512 6526
rect 259460 6462 259512 6468
rect 258816 3052 258868 3058
rect 258816 2994 258868 3000
rect 258724 2984 258776 2990
rect 258724 2926 258776 2932
rect 259840 480 259868 8026
rect 260116 2922 260144 337622
rect 260852 337346 260880 340068
rect 261036 340054 261326 340082
rect 261496 340054 261878 340082
rect 260840 337340 260892 337346
rect 260840 337282 260892 337288
rect 260932 335640 260984 335646
rect 260932 335582 260984 335588
rect 260944 14550 260972 335582
rect 260932 14544 260984 14550
rect 260932 14486 260984 14492
rect 261036 6594 261064 340054
rect 261392 337612 261444 337618
rect 261392 337554 261444 337560
rect 261404 334370 261432 337554
rect 261496 335646 261524 340054
rect 262324 337754 262352 340068
rect 262416 340054 262798 340082
rect 263060 340054 263350 340082
rect 262312 337748 262364 337754
rect 262312 337690 262364 337696
rect 261484 335640 261536 335646
rect 261484 335582 261536 335588
rect 261404 334342 261524 334370
rect 261024 6588 261076 6594
rect 261024 6530 261076 6536
rect 260104 2916 260156 2922
rect 260104 2858 260156 2864
rect 261496 2854 261524 334342
rect 262312 258052 262364 258058
rect 262312 257994 262364 258000
rect 262324 248441 262352 257994
rect 262310 248432 262366 248441
rect 262310 248367 262366 248376
rect 262416 8158 262444 340054
rect 263060 335646 263088 340054
rect 263796 337074 263824 340068
rect 263888 340054 264270 340082
rect 264440 340054 264822 340082
rect 263784 337068 263836 337074
rect 263784 337010 263836 337016
rect 262588 335640 262640 335646
rect 262588 335582 262640 335588
rect 263048 335640 263100 335646
rect 263048 335582 263100 335588
rect 263692 335640 263744 335646
rect 263692 335582 263744 335588
rect 262600 331226 262628 335582
rect 262588 331220 262640 331226
rect 262588 331162 262640 331168
rect 262772 331220 262824 331226
rect 262772 331162 262824 331168
rect 262784 321638 262812 331162
rect 262772 321632 262824 321638
rect 262772 321574 262824 321580
rect 262864 321496 262916 321502
rect 262864 321438 262916 321444
rect 262876 309210 262904 321438
rect 262692 309182 262904 309210
rect 262692 299674 262720 309182
rect 262680 299668 262732 299674
rect 262680 299610 262732 299616
rect 262588 296744 262640 296750
rect 262588 296686 262640 296692
rect 262600 269113 262628 296686
rect 262586 269104 262642 269113
rect 262586 269039 262642 269048
rect 262678 268968 262734 268977
rect 262678 268903 262734 268912
rect 262692 263514 262720 268903
rect 262600 263486 262720 263514
rect 262600 258058 262628 263486
rect 262588 258052 262640 258058
rect 262588 257994 262640 258000
rect 262494 248432 262550 248441
rect 262494 248367 262550 248376
rect 262508 240174 262536 248367
rect 262600 240174 262628 240205
rect 262496 240168 262548 240174
rect 262496 240110 262548 240116
rect 262588 240168 262640 240174
rect 262640 240116 262720 240122
rect 262588 240110 262720 240116
rect 262600 240094 262720 240110
rect 262692 212158 262720 240094
rect 262496 212152 262548 212158
rect 262496 212094 262548 212100
rect 262680 212152 262732 212158
rect 262680 212094 262732 212100
rect 262508 202910 262536 212094
rect 262496 202904 262548 202910
rect 262588 202904 262640 202910
rect 262496 202846 262548 202852
rect 262586 202872 262588 202881
rect 262640 202872 262642 202881
rect 262586 202807 262642 202816
rect 262678 202736 262734 202745
rect 262678 202671 262734 202680
rect 262692 186266 262720 202671
rect 262600 186238 262720 186266
rect 262600 183569 262628 186238
rect 262586 183560 262642 183569
rect 262586 183495 262642 183504
rect 262678 183424 262734 183433
rect 262678 183359 262734 183368
rect 262692 157434 262720 183359
rect 262600 157406 262720 157434
rect 262600 157298 262628 157406
rect 262600 157270 262720 157298
rect 262692 149682 262720 157270
rect 262692 149654 262904 149682
rect 262876 147642 262904 149654
rect 262784 147614 262904 147642
rect 262784 144888 262812 147614
rect 262784 144860 262904 144888
rect 262876 135289 262904 144860
rect 262678 135280 262734 135289
rect 262678 135215 262734 135224
rect 262862 135280 262918 135289
rect 262862 135215 262918 135224
rect 262692 132462 262720 135215
rect 262680 132456 262732 132462
rect 262680 132398 262732 132404
rect 262588 122868 262640 122874
rect 262588 122810 262640 122816
rect 262600 109750 262628 122810
rect 262588 109744 262640 109750
rect 262588 109686 262640 109692
rect 262496 104916 262548 104922
rect 262496 104858 262548 104864
rect 262508 95266 262536 104858
rect 262496 95260 262548 95266
rect 262496 95202 262548 95208
rect 262588 95260 262640 95266
rect 262588 95202 262640 95208
rect 262600 93838 262628 95202
rect 262588 93832 262640 93838
rect 262588 93774 262640 93780
rect 262680 84244 262732 84250
rect 262680 84186 262732 84192
rect 262692 66201 262720 84186
rect 262678 66192 262734 66201
rect 262678 66127 262734 66136
rect 262954 66192 263010 66201
rect 262954 66127 263010 66136
rect 262968 61470 262996 66127
rect 262772 61464 262824 61470
rect 262772 61406 262824 61412
rect 262956 61464 263008 61470
rect 262956 61406 263008 61412
rect 262784 29034 262812 61406
rect 262680 29028 262732 29034
rect 262680 28970 262732 28976
rect 262772 29028 262824 29034
rect 262772 28970 262824 28976
rect 262692 22114 262720 28970
rect 262600 22086 262720 22114
rect 262600 14618 262628 22086
rect 263704 14686 263732 335582
rect 263692 14680 263744 14686
rect 263692 14622 263744 14628
rect 262588 14612 262640 14618
rect 262588 14554 262640 14560
rect 263888 8226 263916 340054
rect 264440 335646 264468 340054
rect 265268 336938 265296 340068
rect 265452 340054 265742 340082
rect 265912 340054 266294 340082
rect 265256 336932 265308 336938
rect 265256 336874 265308 336880
rect 264428 335640 264480 335646
rect 264428 335582 264480 335588
rect 265072 335640 265124 335646
rect 265452 335594 265480 340054
rect 265912 335646 265940 340054
rect 266740 337414 266768 340068
rect 266924 340054 267214 340082
rect 267384 340054 267674 340082
rect 266728 337408 266780 337414
rect 266728 337350 266780 337356
rect 265072 335582 265124 335588
rect 264978 193216 265034 193225
rect 264978 193151 265034 193160
rect 264992 183598 265020 193151
rect 264980 183592 265032 183598
rect 264980 183534 265032 183540
rect 264980 17944 265032 17950
rect 264980 17886 265032 17892
rect 264992 8401 265020 17886
rect 265084 14754 265112 335582
rect 265268 335566 265480 335594
rect 265900 335640 265952 335646
rect 265900 335582 265952 335588
rect 266452 335640 266504 335646
rect 266924 335594 266952 340054
rect 267384 335646 267412 340054
rect 268212 337210 268240 340068
rect 268396 340054 268686 340082
rect 269146 340054 269252 340082
rect 268200 337204 268252 337210
rect 268200 337146 268252 337152
rect 266452 335582 266504 335588
rect 265268 328438 265296 335566
rect 265256 328432 265308 328438
rect 265256 328374 265308 328380
rect 265348 328432 265400 328438
rect 265348 328374 265400 328380
rect 265360 327078 265388 328374
rect 265348 327072 265400 327078
rect 265348 327014 265400 327020
rect 265256 317484 265308 317490
rect 265256 317426 265308 317432
rect 265268 309126 265296 317426
rect 265256 309120 265308 309126
rect 265256 309062 265308 309068
rect 265348 300144 265400 300150
rect 265348 300086 265400 300092
rect 265360 293962 265388 300086
rect 265348 293956 265400 293962
rect 265348 293898 265400 293904
rect 265532 293956 265584 293962
rect 265532 293898 265584 293904
rect 265544 276049 265572 293898
rect 265254 276040 265310 276049
rect 265254 275975 265310 275984
rect 265530 276040 265586 276049
rect 265530 275975 265586 275984
rect 265268 269142 265296 275975
rect 265256 269136 265308 269142
rect 265256 269078 265308 269084
rect 265164 269068 265216 269074
rect 265164 269010 265216 269016
rect 265176 266393 265204 269010
rect 265162 266384 265218 266393
rect 265162 266319 265218 266328
rect 265346 266384 265402 266393
rect 265346 266319 265402 266328
rect 265360 259434 265388 266319
rect 265268 259406 265388 259434
rect 265268 248418 265296 259406
rect 265176 248390 265296 248418
rect 265176 234410 265204 248390
rect 265176 234382 265296 234410
rect 265268 227202 265296 234382
rect 265268 227174 265388 227202
rect 265360 222222 265388 227174
rect 265164 222216 265216 222222
rect 265162 222184 265164 222193
rect 265348 222216 265400 222222
rect 265216 222184 265218 222193
rect 265162 222119 265218 222128
rect 265346 222184 265348 222193
rect 265400 222184 265402 222193
rect 265346 222119 265402 222128
rect 265360 212548 265388 222119
rect 265268 212520 265388 212548
rect 265268 212514 265296 212520
rect 265176 212486 265296 212514
rect 265176 202881 265204 212486
rect 265162 202872 265218 202881
rect 265162 202807 265218 202816
rect 265346 202872 265402 202881
rect 265346 202807 265402 202816
rect 265360 193254 265388 202807
rect 265256 193248 265308 193254
rect 265254 193216 265256 193225
rect 265348 193248 265400 193254
rect 265308 193216 265310 193225
rect 265348 193190 265400 193196
rect 265254 193151 265310 193160
rect 265164 183592 265216 183598
rect 265162 183560 265164 183569
rect 265216 183560 265218 183569
rect 265162 183495 265218 183504
rect 265346 183560 265402 183569
rect 265346 183495 265402 183504
rect 265360 173942 265388 183495
rect 265256 173936 265308 173942
rect 265256 173878 265308 173884
rect 265348 173936 265400 173942
rect 265348 173878 265400 173884
rect 265268 161498 265296 173878
rect 265164 161492 265216 161498
rect 265164 161434 265216 161440
rect 265256 161492 265308 161498
rect 265256 161434 265308 161440
rect 265176 160070 265204 161434
rect 265164 160064 265216 160070
rect 265164 160006 265216 160012
rect 265348 150476 265400 150482
rect 265348 150418 265400 150424
rect 265360 137714 265388 150418
rect 265268 137686 265388 137714
rect 265268 125769 265296 137686
rect 265254 125760 265310 125769
rect 265254 125695 265310 125704
rect 265254 125624 265310 125633
rect 265254 125559 265310 125568
rect 265268 114578 265296 125559
rect 265164 114572 265216 114578
rect 265164 114514 265216 114520
rect 265256 114572 265308 114578
rect 265256 114514 265308 114520
rect 265176 109070 265204 114514
rect 265164 109064 265216 109070
rect 265164 109006 265216 109012
rect 265256 108996 265308 109002
rect 265256 108938 265308 108944
rect 265268 95334 265296 108938
rect 265256 95328 265308 95334
rect 265256 95270 265308 95276
rect 265256 92540 265308 92546
rect 265256 92482 265308 92488
rect 265268 67658 265296 92482
rect 265164 67652 265216 67658
rect 265164 67594 265216 67600
rect 265256 67652 265308 67658
rect 265256 67594 265308 67600
rect 265176 66230 265204 67594
rect 265164 66224 265216 66230
rect 265164 66166 265216 66172
rect 265164 50924 265216 50930
rect 265164 50866 265216 50872
rect 265176 46918 265204 50866
rect 265164 46912 265216 46918
rect 265164 46854 265216 46860
rect 265164 37324 265216 37330
rect 265164 37266 265216 37272
rect 265176 29034 265204 37266
rect 265164 29028 265216 29034
rect 265164 28970 265216 28976
rect 265256 29028 265308 29034
rect 265256 28970 265308 28976
rect 265268 27606 265296 28970
rect 265256 27600 265308 27606
rect 265256 27542 265308 27548
rect 265622 16960 265678 16969
rect 265622 16895 265678 16904
rect 265636 16425 265664 16895
rect 265622 16416 265678 16425
rect 265622 16351 265678 16360
rect 266464 14822 266492 335582
rect 266740 335566 266952 335594
rect 267372 335640 267424 335646
rect 268396 335594 268424 340054
rect 269028 337408 269080 337414
rect 269028 337350 269080 337356
rect 267372 335582 267424 335588
rect 267844 335566 268424 335594
rect 266740 321638 266768 335566
rect 267844 321638 267872 335566
rect 266728 321632 266780 321638
rect 266728 321574 266780 321580
rect 267832 321632 267884 321638
rect 267832 321574 267884 321580
rect 266636 318844 266688 318850
rect 266636 318786 266688 318792
rect 267740 318844 267792 318850
rect 267740 318786 267792 318792
rect 266648 309262 266676 318786
rect 267752 315994 267780 318786
rect 267740 315988 267792 315994
rect 267740 315930 267792 315936
rect 267832 311160 267884 311166
rect 267832 311102 267884 311108
rect 266636 309256 266688 309262
rect 266636 309198 266688 309204
rect 267844 306377 267872 311102
rect 267830 306368 267886 306377
rect 267830 306303 267886 306312
rect 268014 306368 268070 306377
rect 268014 306303 268070 306312
rect 266636 305040 266688 305046
rect 266636 304982 266688 304988
rect 266648 299538 266676 304982
rect 266636 299532 266688 299538
rect 266636 299474 266688 299480
rect 266728 299532 266780 299538
rect 266728 299474 266780 299480
rect 266740 298110 266768 299474
rect 266728 298104 266780 298110
rect 266728 298046 266780 298052
rect 268028 296750 268056 306303
rect 267740 296744 267792 296750
rect 267740 296686 267792 296692
rect 268016 296744 268068 296750
rect 268016 296686 268068 296692
rect 267752 296614 267780 296686
rect 267740 296608 267792 296614
rect 267740 296550 267792 296556
rect 266820 288448 266872 288454
rect 266820 288390 266872 288396
rect 266832 280226 266860 288390
rect 267740 287088 267792 287094
rect 267740 287030 267792 287036
rect 266728 280220 266780 280226
rect 266728 280162 266780 280168
rect 266820 280220 266872 280226
rect 266820 280162 266872 280168
rect 266740 263634 266768 280162
rect 267752 269113 267780 287030
rect 267738 269104 267794 269113
rect 267738 269039 267794 269048
rect 267830 268968 267886 268977
rect 267830 268903 267886 268912
rect 266728 263628 266780 263634
rect 266728 263570 266780 263576
rect 266740 259486 266768 259517
rect 266728 259480 266780 259486
rect 266648 259428 266728 259434
rect 266648 259422 266780 259428
rect 266648 259406 266768 259422
rect 266648 241534 266676 259406
rect 266636 241528 266688 241534
rect 266636 241470 266688 241476
rect 266728 241528 266780 241534
rect 266728 241470 266780 241476
rect 266740 235362 266768 241470
rect 267844 240174 267872 268903
rect 267740 240168 267792 240174
rect 267740 240110 267792 240116
rect 267832 240168 267884 240174
rect 267832 240110 267884 240116
rect 266740 235334 266860 235362
rect 266832 220833 266860 235334
rect 267752 234734 267780 240110
rect 267740 234728 267792 234734
rect 267740 234670 267792 234676
rect 267740 234592 267792 234598
rect 267740 234534 267792 234540
rect 267752 222193 267780 234534
rect 267738 222184 267794 222193
rect 267738 222119 267794 222128
rect 267738 222048 267794 222057
rect 267738 221983 267794 221992
rect 266634 220824 266690 220833
rect 266634 220759 266690 220768
rect 266818 220824 266874 220833
rect 266818 220759 266874 220768
rect 266648 215914 266676 220759
rect 266648 215886 266768 215914
rect 266740 198150 266768 215886
rect 267752 212548 267780 221983
rect 267752 212520 267872 212548
rect 267844 202892 267872 212520
rect 267752 202881 267872 202892
rect 267738 202872 267872 202881
rect 267794 202864 267872 202872
rect 267922 202872 267978 202881
rect 267738 202807 267794 202816
rect 267922 202807 267978 202816
rect 266728 198144 266780 198150
rect 266728 198086 266780 198092
rect 266728 198008 266780 198014
rect 266728 197950 266780 197956
rect 266740 193236 266768 197950
rect 267936 193254 267964 202807
rect 266648 193208 266768 193236
rect 267832 193248 267884 193254
rect 266648 186386 266676 193208
rect 267832 193190 267884 193196
rect 267924 193248 267976 193254
rect 267924 193190 267976 193196
rect 267844 190466 267872 193190
rect 267740 190460 267792 190466
rect 267740 190402 267792 190408
rect 267832 190460 267884 190466
rect 267832 190402 267884 190408
rect 266636 186380 266688 186386
rect 266636 186322 266688 186328
rect 266728 186244 266780 186250
rect 266728 186186 266780 186192
rect 266740 178838 266768 186186
rect 267752 180849 267780 190402
rect 267738 180840 267794 180849
rect 267922 180840 267978 180849
rect 267738 180775 267794 180784
rect 267832 180804 267884 180810
rect 267922 180775 267924 180784
rect 267832 180746 267884 180752
rect 267976 180775 267978 180784
rect 267924 180746 267976 180752
rect 267844 179382 267872 180746
rect 267832 179376 267884 179382
rect 267832 179318 267884 179324
rect 266728 178832 266780 178838
rect 266728 178774 266780 178780
rect 266728 178696 266780 178702
rect 266728 178638 266780 178644
rect 266740 173924 266768 178638
rect 266648 173896 266768 173924
rect 266648 171086 266676 173896
rect 266636 171080 266688 171086
rect 266636 171022 266688 171028
rect 267832 169788 267884 169794
rect 267832 169730 267884 169736
rect 267844 161514 267872 169730
rect 266820 161492 266872 161498
rect 266820 161434 266872 161440
rect 267752 161486 267872 161514
rect 266832 151842 266860 161434
rect 267752 157486 267780 161486
rect 267740 157480 267792 157486
rect 267740 157422 267792 157428
rect 267740 157344 267792 157350
rect 267740 157286 267792 157292
rect 266820 151836 266872 151842
rect 266820 151778 266872 151784
rect 266820 151700 266872 151706
rect 266820 151642 266872 151648
rect 266832 139890 266860 151642
rect 267752 144906 267780 157286
rect 267740 144900 267792 144906
rect 267740 144842 267792 144848
rect 267924 144900 267976 144906
rect 267924 144842 267976 144848
rect 267936 139890 267964 144842
rect 266740 139862 266860 139890
rect 267844 139862 267964 139890
rect 266740 125769 266768 139862
rect 267646 134600 267702 134609
rect 267646 134535 267702 134544
rect 267660 134337 267688 134535
rect 267646 134328 267702 134337
rect 267646 134263 267702 134272
rect 267844 125769 267872 139862
rect 266726 125760 266782 125769
rect 266726 125695 266782 125704
rect 267830 125760 267886 125769
rect 267830 125695 267886 125704
rect 266634 125624 266690 125633
rect 266634 125559 266690 125568
rect 267738 125624 267794 125633
rect 267738 125559 267794 125568
rect 266648 77314 266676 125559
rect 267648 110628 267700 110634
rect 267648 110570 267700 110576
rect 267660 110537 267688 110570
rect 267646 110528 267702 110537
rect 267646 110463 267702 110472
rect 267752 104922 267780 125559
rect 267740 104916 267792 104922
rect 267740 104858 267792 104864
rect 267832 104916 267884 104922
rect 267832 104858 267884 104864
rect 267844 99482 267872 104858
rect 267832 99476 267884 99482
rect 267832 99418 267884 99424
rect 267740 99340 267792 99346
rect 267740 99282 267792 99288
rect 267752 85610 267780 99282
rect 267740 85604 267792 85610
rect 267740 85546 267792 85552
rect 267832 85468 267884 85474
rect 267832 85410 267884 85416
rect 267844 82822 267872 85410
rect 267832 82816 267884 82822
rect 267832 82758 267884 82764
rect 266636 77308 266688 77314
rect 266636 77250 266688 77256
rect 266728 77308 266780 77314
rect 266728 77250 266780 77256
rect 266740 67674 266768 77250
rect 267924 73228 267976 73234
rect 267924 73170 267976 73176
rect 266648 67646 266768 67674
rect 266648 60790 266676 67646
rect 267936 65006 267964 73170
rect 267924 65000 267976 65006
rect 267924 64942 267976 64948
rect 267740 64932 267792 64938
rect 267740 64874 267792 64880
rect 267752 60858 267780 64874
rect 267740 60852 267792 60858
rect 267740 60794 267792 60800
rect 266636 60784 266688 60790
rect 266636 60726 266688 60732
rect 267740 60716 267792 60722
rect 267740 60658 267792 60664
rect 266728 60648 266780 60654
rect 266728 60590 266780 60596
rect 266740 46918 266768 60590
rect 267752 48385 267780 60658
rect 267738 48376 267794 48385
rect 267738 48311 267794 48320
rect 267922 48240 267978 48249
rect 267922 48175 267978 48184
rect 266728 46912 266780 46918
rect 266728 46854 266780 46860
rect 267936 38758 267964 48175
rect 267924 38752 267976 38758
rect 267924 38694 267976 38700
rect 267924 38616 267976 38622
rect 267924 38558 267976 38564
rect 266728 37324 266780 37330
rect 266728 37266 266780 37272
rect 266740 19446 266768 37266
rect 267936 29034 267964 38558
rect 267832 29028 267884 29034
rect 267832 28970 267884 28976
rect 267924 29028 267976 29034
rect 267924 28970 267976 28976
rect 267844 22642 267872 28970
rect 267832 22636 267884 22642
rect 267832 22578 267884 22584
rect 266728 19440 266780 19446
rect 266728 19382 266780 19388
rect 266636 19304 266688 19310
rect 266636 19246 266688 19252
rect 266452 14816 266504 14822
rect 266452 14758 266504 14764
rect 265072 14748 265124 14754
rect 265072 14690 265124 14696
rect 266648 10606 266676 19246
rect 266636 10600 266688 10606
rect 266636 10542 266688 10548
rect 264978 8392 265034 8401
rect 264978 8327 265034 8336
rect 265162 8392 265218 8401
rect 265162 8327 265218 8336
rect 265176 8294 265204 8327
rect 265164 8288 265216 8294
rect 265164 8230 265216 8236
rect 263876 8220 263928 8226
rect 263876 8162 263928 8168
rect 267004 8220 267056 8226
rect 267004 8162 267056 8168
rect 262404 8152 262456 8158
rect 262404 8094 262456 8100
rect 263416 8152 263468 8158
rect 263416 8094 263468 8100
rect 262220 3664 262272 3670
rect 262220 3606 262272 3612
rect 261484 2848 261536 2854
rect 261484 2790 261536 2796
rect 261024 1148 261076 1154
rect 261024 1090 261076 1096
rect 261036 480 261064 1090
rect 262232 480 262260 3606
rect 263428 480 263456 8094
rect 264612 3868 264664 3874
rect 264612 3810 264664 3816
rect 264624 480 264652 3810
rect 265808 3596 265860 3602
rect 265808 3538 265860 3544
rect 265820 480 265848 3538
rect 267016 480 267044 8162
rect 269040 4146 269068 337350
rect 269224 14890 269252 340054
rect 269684 337482 269712 340068
rect 269868 340054 270158 340082
rect 269672 337476 269724 337482
rect 269672 337418 269724 337424
rect 269868 335594 269896 340054
rect 269316 335566 269896 335594
rect 269212 14884 269264 14890
rect 269212 14826 269264 14832
rect 269316 10742 269344 335566
rect 270498 212528 270554 212537
rect 270498 212463 270554 212472
rect 270512 202910 270540 212463
rect 270500 202904 270552 202910
rect 270498 202872 270500 202881
rect 270552 202872 270554 202881
rect 270498 202807 270554 202816
rect 270512 193254 270540 202807
rect 270500 193248 270552 193254
rect 270498 193216 270500 193225
rect 270552 193216 270554 193225
rect 270498 193151 270554 193160
rect 270512 183598 270540 193151
rect 270500 183592 270552 183598
rect 270498 183560 270500 183569
rect 270552 183560 270554 183569
rect 270498 183495 270554 183504
rect 270512 173942 270540 183495
rect 270500 173936 270552 173942
rect 270500 173878 270552 173884
rect 270314 134328 270370 134337
rect 270498 134328 270554 134337
rect 270370 134286 270498 134314
rect 270314 134263 270370 134272
rect 270498 134263 270554 134272
rect 270500 76016 270552 76022
rect 270498 75984 270500 75993
rect 270552 75984 270554 75993
rect 270498 75919 270554 75928
rect 270406 40216 270462 40225
rect 270406 40151 270462 40160
rect 270420 40089 270448 40151
rect 270406 40080 270462 40089
rect 270406 40015 270462 40024
rect 269856 22160 269908 22166
rect 269856 22102 269908 22108
rect 269868 10810 269896 22102
rect 270604 14958 270632 340068
rect 271156 337142 271184 340068
rect 271248 340054 271630 340082
rect 271984 340054 272090 340082
rect 271144 337136 271196 337142
rect 271144 337078 271196 337084
rect 271248 334354 271276 340054
rect 271328 337272 271380 337278
rect 271328 337214 271380 337220
rect 270776 334348 270828 334354
rect 270776 334290 270828 334296
rect 271236 334348 271288 334354
rect 271236 334290 271288 334296
rect 270788 317422 270816 334290
rect 271340 334234 271368 337214
rect 271788 337204 271840 337210
rect 271788 337146 271840 337152
rect 271156 334206 271368 334234
rect 270776 317416 270828 317422
rect 270776 317358 270828 317364
rect 270776 307828 270828 307834
rect 270776 307770 270828 307776
rect 270788 299470 270816 307770
rect 270776 299464 270828 299470
rect 270776 299406 270828 299412
rect 270776 289876 270828 289882
rect 270776 289818 270828 289824
rect 270788 283014 270816 289818
rect 270776 283008 270828 283014
rect 270776 282950 270828 282956
rect 270684 282872 270736 282878
rect 270684 282814 270736 282820
rect 270696 280158 270724 282814
rect 270684 280152 270736 280158
rect 270684 280094 270736 280100
rect 270684 275324 270736 275330
rect 270684 275266 270736 275272
rect 270696 263634 270724 275266
rect 270684 263628 270736 263634
rect 270684 263570 270736 263576
rect 270684 263492 270736 263498
rect 270684 263434 270736 263440
rect 270696 260846 270724 263434
rect 270684 260840 270736 260846
rect 270684 260782 270736 260788
rect 270684 256012 270736 256018
rect 270684 255954 270736 255960
rect 270696 241466 270724 255954
rect 270684 241460 270736 241466
rect 270684 241402 270736 241408
rect 270868 241460 270920 241466
rect 270868 241402 270920 241408
rect 270880 240122 270908 241402
rect 270788 240094 270908 240122
rect 270788 230518 270816 240094
rect 270684 230512 270736 230518
rect 270684 230454 270736 230460
rect 270776 230512 270828 230518
rect 270776 230454 270828 230460
rect 270696 225010 270724 230454
rect 270684 225004 270736 225010
rect 270684 224946 270736 224952
rect 270684 224868 270736 224874
rect 270684 224810 270736 224816
rect 270696 222154 270724 224810
rect 270684 222148 270736 222154
rect 270684 222090 270736 222096
rect 270776 212560 270828 212566
rect 270774 212528 270776 212537
rect 270828 212528 270830 212537
rect 270774 212463 270830 212472
rect 270684 202904 270736 202910
rect 270682 202872 270684 202881
rect 270736 202872 270738 202881
rect 270682 202807 270738 202816
rect 270776 193248 270828 193254
rect 270774 193216 270776 193225
rect 270828 193216 270830 193225
rect 270774 193151 270830 193160
rect 270684 183592 270736 183598
rect 270682 183560 270684 183569
rect 270736 183560 270738 183569
rect 270682 183495 270738 183504
rect 270776 173936 270828 173942
rect 270776 173878 270828 173884
rect 270788 169130 270816 173878
rect 270696 169102 270816 169130
rect 270696 164218 270724 169102
rect 270684 164212 270736 164218
rect 270684 164154 270736 164160
rect 270776 164144 270828 164150
rect 270776 164086 270828 164092
rect 270788 153202 270816 164086
rect 270776 153196 270828 153202
rect 270776 153138 270828 153144
rect 270868 153196 270920 153202
rect 270868 153138 270920 153144
rect 270880 137850 270908 153138
rect 270788 137822 270908 137850
rect 270788 133890 270816 137822
rect 270776 133884 270828 133890
rect 270776 133826 270828 133832
rect 271052 133884 271104 133890
rect 271052 133826 271104 133832
rect 271064 124250 271092 133826
rect 270880 124222 271092 124250
rect 270880 122806 270908 124222
rect 270868 122800 270920 122806
rect 270868 122742 270920 122748
rect 270776 113212 270828 113218
rect 270776 113154 270828 113160
rect 270788 104922 270816 113154
rect 270684 104916 270736 104922
rect 270684 104858 270736 104864
rect 270776 104916 270828 104922
rect 270776 104858 270828 104864
rect 270696 95266 270724 104858
rect 270684 95260 270736 95266
rect 270684 95202 270736 95208
rect 270776 95260 270828 95266
rect 270776 95202 270828 95208
rect 270788 90438 270816 95202
rect 270776 90432 270828 90438
rect 270776 90374 270828 90380
rect 270776 77308 270828 77314
rect 270776 77250 270828 77256
rect 270788 70514 270816 77250
rect 270776 70508 270828 70514
rect 270776 70450 270828 70456
rect 270684 70372 270736 70378
rect 270684 70314 270736 70320
rect 270696 58070 270724 70314
rect 270684 58064 270736 58070
rect 270684 58006 270736 58012
rect 270684 57928 270736 57934
rect 270684 57870 270736 57876
rect 270696 38690 270724 57870
rect 270684 38684 270736 38690
rect 270684 38626 270736 38632
rect 270776 38684 270828 38690
rect 270776 38626 270828 38632
rect 270788 37262 270816 38626
rect 270776 37256 270828 37262
rect 270776 37198 270828 37204
rect 270868 37256 270920 37262
rect 270868 37198 270920 37204
rect 270880 35902 270908 37198
rect 270868 35896 270920 35902
rect 270868 35838 270920 35844
rect 270776 26308 270828 26314
rect 270776 26250 270828 26256
rect 270788 26194 270816 26250
rect 270696 26166 270816 26194
rect 270696 22166 270724 26166
rect 270684 22160 270736 22166
rect 270684 22102 270736 22108
rect 270592 14952 270644 14958
rect 270592 14894 270644 14900
rect 269856 10804 269908 10810
rect 269856 10746 269908 10752
rect 269304 10736 269356 10742
rect 269304 10678 269356 10684
rect 270500 8288 270552 8294
rect 270500 8230 270552 8236
rect 268108 4140 268160 4146
rect 268108 4082 268160 4088
rect 269028 4140 269080 4146
rect 269028 4082 269080 4088
rect 268120 480 268148 4082
rect 269304 3256 269356 3262
rect 269304 3198 269356 3204
rect 269316 480 269344 3198
rect 270512 480 270540 8230
rect 271156 4418 271184 334206
rect 271144 4412 271196 4418
rect 271144 4354 271196 4360
rect 271800 626 271828 337146
rect 271984 15026 272012 340054
rect 272628 337890 272656 340068
rect 272720 340054 273102 340082
rect 273364 340054 273562 340082
rect 272616 337884 272668 337890
rect 272616 337826 272668 337832
rect 272720 334354 272748 340054
rect 272800 337340 272852 337346
rect 272800 337282 272852 337288
rect 272248 334348 272300 334354
rect 272248 334290 272300 334296
rect 272708 334348 272760 334354
rect 272708 334290 272760 334296
rect 272260 317422 272288 334290
rect 272812 334234 272840 337282
rect 272536 334206 272840 334234
rect 272248 317416 272300 317422
rect 272248 317358 272300 317364
rect 272248 307828 272300 307834
rect 272248 307770 272300 307776
rect 272260 299470 272288 307770
rect 272248 299464 272300 299470
rect 272248 299406 272300 299412
rect 272248 289332 272300 289338
rect 272248 289274 272300 289280
rect 272260 288386 272288 289274
rect 272248 288380 272300 288386
rect 272248 288322 272300 288328
rect 272340 288380 272392 288386
rect 272340 288322 272392 288328
rect 272352 278769 272380 288322
rect 272154 278760 272210 278769
rect 272154 278695 272210 278704
rect 272338 278760 272394 278769
rect 272338 278695 272394 278704
rect 272168 270042 272196 278695
rect 272168 270014 272380 270042
rect 272352 260982 272380 270014
rect 272340 260976 272392 260982
rect 272340 260918 272392 260924
rect 272156 260772 272208 260778
rect 272156 260714 272208 260720
rect 272168 241466 272196 260714
rect 272156 241460 272208 241466
rect 272156 241402 272208 241408
rect 272340 241460 272392 241466
rect 272340 241402 272392 241408
rect 272352 240145 272380 241402
rect 272154 240136 272210 240145
rect 272154 240071 272210 240080
rect 272338 240136 272394 240145
rect 272338 240071 272394 240080
rect 272168 231554 272196 240071
rect 272168 231526 272380 231554
rect 272352 224890 272380 231526
rect 272168 224862 272380 224890
rect 272168 222154 272196 224862
rect 272156 222148 272208 222154
rect 272156 222090 272208 222096
rect 272248 222148 272300 222154
rect 272248 222090 272300 222096
rect 272260 220833 272288 222090
rect 272062 220824 272118 220833
rect 272062 220759 272118 220768
rect 272246 220824 272302 220833
rect 272246 220759 272302 220768
rect 272076 211177 272104 220759
rect 272062 211168 272118 211177
rect 272062 211103 272118 211112
rect 272246 211168 272302 211177
rect 272246 211103 272302 211112
rect 272260 207754 272288 211103
rect 272076 207726 272288 207754
rect 272076 205578 272104 207726
rect 272076 205550 272196 205578
rect 272168 202881 272196 205550
rect 272154 202872 272210 202881
rect 272154 202807 272210 202816
rect 272338 202736 272394 202745
rect 272338 202671 272394 202680
rect 272352 193202 272380 202671
rect 272076 193174 272380 193202
rect 272076 186266 272104 193174
rect 272076 186238 272196 186266
rect 272168 183569 272196 186238
rect 272154 183560 272210 183569
rect 272154 183495 272210 183504
rect 272338 183424 272394 183433
rect 272338 183359 272394 183368
rect 272352 182170 272380 183359
rect 272064 182164 272116 182170
rect 272064 182106 272116 182112
rect 272340 182164 272392 182170
rect 272340 182106 272392 182112
rect 272076 172553 272104 182106
rect 272062 172544 272118 172553
rect 272062 172479 272118 172488
rect 272246 172544 272302 172553
rect 272246 172479 272302 172488
rect 272260 166274 272288 172479
rect 272168 166246 272288 166274
rect 272168 160070 272196 166246
rect 272156 160064 272208 160070
rect 272156 160006 272208 160012
rect 272340 148300 272392 148306
rect 272340 148242 272392 148248
rect 272352 139890 272380 148242
rect 272260 139862 272380 139890
rect 272260 125769 272288 139862
rect 272246 125760 272302 125769
rect 272246 125695 272302 125704
rect 272154 125624 272210 125633
rect 272154 125559 272210 125568
rect 272168 119354 272196 125559
rect 272168 119326 272288 119354
rect 272260 114510 272288 119326
rect 272248 114504 272300 114510
rect 272248 114446 272300 114452
rect 272340 114504 272392 114510
rect 272340 114446 272392 114452
rect 272352 95334 272380 114446
rect 272340 95328 272392 95334
rect 272340 95270 272392 95276
rect 272248 95260 272300 95266
rect 272248 95202 272300 95208
rect 272260 90438 272288 95202
rect 272248 90432 272300 90438
rect 272248 90374 272300 90380
rect 272248 77308 272300 77314
rect 272248 77250 272300 77256
rect 272260 70582 272288 77250
rect 272248 70576 272300 70582
rect 272248 70518 272300 70524
rect 272156 67652 272208 67658
rect 272156 67594 272208 67600
rect 272168 58002 272196 67594
rect 272156 57996 272208 58002
rect 272156 57938 272208 57944
rect 272248 57996 272300 58002
rect 272248 57938 272300 57944
rect 272260 53122 272288 57938
rect 272168 53094 272288 53122
rect 272168 38690 272196 53094
rect 272156 38684 272208 38690
rect 272156 38626 272208 38632
rect 272248 38684 272300 38690
rect 272248 38626 272300 38632
rect 272260 26246 272288 38626
rect 272248 26240 272300 26246
rect 272248 26182 272300 26188
rect 271972 15020 272024 15026
rect 271972 14962 272024 14968
rect 272536 4350 272564 334206
rect 273074 87136 273130 87145
rect 273258 87136 273314 87145
rect 273130 87094 273258 87122
rect 273074 87071 273130 87080
rect 273258 87071 273314 87080
rect 273074 29200 273130 29209
rect 273258 29200 273314 29209
rect 273130 29158 273258 29186
rect 273074 29135 273130 29144
rect 273258 29135 273314 29144
rect 273364 15094 273392 340054
rect 274100 337006 274128 340068
rect 274284 340054 274574 340082
rect 274744 340054 275034 340082
rect 274088 337000 274140 337006
rect 274088 336942 274140 336948
rect 274284 331242 274312 340054
rect 273548 331214 274312 331242
rect 273548 321774 273576 331214
rect 273536 321768 273588 321774
rect 273536 321710 273588 321716
rect 273536 317552 273588 317558
rect 273536 317494 273588 317500
rect 273548 317422 273576 317494
rect 273536 317416 273588 317422
rect 273536 317358 273588 317364
rect 273628 317348 273680 317354
rect 273628 317290 273680 317296
rect 273640 309074 273668 317290
rect 273548 309046 273668 309074
rect 273548 299470 273576 309046
rect 273536 299464 273588 299470
rect 273536 299406 273588 299412
rect 273536 299328 273588 299334
rect 273536 299270 273588 299276
rect 273548 280158 273576 299270
rect 273536 280152 273588 280158
rect 273536 280094 273588 280100
rect 273536 270564 273588 270570
rect 273536 270506 273588 270512
rect 273548 260846 273576 270506
rect 273536 260840 273588 260846
rect 273536 260782 273588 260788
rect 273536 251252 273588 251258
rect 273536 251194 273588 251200
rect 273548 241505 273576 251194
rect 273534 241496 273590 241505
rect 273534 241431 273590 241440
rect 273718 241496 273774 241505
rect 273718 241431 273774 241440
rect 273732 231878 273760 241431
rect 273536 231872 273588 231878
rect 273536 231814 273588 231820
rect 273720 231872 273772 231878
rect 273720 231814 273772 231820
rect 273548 222193 273576 231814
rect 273534 222184 273590 222193
rect 273534 222119 273590 222128
rect 273718 222184 273774 222193
rect 273718 222119 273774 222128
rect 273732 212566 273760 222119
rect 273536 212560 273588 212566
rect 273536 212502 273588 212508
rect 273720 212560 273772 212566
rect 273720 212502 273772 212508
rect 273548 202881 273576 212502
rect 273534 202872 273590 202881
rect 273534 202807 273590 202816
rect 273718 202872 273774 202881
rect 273718 202807 273774 202816
rect 273732 193254 273760 202807
rect 273536 193248 273588 193254
rect 273536 193190 273588 193196
rect 273720 193248 273772 193254
rect 273720 193190 273772 193196
rect 273548 183569 273576 193190
rect 273534 183560 273590 183569
rect 273534 183495 273590 183504
rect 273718 183560 273774 183569
rect 273718 183495 273774 183504
rect 273732 182170 273760 183495
rect 273720 182164 273772 182170
rect 273720 182106 273772 182112
rect 273536 172576 273588 172582
rect 273536 172518 273588 172524
rect 273548 153202 273576 172518
rect 273536 153196 273588 153202
rect 273536 153138 273588 153144
rect 273536 144900 273588 144906
rect 273536 144842 273588 144848
rect 273548 143562 273576 144842
rect 273548 143534 273668 143562
rect 273640 135318 273668 143534
rect 273536 135312 273588 135318
rect 273536 135254 273588 135260
rect 273628 135312 273680 135318
rect 273628 135254 273680 135260
rect 273548 125769 273576 135254
rect 273534 125760 273590 125769
rect 273534 125695 273590 125704
rect 273534 125624 273590 125633
rect 273534 125559 273590 125568
rect 273548 118810 273576 125559
rect 273718 123312 273774 123321
rect 273902 123312 273958 123321
rect 273774 123270 273902 123298
rect 273718 123247 273774 123256
rect 273902 123247 273958 123256
rect 273548 118782 273668 118810
rect 273640 118538 273668 118782
rect 273548 118510 273668 118538
rect 273548 99498 273576 118510
rect 273456 99470 273576 99498
rect 273456 99362 273484 99470
rect 273456 99334 273576 99362
rect 273548 80034 273576 99334
rect 273536 80028 273588 80034
rect 273536 79970 273588 79976
rect 273536 75948 273588 75954
rect 273536 75890 273588 75896
rect 273548 66230 273576 75890
rect 273536 66224 273588 66230
rect 273536 66166 273588 66172
rect 273536 56636 273588 56642
rect 273536 56578 273588 56584
rect 273548 51134 273576 56578
rect 273536 51128 273588 51134
rect 273536 51070 273588 51076
rect 273536 50924 273588 50930
rect 273536 50866 273588 50872
rect 273548 22114 273576 50866
rect 273456 22086 273576 22114
rect 273456 17950 273484 22086
rect 273444 17944 273496 17950
rect 273444 17886 273496 17892
rect 274744 15162 274772 340054
rect 275572 337550 275600 340068
rect 275560 337544 275612 337550
rect 275560 337486 275612 337492
rect 275928 337544 275980 337550
rect 275928 337486 275980 337492
rect 275374 76120 275430 76129
rect 275374 76055 275430 76064
rect 275388 76022 275416 76055
rect 275376 76016 275428 76022
rect 275376 75958 275428 75964
rect 274732 15156 274784 15162
rect 274732 15098 274784 15104
rect 273352 15088 273404 15094
rect 273352 15030 273404 15036
rect 274088 6180 274140 6186
rect 274088 6122 274140 6128
rect 272524 4344 272576 4350
rect 272524 4286 272576 4292
rect 272892 3188 272944 3194
rect 272892 3130 272944 3136
rect 271708 598 271828 626
rect 271708 480 271736 598
rect 272904 480 272932 3130
rect 274100 480 274128 6122
rect 275940 2922 275968 337486
rect 276032 11014 276060 340068
rect 276124 340054 276506 340082
rect 276124 14414 276152 340054
rect 277044 337686 277072 340068
rect 277518 340054 277624 340082
rect 277032 337680 277084 337686
rect 277032 337622 277084 337628
rect 276112 14408 276164 14414
rect 276112 14350 276164 14356
rect 276020 11008 276072 11014
rect 276020 10950 276072 10956
rect 277596 10266 277624 340054
rect 277688 340054 277978 340082
rect 277688 14346 277716 340054
rect 278516 336870 278544 340068
rect 278884 340054 278990 340082
rect 279068 340054 279450 340082
rect 278504 336864 278556 336870
rect 278504 336806 278556 336812
rect 278884 335442 278912 340054
rect 278872 335436 278924 335442
rect 278872 335378 278924 335384
rect 278964 335232 279016 335238
rect 278964 335174 279016 335180
rect 278872 333328 278924 333334
rect 278872 333270 278924 333276
rect 278884 302274 278912 333270
rect 278792 302246 278912 302274
rect 278792 302138 278820 302246
rect 278792 302110 278912 302138
rect 278884 282962 278912 302110
rect 278792 282934 278912 282962
rect 278792 282826 278820 282934
rect 278792 282798 278912 282826
rect 278884 263650 278912 282798
rect 278792 263622 278912 263650
rect 278792 263514 278820 263622
rect 278792 263486 278912 263514
rect 278884 244338 278912 263486
rect 278792 244310 278912 244338
rect 278792 244202 278820 244310
rect 278792 244174 278912 244202
rect 278884 225026 278912 244174
rect 278792 224998 278912 225026
rect 278792 224890 278820 224998
rect 278792 224862 278912 224890
rect 278884 205714 278912 224862
rect 278792 205686 278912 205714
rect 278792 205578 278820 205686
rect 278792 205550 278912 205578
rect 278884 186402 278912 205550
rect 278792 186374 278912 186402
rect 278792 186266 278820 186374
rect 278792 186238 278912 186266
rect 278884 167074 278912 186238
rect 278872 167068 278924 167074
rect 278872 167010 278924 167016
rect 278780 166932 278832 166938
rect 278780 166874 278832 166880
rect 278792 140026 278820 166874
rect 278792 139998 278912 140026
rect 278884 118794 278912 139998
rect 278872 118788 278924 118794
rect 278872 118730 278924 118736
rect 278872 118652 278924 118658
rect 278872 118594 278924 118600
rect 278884 80170 278912 118594
rect 278872 80164 278924 80170
rect 278872 80106 278924 80112
rect 278872 80028 278924 80034
rect 278872 79970 278924 79976
rect 278884 51202 278912 79970
rect 278872 51196 278924 51202
rect 278872 51138 278924 51144
rect 278872 48340 278924 48346
rect 278872 48282 278924 48288
rect 278884 31770 278912 48282
rect 278792 31742 278912 31770
rect 277676 14340 277728 14346
rect 277676 14282 277728 14288
rect 278792 14278 278820 31742
rect 278780 14272 278832 14278
rect 278780 14214 278832 14220
rect 277584 10260 277636 10266
rect 277584 10202 277636 10208
rect 278976 10198 279004 335174
rect 279068 333334 279096 340054
rect 279988 337618 280016 340068
rect 280356 340054 280462 340082
rect 280632 340054 280922 340082
rect 281184 340054 281474 340082
rect 281552 340054 281934 340082
rect 279976 337612 280028 337618
rect 279976 337554 280028 337560
rect 280252 335640 280304 335646
rect 280252 335582 280304 335588
rect 279056 333328 279108 333334
rect 279056 333270 279108 333276
rect 280264 14210 280292 335582
rect 280252 14204 280304 14210
rect 280252 14146 280304 14152
rect 278964 10192 279016 10198
rect 278964 10134 279016 10140
rect 280356 10130 280384 340054
rect 280632 335646 280660 340054
rect 281184 336802 281212 340054
rect 281448 337612 281500 337618
rect 281448 337554 281500 337560
rect 281172 336796 281224 336802
rect 281172 336738 281224 336744
rect 280620 335640 280672 335646
rect 280620 335582 280672 335588
rect 280344 10124 280396 10130
rect 280344 10066 280396 10072
rect 280068 6248 280120 6254
rect 280068 6190 280120 6196
rect 278872 3800 278924 3806
rect 278872 3742 278924 3748
rect 276480 3256 276532 3262
rect 276480 3198 276532 3204
rect 275284 2916 275336 2922
rect 275284 2858 275336 2864
rect 275928 2916 275980 2922
rect 275928 2858 275980 2864
rect 275296 480 275324 2858
rect 276492 480 276520 3198
rect 277676 3188 277728 3194
rect 277676 3130 277728 3136
rect 277688 480 277716 3130
rect 278884 480 278912 3742
rect 280080 480 280108 6190
rect 281460 610 281488 337554
rect 281552 11830 281580 340054
rect 282012 335628 282040 340190
rect 282946 340054 283144 340082
rect 281828 335600 282040 335628
rect 283012 335640 283064 335646
rect 281828 321638 281856 335600
rect 283012 335582 283064 335588
rect 281816 321632 281868 321638
rect 281816 321574 281868 321580
rect 281724 316056 281776 316062
rect 281724 315998 281776 316004
rect 281736 311250 281764 315998
rect 281736 311222 281856 311250
rect 281828 299470 281856 311222
rect 281724 299464 281776 299470
rect 281724 299406 281776 299412
rect 281816 299464 281868 299470
rect 281816 299406 281868 299412
rect 281736 298110 281764 299406
rect 281724 298104 281776 298110
rect 281724 298046 281776 298052
rect 281816 298104 281868 298110
rect 281816 298046 281868 298052
rect 281828 280158 281856 298046
rect 281724 280152 281776 280158
rect 281724 280094 281776 280100
rect 281816 280152 281868 280158
rect 281816 280094 281868 280100
rect 281736 278769 281764 280094
rect 281722 278760 281778 278769
rect 281722 278695 281778 278704
rect 281814 278624 281870 278633
rect 281814 278559 281870 278568
rect 281828 260914 281856 278559
rect 281816 260908 281868 260914
rect 281816 260850 281868 260856
rect 281816 259480 281868 259486
rect 281816 259422 281868 259428
rect 281828 251190 281856 259422
rect 281816 251184 281868 251190
rect 281816 251126 281868 251132
rect 281816 241528 281868 241534
rect 281816 241470 281868 241476
rect 281828 234734 281856 241470
rect 281816 234728 281868 234734
rect 281816 234670 281868 234676
rect 281816 234592 281868 234598
rect 281816 234534 281868 234540
rect 281828 217410 281856 234534
rect 281828 217382 281948 217410
rect 281920 212566 281948 217382
rect 281724 212560 281776 212566
rect 281724 212502 281776 212508
rect 281908 212560 281960 212566
rect 281908 212502 281960 212508
rect 281736 205698 281764 212502
rect 281724 205692 281776 205698
rect 281724 205634 281776 205640
rect 281816 205556 281868 205562
rect 281816 205498 281868 205504
rect 281828 198098 281856 205498
rect 281828 198070 281948 198098
rect 281920 193254 281948 198070
rect 281724 193248 281776 193254
rect 281722 193216 281724 193225
rect 281908 193248 281960 193254
rect 281776 193216 281778 193225
rect 281722 193151 281778 193160
rect 281906 193216 281908 193225
rect 281960 193216 281962 193225
rect 281906 193151 281962 193160
rect 281920 186266 281948 193151
rect 281828 186238 281948 186266
rect 281828 178786 281856 186238
rect 281828 178758 281948 178786
rect 281920 173942 281948 178758
rect 281724 173936 281776 173942
rect 281722 173904 281724 173913
rect 281908 173936 281960 173942
rect 281776 173904 281778 173913
rect 281722 173839 281778 173848
rect 281906 173904 281908 173913
rect 281960 173904 281962 173913
rect 281906 173839 281962 173848
rect 281920 166818 281948 173839
rect 281828 166790 281948 166818
rect 281828 157434 281856 166790
rect 281736 157406 281856 157434
rect 281736 148374 281764 157406
rect 281724 148368 281776 148374
rect 281724 148310 281776 148316
rect 281724 143608 281776 143614
rect 281724 143550 281776 143556
rect 281736 125769 281764 143550
rect 281722 125760 281778 125769
rect 281722 125695 281778 125704
rect 281722 125624 281778 125633
rect 281722 125559 281778 125568
rect 281736 122074 281764 125559
rect 281736 122046 281948 122074
rect 281920 118538 281948 122046
rect 281828 118510 281948 118538
rect 281828 100586 281856 118510
rect 281736 100558 281856 100586
rect 281736 89010 281764 100558
rect 281724 89004 281776 89010
rect 281724 88946 281776 88952
rect 281816 75948 281868 75954
rect 281816 75890 281868 75896
rect 281828 67658 281856 75890
rect 281724 67652 281776 67658
rect 281724 67594 281776 67600
rect 281816 67652 281868 67658
rect 281816 67594 281868 67600
rect 281736 61470 281764 67594
rect 281724 61464 281776 61470
rect 281724 61406 281776 61412
rect 281724 48340 281776 48346
rect 281724 48282 281776 48288
rect 281736 38622 281764 48282
rect 281724 38616 281776 38622
rect 281724 38558 281776 38564
rect 281724 29028 281776 29034
rect 281724 28970 281776 28976
rect 281736 19446 281764 28970
rect 281724 19440 281776 19446
rect 281724 19382 281776 19388
rect 281632 19372 281684 19378
rect 281632 19314 281684 19320
rect 281644 11898 281672 19314
rect 281632 11892 281684 11898
rect 281632 11834 281684 11840
rect 281540 11824 281592 11830
rect 281540 11766 281592 11772
rect 283024 6662 283052 335582
rect 283116 7585 283144 340054
rect 283208 340054 283406 340082
rect 283576 340054 283866 340082
rect 284418 340054 284616 340082
rect 283102 7576 283158 7585
rect 283102 7511 283158 7520
rect 283012 6656 283064 6662
rect 283012 6598 283064 6604
rect 283208 5370 283236 340054
rect 283576 335646 283604 340054
rect 284300 336932 284352 336938
rect 284300 336874 284352 336880
rect 283564 335640 283616 335646
rect 283564 335582 283616 335588
rect 284312 5438 284340 336874
rect 284588 335220 284616 340054
rect 284864 336938 284892 340068
rect 285140 340054 285338 340082
rect 285798 340054 285904 340082
rect 284852 336932 284904 336938
rect 284852 336874 284904 336880
rect 284496 335192 284616 335220
rect 284496 8945 284524 335192
rect 285140 331242 285168 340054
rect 285588 337680 285640 337686
rect 285588 337622 285640 337628
rect 284772 331214 285168 331242
rect 284772 311982 284800 331214
rect 284760 311976 284812 311982
rect 284760 311918 284812 311924
rect 284760 311840 284812 311846
rect 284760 311782 284812 311788
rect 284772 299470 284800 311782
rect 284668 299464 284720 299470
rect 284668 299406 284720 299412
rect 284760 299464 284812 299470
rect 284760 299406 284812 299412
rect 284680 298110 284708 299406
rect 284668 298104 284720 298110
rect 284668 298046 284720 298052
rect 284760 298104 284812 298110
rect 284760 298046 284812 298052
rect 284772 280158 284800 298046
rect 284760 280152 284812 280158
rect 284760 280094 284812 280100
rect 284852 280152 284904 280158
rect 284852 280094 284904 280100
rect 284864 278769 284892 280094
rect 284666 278760 284722 278769
rect 284666 278695 284722 278704
rect 284850 278760 284906 278769
rect 284850 278695 284906 278704
rect 284680 269906 284708 278695
rect 284680 269878 284892 269906
rect 284864 259486 284892 269878
rect 284760 259480 284812 259486
rect 284760 259422 284812 259428
rect 284852 259480 284904 259486
rect 284852 259422 284904 259428
rect 284772 251190 284800 259422
rect 284668 251184 284720 251190
rect 284668 251126 284720 251132
rect 284760 251184 284812 251190
rect 284760 251126 284812 251132
rect 284680 248402 284708 251126
rect 284668 248396 284720 248402
rect 284668 248338 284720 248344
rect 284760 238808 284812 238814
rect 284760 238750 284812 238756
rect 284772 217410 284800 238750
rect 284772 217382 284892 217410
rect 284864 212566 284892 217382
rect 284668 212560 284720 212566
rect 284668 212502 284720 212508
rect 284852 212560 284904 212566
rect 284852 212502 284904 212508
rect 284680 205698 284708 212502
rect 284668 205692 284720 205698
rect 284668 205634 284720 205640
rect 284760 205556 284812 205562
rect 284760 205498 284812 205504
rect 284772 198098 284800 205498
rect 284772 198070 284892 198098
rect 284864 193254 284892 198070
rect 284668 193248 284720 193254
rect 284666 193216 284668 193225
rect 284852 193248 284904 193254
rect 284720 193216 284722 193225
rect 284666 193151 284722 193160
rect 284850 193216 284852 193225
rect 284904 193216 284906 193225
rect 284850 193151 284906 193160
rect 284864 186266 284892 193151
rect 284772 186238 284892 186266
rect 284772 178786 284800 186238
rect 284772 178758 284892 178786
rect 284864 173942 284892 178758
rect 284668 173936 284720 173942
rect 284666 173904 284668 173913
rect 284852 173936 284904 173942
rect 284720 173904 284722 173913
rect 284666 173839 284722 173848
rect 284850 173904 284852 173913
rect 284904 173904 284906 173913
rect 284850 173839 284906 173848
rect 284864 166818 284892 173839
rect 284772 166790 284892 166818
rect 284772 157434 284800 166790
rect 284680 157406 284800 157434
rect 284680 149682 284708 157406
rect 284588 149654 284708 149682
rect 284588 147370 284616 149654
rect 284588 147342 284800 147370
rect 284772 144906 284800 147342
rect 284668 144900 284720 144906
rect 284668 144842 284720 144848
rect 284760 144900 284812 144906
rect 284760 144842 284812 144848
rect 284680 139890 284708 144842
rect 284680 139862 284800 139890
rect 284772 125769 284800 139862
rect 284758 125760 284814 125769
rect 284758 125695 284814 125704
rect 284666 125624 284722 125633
rect 284666 125559 284722 125568
rect 284680 119490 284708 125559
rect 284680 119462 284892 119490
rect 284864 118674 284892 119462
rect 284772 118646 284892 118674
rect 284772 106282 284800 118646
rect 284760 106276 284812 106282
rect 284760 106218 284812 106224
rect 284852 106276 284904 106282
rect 284852 106218 284904 106224
rect 284864 96694 284892 106218
rect 284852 96688 284904 96694
rect 284852 96630 284904 96636
rect 284760 96620 284812 96626
rect 284760 96562 284812 96568
rect 284772 86970 284800 96562
rect 284576 86964 284628 86970
rect 284576 86906 284628 86912
rect 284760 86964 284812 86970
rect 284760 86906 284812 86912
rect 284588 72434 284616 86906
rect 284666 76120 284722 76129
rect 284722 76078 284800 76106
rect 284666 76055 284722 76064
rect 284772 75993 284800 76078
rect 284758 75984 284814 75993
rect 284758 75919 284814 75928
rect 284588 72406 284800 72434
rect 284772 58070 284800 72406
rect 284760 58064 284812 58070
rect 284760 58006 284812 58012
rect 284760 57928 284812 57934
rect 284760 57870 284812 57876
rect 284772 48346 284800 57870
rect 284668 48340 284720 48346
rect 284668 48282 284720 48288
rect 284760 48340 284812 48346
rect 284760 48282 284812 48288
rect 284680 46918 284708 48282
rect 284668 46912 284720 46918
rect 284668 46854 284720 46860
rect 284760 37324 284812 37330
rect 284760 37266 284812 37272
rect 284772 28966 284800 37266
rect 284576 28960 284628 28966
rect 284576 28902 284628 28908
rect 284760 28960 284812 28966
rect 284760 28902 284812 28908
rect 284588 19394 284616 28902
rect 284588 19366 284708 19394
rect 284680 12458 284708 19366
rect 284680 12430 284800 12458
rect 284772 12322 284800 12430
rect 284588 12294 284800 12322
rect 284482 8936 284538 8945
rect 284482 8871 284538 8880
rect 284588 7546 284616 12294
rect 284576 7540 284628 7546
rect 284576 7482 284628 7488
rect 284300 5432 284352 5438
rect 284300 5374 284352 5380
rect 283196 5364 283248 5370
rect 283196 5306 283248 5312
rect 283656 5296 283708 5302
rect 283656 5238 283708 5244
rect 282460 3936 282512 3942
rect 282460 3878 282512 3884
rect 281264 604 281316 610
rect 281264 546 281316 552
rect 281448 604 281500 610
rect 281448 546 281500 552
rect 281276 480 281304 546
rect 282472 480 282500 3878
rect 283668 480 283696 5238
rect 285600 4146 285628 337622
rect 285680 335640 285732 335646
rect 285680 335582 285732 335588
rect 285692 5506 285720 335582
rect 285770 325680 285826 325689
rect 285770 325615 285826 325624
rect 285784 316062 285812 325615
rect 285772 316056 285824 316062
rect 285772 315998 285824 316004
rect 285772 137760 285824 137766
rect 285772 137702 285824 137708
rect 285784 124273 285812 137702
rect 285770 124264 285826 124273
rect 285770 124199 285826 124208
rect 285876 9314 285904 340054
rect 285968 340054 286350 340082
rect 286612 340054 286810 340082
rect 287164 340054 287270 340082
rect 287348 340054 287822 340082
rect 287992 340054 288282 340082
rect 288544 340054 288742 340082
rect 289004 340054 289294 340082
rect 289464 340054 289754 340082
rect 289832 340054 290214 340082
rect 285968 335646 285996 340054
rect 285956 335640 286008 335646
rect 285956 335582 286008 335588
rect 286612 335510 286640 340054
rect 287060 335640 287112 335646
rect 287060 335582 287112 335588
rect 285956 335504 286008 335510
rect 285956 335446 286008 335452
rect 286600 335504 286652 335510
rect 286600 335446 286652 335452
rect 285968 325689 285996 335446
rect 285954 325680 286010 325689
rect 285954 325615 286010 325624
rect 286048 316056 286100 316062
rect 286046 316024 286048 316033
rect 286100 316024 286102 316033
rect 286046 315959 286102 315968
rect 286230 316024 286286 316033
rect 286230 315959 286286 315968
rect 286244 306406 286272 315959
rect 286140 306400 286192 306406
rect 286140 306342 286192 306348
rect 286232 306400 286284 306406
rect 286232 306342 286284 306348
rect 286152 298246 286180 306342
rect 286048 298240 286100 298246
rect 286048 298182 286100 298188
rect 286140 298240 286192 298246
rect 286140 298182 286192 298188
rect 286060 298110 286088 298182
rect 286048 298104 286100 298110
rect 286048 298046 286100 298052
rect 286140 298104 286192 298110
rect 286140 298046 286192 298052
rect 286152 275210 286180 298046
rect 286060 275182 286180 275210
rect 286060 270502 286088 275182
rect 286048 270496 286100 270502
rect 286048 270438 286100 270444
rect 286140 270496 286192 270502
rect 286140 270438 286192 270444
rect 286152 255950 286180 270438
rect 286140 255944 286192 255950
rect 286140 255886 286192 255892
rect 286048 247104 286100 247110
rect 286048 247046 286100 247052
rect 286060 238921 286088 247046
rect 286046 238912 286102 238921
rect 286046 238847 286102 238856
rect 285954 238776 286010 238785
rect 285954 238711 285956 238720
rect 286008 238711 286010 238720
rect 285956 238682 286008 238688
rect 286140 238604 286192 238610
rect 286140 238546 286192 238552
rect 286152 217274 286180 238546
rect 286060 217246 286180 217274
rect 286060 212498 286088 217246
rect 286048 212492 286100 212498
rect 286048 212434 286100 212440
rect 286140 202904 286192 202910
rect 286140 202846 286192 202852
rect 286152 197962 286180 202846
rect 286060 197934 286180 197962
rect 286060 191826 286088 197934
rect 285956 191820 286008 191826
rect 285956 191762 286008 191768
rect 286048 191820 286100 191826
rect 286048 191762 286100 191768
rect 285968 182209 285996 191762
rect 285954 182200 286010 182209
rect 285954 182135 286010 182144
rect 286138 182200 286194 182209
rect 286138 182135 286194 182144
rect 286152 173913 286180 182135
rect 285954 173904 286010 173913
rect 285954 173839 286010 173848
rect 286138 173904 286194 173913
rect 286138 173839 286194 173848
rect 285968 164286 285996 173839
rect 285956 164280 286008 164286
rect 285956 164222 286008 164228
rect 286140 164144 286192 164150
rect 286140 164086 286192 164092
rect 286152 161430 286180 164086
rect 286140 161424 286192 161430
rect 286140 161366 286192 161372
rect 285956 151836 286008 151842
rect 285956 151778 286008 151784
rect 285968 147778 285996 151778
rect 285968 147750 286088 147778
rect 286060 143562 286088 147750
rect 286060 143534 286180 143562
rect 286152 137766 286180 143534
rect 286140 137760 286192 137766
rect 286140 137702 286192 137708
rect 286966 134192 287022 134201
rect 286966 134127 287022 134136
rect 286980 133793 287008 134127
rect 286966 133784 287022 133793
rect 286966 133719 287022 133728
rect 285954 124264 286010 124273
rect 285954 124199 286010 124208
rect 285968 122806 285996 124199
rect 285956 122800 286008 122806
rect 285956 122742 286008 122748
rect 286048 122800 286100 122806
rect 286048 122742 286100 122748
rect 286060 113234 286088 122742
rect 285968 113206 286088 113234
rect 285968 113150 285996 113206
rect 285956 113144 286008 113150
rect 285956 113086 286008 113092
rect 286048 103556 286100 103562
rect 286048 103498 286100 103504
rect 286060 93786 286088 103498
rect 286060 93758 286180 93786
rect 286152 84998 286180 93758
rect 286230 87272 286286 87281
rect 286230 87207 286286 87216
rect 286244 87009 286272 87207
rect 286230 87000 286286 87009
rect 286230 86935 286286 86944
rect 286140 84992 286192 84998
rect 286140 84934 286192 84940
rect 286140 75948 286192 75954
rect 286140 75890 286192 75896
rect 286152 75834 286180 75890
rect 286152 75806 286272 75834
rect 286244 56681 286272 75806
rect 286046 56672 286102 56681
rect 286046 56607 286102 56616
rect 286230 56672 286286 56681
rect 286230 56607 286286 56616
rect 286060 46918 286088 56607
rect 286048 46912 286100 46918
rect 286048 46854 286100 46860
rect 286140 46912 286192 46918
rect 286140 46854 286192 46860
rect 286152 26058 286180 46854
rect 286060 26030 286180 26058
rect 286060 12322 286088 26030
rect 285968 12294 286088 12322
rect 285864 9308 285916 9314
rect 285864 9250 285916 9256
rect 285968 7478 285996 12294
rect 285956 7472 286008 7478
rect 285956 7414 286008 7420
rect 287072 7410 287100 335582
rect 287164 9382 287192 340054
rect 287348 11966 287376 340054
rect 287992 335646 288020 340054
rect 288256 337816 288308 337822
rect 288256 337758 288308 337764
rect 287980 335640 288032 335646
rect 287980 335582 288032 335588
rect 287336 11960 287388 11966
rect 287336 11902 287388 11908
rect 287152 9376 287204 9382
rect 287152 9318 287204 9324
rect 287060 7404 287112 7410
rect 287060 7346 287112 7352
rect 285680 5500 285732 5506
rect 285680 5442 285732 5448
rect 287152 5364 287204 5370
rect 287152 5306 287204 5312
rect 284760 4140 284812 4146
rect 284760 4082 284812 4088
rect 285588 4140 285640 4146
rect 285588 4082 285640 4088
rect 284772 480 284800 4082
rect 285956 3800 286008 3806
rect 285956 3742 286008 3748
rect 285968 480 285996 3742
rect 287164 480 287192 5306
rect 288268 626 288296 337758
rect 288440 335640 288492 335646
rect 288440 335582 288492 335588
rect 288346 16960 288402 16969
rect 288346 16895 288402 16904
rect 288360 16833 288388 16895
rect 288346 16824 288402 16833
rect 288346 16759 288402 16768
rect 288452 7342 288480 335582
rect 288544 10062 288572 340054
rect 289004 335345 289032 340054
rect 289464 335646 289492 340054
rect 289452 335640 289504 335646
rect 289452 335582 289504 335588
rect 288714 335336 288770 335345
rect 288714 335271 288770 335280
rect 288990 335336 289046 335345
rect 288990 335271 289046 335280
rect 288728 325718 288756 335271
rect 288716 325712 288768 325718
rect 288716 325654 288768 325660
rect 288808 325712 288860 325718
rect 288808 325654 288860 325660
rect 288820 307766 288848 325654
rect 288808 307760 288860 307766
rect 288808 307702 288860 307708
rect 288716 306400 288768 306406
rect 288714 306368 288716 306377
rect 288768 306368 288770 306377
rect 288714 306303 288770 306312
rect 288898 306368 288954 306377
rect 288898 306303 288954 306312
rect 288912 298178 288940 306303
rect 288900 298172 288952 298178
rect 288900 298114 288952 298120
rect 288900 298036 288952 298042
rect 288900 297978 288952 297984
rect 288912 289796 288940 297978
rect 288912 289768 289032 289796
rect 289004 289626 289032 289768
rect 288912 289598 289032 289626
rect 288912 288402 288940 289598
rect 288912 288374 289032 288402
rect 289004 284306 289032 288374
rect 288992 284300 289044 284306
rect 288992 284242 289044 284248
rect 288900 274712 288952 274718
rect 288900 274654 288952 274660
rect 288912 259146 288940 274654
rect 288900 259140 288952 259146
rect 288900 259082 288952 259088
rect 288808 241528 288860 241534
rect 288808 241470 288860 241476
rect 288820 230518 288848 241470
rect 288716 230512 288768 230518
rect 288716 230454 288768 230460
rect 288808 230512 288860 230518
rect 288808 230454 288860 230460
rect 288728 225010 288756 230454
rect 288716 225004 288768 225010
rect 288716 224946 288768 224952
rect 288808 224868 288860 224874
rect 288808 224810 288860 224816
rect 288820 220833 288848 224810
rect 288806 220824 288862 220833
rect 288806 220759 288862 220768
rect 288714 220688 288770 220697
rect 288714 220623 288770 220632
rect 288728 205698 288756 220623
rect 288716 205692 288768 205698
rect 288716 205634 288768 205640
rect 288808 205624 288860 205630
rect 288808 205566 288860 205572
rect 288820 198098 288848 205566
rect 288820 198070 288940 198098
rect 288912 193254 288940 198070
rect 288716 193248 288768 193254
rect 288714 193216 288716 193225
rect 288900 193248 288952 193254
rect 288768 193216 288770 193225
rect 288714 193151 288770 193160
rect 288898 193216 288900 193225
rect 288952 193216 288954 193225
rect 288898 193151 288954 193160
rect 288912 186266 288940 193151
rect 288820 186238 288940 186266
rect 288820 178786 288848 186238
rect 288820 178758 288940 178786
rect 288912 173942 288940 178758
rect 288716 173936 288768 173942
rect 288716 173878 288768 173884
rect 288900 173936 288952 173942
rect 288900 173878 288952 173884
rect 288728 169130 288756 173878
rect 288728 169102 288848 169130
rect 288820 156754 288848 169102
rect 288728 156726 288848 156754
rect 288728 129010 288756 156726
rect 288728 128982 288848 129010
rect 288820 122806 288848 128982
rect 288716 122800 288768 122806
rect 288716 122742 288768 122748
rect 288808 122800 288860 122806
rect 288808 122742 288860 122748
rect 288728 67946 288756 122742
rect 288636 67918 288756 67946
rect 288636 67674 288664 67918
rect 288636 67646 288756 67674
rect 288728 57050 288756 67646
rect 288716 57044 288768 57050
rect 288716 56986 288768 56992
rect 288716 48340 288768 48346
rect 288716 48282 288768 48288
rect 288728 42106 288756 48282
rect 288728 42078 288940 42106
rect 288912 38570 288940 42078
rect 288820 38542 288940 38570
rect 288820 37262 288848 38542
rect 288808 37256 288860 37262
rect 288808 37198 288860 37204
rect 288900 37256 288952 37262
rect 288900 37198 288952 37204
rect 288912 12034 288940 37198
rect 288900 12028 288952 12034
rect 288900 11970 288952 11976
rect 288532 10056 288584 10062
rect 288532 9998 288584 10004
rect 289832 9994 289860 340054
rect 290292 335594 290320 340190
rect 290464 336796 290516 336802
rect 290464 336738 290516 336744
rect 290108 335566 290320 335594
rect 290108 317422 290136 335566
rect 290096 317416 290148 317422
rect 290096 317358 290148 317364
rect 290188 317416 290240 317422
rect 290188 317358 290240 317364
rect 290200 294642 290228 317358
rect 290004 294636 290056 294642
rect 290004 294578 290056 294584
rect 290188 294636 290240 294642
rect 290188 294578 290240 294584
rect 290016 289814 290044 294578
rect 290004 289808 290056 289814
rect 290004 289750 290056 289756
rect 290188 289808 290240 289814
rect 290188 289750 290240 289756
rect 290200 269142 290228 289750
rect 290096 269136 290148 269142
rect 290096 269078 290148 269084
rect 290188 269136 290240 269142
rect 290188 269078 290240 269084
rect 290108 251258 290136 269078
rect 290004 251252 290056 251258
rect 290004 251194 290056 251200
rect 290096 251252 290148 251258
rect 290096 251194 290148 251200
rect 290016 241534 290044 251194
rect 290004 241528 290056 241534
rect 290004 241470 290056 241476
rect 290188 241528 290240 241534
rect 290188 241470 290240 241476
rect 290200 235362 290228 241470
rect 290200 235334 290412 235362
rect 290384 220930 290412 235334
rect 290372 220924 290424 220930
rect 290372 220866 290424 220872
rect 290188 220856 290240 220862
rect 290186 220824 290188 220833
rect 290240 220824 290242 220833
rect 290186 220759 290242 220768
rect 290186 220688 290242 220697
rect 290186 220623 290242 220632
rect 290200 219434 290228 220623
rect 290188 219428 290240 219434
rect 290188 219370 290240 219376
rect 290188 211132 290240 211138
rect 290188 211074 290240 211080
rect 290200 209794 290228 211074
rect 290200 209766 290320 209794
rect 290292 204218 290320 209766
rect 290200 204190 290320 204218
rect 290200 200122 290228 204190
rect 290188 200116 290240 200122
rect 290188 200058 290240 200064
rect 290004 190528 290056 190534
rect 290004 190470 290056 190476
rect 290016 188358 290044 190470
rect 290004 188352 290056 188358
rect 290004 188294 290056 188300
rect 290004 188216 290056 188222
rect 290004 188158 290056 188164
rect 290016 182170 290044 188158
rect 290004 182164 290056 182170
rect 290004 182106 290056 182112
rect 290004 172576 290056 172582
rect 290004 172518 290056 172524
rect 290016 153202 290044 172518
rect 290004 153196 290056 153202
rect 290004 153138 290056 153144
rect 290096 153196 290148 153202
rect 290096 153138 290148 153144
rect 290108 132530 290136 153138
rect 289912 132524 289964 132530
rect 289912 132466 289964 132472
rect 290096 132524 290148 132530
rect 290096 132466 290148 132472
rect 289924 124234 289952 132466
rect 289912 124228 289964 124234
rect 289912 124170 289964 124176
rect 290004 124228 290056 124234
rect 290004 124170 290056 124176
rect 290016 119898 290044 124170
rect 289924 119870 290044 119898
rect 289924 114458 289952 119870
rect 289924 114430 290136 114458
rect 290108 111790 290136 114430
rect 290096 111784 290148 111790
rect 290096 111726 290148 111732
rect 290004 104236 290056 104242
rect 290004 104178 290056 104184
rect 290016 97986 290044 104178
rect 290004 97980 290056 97986
rect 290004 97922 290056 97928
rect 290004 93832 290056 93838
rect 290004 93774 290056 93780
rect 290016 88346 290044 93774
rect 290016 88318 290136 88346
rect 290108 84250 290136 88318
rect 290096 84244 290148 84250
rect 290096 84186 290148 84192
rect 290188 84108 290240 84114
rect 290188 84050 290240 84056
rect 290200 60761 290228 84050
rect 290002 60752 290058 60761
rect 290002 60687 290058 60696
rect 290186 60752 290242 60761
rect 290186 60687 290242 60696
rect 290016 12102 290044 60687
rect 290004 12096 290056 12102
rect 290004 12038 290056 12044
rect 289820 9988 289872 9994
rect 289820 9930 289872 9936
rect 288440 7336 288492 7342
rect 288440 7278 288492 7284
rect 289820 6520 289872 6526
rect 289820 6462 289872 6468
rect 288440 6452 288492 6458
rect 288440 6394 288492 6400
rect 288452 3330 288480 6394
rect 288532 6384 288584 6390
rect 288532 6326 288584 6332
rect 288440 3324 288492 3330
rect 288440 3266 288492 3272
rect 288544 3262 288572 6326
rect 289544 3868 289596 3874
rect 289544 3810 289596 3816
rect 288532 3256 288584 3262
rect 288532 3198 288584 3204
rect 288268 598 288388 626
rect 288360 480 288388 598
rect 289556 480 289584 3810
rect 289832 3398 289860 6462
rect 289820 3392 289872 3398
rect 289820 3334 289872 3340
rect 290476 3194 290504 336738
rect 291212 7274 291240 340068
rect 291304 340054 291686 340082
rect 291304 9926 291332 340054
rect 291764 335594 291792 340190
rect 291580 335566 291792 335594
rect 292592 340054 292698 340082
rect 292868 340054 293158 340082
rect 293328 340054 293710 340082
rect 293972 340054 294170 340082
rect 294248 340054 294630 340082
rect 291580 319410 291608 335566
rect 291488 319382 291608 319410
rect 291488 319138 291516 319382
rect 291488 319110 291608 319138
rect 291580 317422 291608 319110
rect 291568 317416 291620 317422
rect 291568 317358 291620 317364
rect 291660 317416 291712 317422
rect 291660 317358 291712 317364
rect 291672 306377 291700 317358
rect 291658 306368 291714 306377
rect 291658 306303 291714 306312
rect 291842 306368 291898 306377
rect 291842 306303 291898 306312
rect 291856 304978 291884 306303
rect 291752 304972 291804 304978
rect 291752 304914 291804 304920
rect 291844 304972 291896 304978
rect 291844 304914 291896 304920
rect 291764 303618 291792 304914
rect 291752 303612 291804 303618
rect 291752 303554 291804 303560
rect 291568 296540 291620 296546
rect 291568 296482 291620 296488
rect 291580 292534 291608 296482
rect 291568 292528 291620 292534
rect 291568 292470 291620 292476
rect 291384 274712 291436 274718
rect 291384 274654 291436 274660
rect 291396 258097 291424 274654
rect 291382 258088 291438 258097
rect 291566 258088 291622 258097
rect 291382 258023 291438 258032
rect 291476 258052 291528 258058
rect 291566 258023 291568 258032
rect 291476 257994 291528 258000
rect 291620 258023 291622 258032
rect 291568 257994 291620 258000
rect 291488 241534 291516 257994
rect 291476 241528 291528 241534
rect 291476 241470 291528 241476
rect 291660 241528 291712 241534
rect 291660 241470 291712 241476
rect 291672 235362 291700 241470
rect 291672 235334 291884 235362
rect 291856 220998 291884 235334
rect 291844 220992 291896 220998
rect 291844 220934 291896 220940
rect 291660 220856 291712 220862
rect 291660 220798 291712 220804
rect 291672 219434 291700 220798
rect 291660 219428 291712 219434
rect 291660 219370 291712 219376
rect 291660 204332 291712 204338
rect 291660 204274 291712 204280
rect 291672 193202 291700 204274
rect 291580 193174 291700 193202
rect 291580 183598 291608 193174
rect 291568 183592 291620 183598
rect 291568 183534 291620 183540
rect 291660 183592 291712 183598
rect 291660 183534 291712 183540
rect 291672 182170 291700 183534
rect 291660 182164 291712 182170
rect 291660 182106 291712 182112
rect 291660 173732 291712 173738
rect 291660 173674 291712 173680
rect 291672 164257 291700 173674
rect 291474 164248 291530 164257
rect 291474 164183 291530 164192
rect 291658 164248 291714 164257
rect 291658 164183 291714 164192
rect 291488 153202 291516 164183
rect 291476 153196 291528 153202
rect 291476 153138 291528 153144
rect 291568 153196 291620 153202
rect 291568 153138 291620 153144
rect 291580 129946 291608 153138
rect 291842 134056 291898 134065
rect 291842 133991 291898 134000
rect 291856 133793 291884 133991
rect 291842 133784 291898 133793
rect 291842 133719 291898 133728
rect 291568 129940 291620 129946
rect 291568 129882 291620 129888
rect 291476 129668 291528 129674
rect 291476 129610 291528 129616
rect 291488 120086 291516 129610
rect 291476 120080 291528 120086
rect 291476 120022 291528 120028
rect 291476 110492 291528 110498
rect 291476 110434 291528 110440
rect 291488 103562 291516 110434
rect 291476 103556 291528 103562
rect 291476 103498 291528 103504
rect 291660 103488 291712 103494
rect 291660 103430 291712 103436
rect 291672 85610 291700 103430
rect 291568 85604 291620 85610
rect 291568 85546 291620 85552
rect 291660 85604 291712 85610
rect 291660 85546 291712 85552
rect 291580 74594 291608 85546
rect 291384 74588 291436 74594
rect 291384 74530 291436 74536
rect 291568 74588 291620 74594
rect 291568 74530 291620 74536
rect 291396 67658 291424 74530
rect 291384 67652 291436 67658
rect 291384 67594 291436 67600
rect 291476 67652 291528 67658
rect 291476 67594 291528 67600
rect 291488 58070 291516 67594
rect 291476 58064 291528 58070
rect 291476 58006 291528 58012
rect 291384 57928 291436 57934
rect 291384 57870 291436 57876
rect 291396 48346 291424 57870
rect 291384 48340 291436 48346
rect 291384 48282 291436 48288
rect 291476 48340 291528 48346
rect 291476 48282 291528 48288
rect 291488 46918 291516 48282
rect 291476 46912 291528 46918
rect 291476 46854 291528 46860
rect 291568 35964 291620 35970
rect 291568 35906 291620 35912
rect 291580 27674 291608 35906
rect 291568 27668 291620 27674
rect 291568 27610 291620 27616
rect 291660 27668 291712 27674
rect 291660 27610 291712 27616
rect 291672 26246 291700 27610
rect 291660 26240 291712 26246
rect 291660 26182 291712 26188
rect 291568 16652 291620 16658
rect 291568 16594 291620 16600
rect 291580 12170 291608 16594
rect 291568 12164 291620 12170
rect 291568 12106 291620 12112
rect 291292 9920 291344 9926
rect 291292 9862 291344 9868
rect 291200 7268 291252 7274
rect 291200 7210 291252 7216
rect 292592 7206 292620 340054
rect 292764 335640 292816 335646
rect 292764 335582 292816 335588
rect 292776 13258 292804 335582
rect 292764 13252 292816 13258
rect 292764 13194 292816 13200
rect 292868 9858 292896 340054
rect 293328 335646 293356 340054
rect 293316 335640 293368 335646
rect 293316 335582 293368 335588
rect 292856 9852 292908 9858
rect 292856 9794 292908 9800
rect 292580 7200 292632 7206
rect 292580 7142 292632 7148
rect 293972 7138 294000 340054
rect 294248 335696 294276 340054
rect 294064 335668 294276 335696
rect 294064 9790 294092 335668
rect 294708 335594 294736 340190
rect 294248 335566 294736 335594
rect 295352 340054 295642 340082
rect 295720 340054 296102 340082
rect 296272 340054 296654 340082
rect 296732 340054 297114 340082
rect 297284 340054 297574 340082
rect 298126 340054 298232 340082
rect 294248 328438 294276 335566
rect 294236 328432 294288 328438
rect 294236 328374 294288 328380
rect 294420 328432 294472 328438
rect 294420 328374 294472 328380
rect 294432 323490 294460 328374
rect 294340 323462 294460 323490
rect 294340 312610 294368 323462
rect 294340 312582 294460 312610
rect 294432 304298 294460 312582
rect 294236 304292 294288 304298
rect 294236 304234 294288 304240
rect 294420 304292 294472 304298
rect 294420 304234 294472 304240
rect 294248 293298 294276 304234
rect 294248 293270 294460 293298
rect 294432 289796 294460 293270
rect 294340 289768 294460 289796
rect 294340 280226 294368 289768
rect 294236 280220 294288 280226
rect 294236 280162 294288 280168
rect 294328 280220 294380 280226
rect 294328 280162 294380 280168
rect 294248 276010 294276 280162
rect 294236 276004 294288 276010
rect 294236 275946 294288 275952
rect 294328 276004 294380 276010
rect 294328 275946 294380 275952
rect 294340 266354 294368 275946
rect 294328 266348 294380 266354
rect 294328 266290 294380 266296
rect 294420 266348 294472 266354
rect 294420 266290 294472 266296
rect 294432 251870 294460 266290
rect 294420 251864 294472 251870
rect 294420 251806 294472 251812
rect 294420 238808 294472 238814
rect 294420 238750 294472 238756
rect 294432 222222 294460 238750
rect 294328 222216 294380 222222
rect 294328 222158 294380 222164
rect 294420 222216 294472 222222
rect 294420 222158 294472 222164
rect 294248 202910 294276 202941
rect 294340 202910 294368 222158
rect 294236 202904 294288 202910
rect 294328 202904 294380 202910
rect 294288 202852 294328 202858
rect 294236 202846 294380 202852
rect 294248 202830 294368 202846
rect 294340 188442 294368 202830
rect 294248 188414 294368 188442
rect 294248 178770 294276 188414
rect 294236 178764 294288 178770
rect 294236 178706 294288 178712
rect 294420 178764 294472 178770
rect 294420 178706 294472 178712
rect 294432 161498 294460 178706
rect 294328 161492 294380 161498
rect 294328 161434 294380 161440
rect 294420 161492 294472 161498
rect 294420 161434 294472 161440
rect 294340 153202 294368 161434
rect 294236 153196 294288 153202
rect 294236 153138 294288 153144
rect 294328 153196 294380 153202
rect 294328 153138 294380 153144
rect 294248 137306 294276 153138
rect 294248 137278 294460 137306
rect 294432 122806 294460 137278
rect 294420 122800 294472 122806
rect 294420 122742 294472 122748
rect 294420 113212 294472 113218
rect 294420 113154 294472 113160
rect 294432 103562 294460 113154
rect 294420 103556 294472 103562
rect 294420 103498 294472 103504
rect 294604 103488 294656 103494
rect 294604 103430 294656 103436
rect 294616 85610 294644 103430
rect 294420 85604 294472 85610
rect 294420 85546 294472 85552
rect 294604 85604 294656 85610
rect 294604 85546 294656 85552
rect 294432 74526 294460 85546
rect 294420 74520 294472 74526
rect 294420 74462 294472 74468
rect 294236 64932 294288 64938
rect 294236 64874 294288 64880
rect 294248 45529 294276 64874
rect 294234 45520 294290 45529
rect 294234 45455 294290 45464
rect 294142 36000 294198 36009
rect 294142 35935 294198 35944
rect 294156 35902 294184 35935
rect 294144 35896 294196 35902
rect 294144 35838 294196 35844
rect 294512 35896 294564 35902
rect 294512 35838 294564 35844
rect 294524 19292 294552 35838
rect 294432 19264 294552 19292
rect 294432 13326 294460 19264
rect 294420 13320 294472 13326
rect 294420 13262 294472 13268
rect 294052 9784 294104 9790
rect 294052 9726 294104 9732
rect 293960 7132 294012 7138
rect 293960 7074 294012 7080
rect 295352 7070 295380 340054
rect 295720 335696 295748 340054
rect 295444 335668 295748 335696
rect 295444 9722 295472 335668
rect 296272 335594 296300 340054
rect 295536 335566 296300 335594
rect 295536 328438 295564 335566
rect 295524 328432 295576 328438
rect 295524 328374 295576 328380
rect 295708 328432 295760 328438
rect 295708 328374 295760 328380
rect 295720 323490 295748 328374
rect 295628 323462 295748 323490
rect 295628 312610 295656 323462
rect 295628 312582 295748 312610
rect 295720 304298 295748 312582
rect 295524 304292 295576 304298
rect 295524 304234 295576 304240
rect 295708 304292 295760 304298
rect 295708 304234 295760 304240
rect 295536 292602 295564 304234
rect 295524 292596 295576 292602
rect 295524 292538 295576 292544
rect 295616 292528 295668 292534
rect 295616 292470 295668 292476
rect 295628 283014 295656 292470
rect 295616 283008 295668 283014
rect 295616 282950 295668 282956
rect 295524 282872 295576 282878
rect 295524 282814 295576 282820
rect 295536 269142 295564 282814
rect 295524 269136 295576 269142
rect 295524 269078 295576 269084
rect 295800 269136 295852 269142
rect 295800 269078 295852 269084
rect 295812 260930 295840 269078
rect 295812 260902 295932 260930
rect 295904 258097 295932 260902
rect 295706 258088 295762 258097
rect 295524 258052 295576 258058
rect 295706 258023 295708 258032
rect 295524 257994 295576 258000
rect 295760 258023 295762 258032
rect 295890 258088 295946 258097
rect 295890 258023 295946 258032
rect 295708 257994 295760 258000
rect 295536 241482 295564 257994
rect 295536 241454 295656 241482
rect 295536 222222 295564 222253
rect 295628 222222 295656 241454
rect 295524 222216 295576 222222
rect 295616 222216 295668 222222
rect 295576 222164 295616 222170
rect 295524 222158 295668 222164
rect 295536 222142 295656 222158
rect 295536 202910 295564 202941
rect 295628 202910 295656 222142
rect 295524 202904 295576 202910
rect 295616 202904 295668 202910
rect 295576 202852 295616 202858
rect 295524 202846 295668 202852
rect 295536 202830 295656 202846
rect 295628 186386 295656 202830
rect 295616 186380 295668 186386
rect 295616 186322 295668 186328
rect 295524 186312 295576 186318
rect 295524 186254 295576 186260
rect 295536 178770 295564 186254
rect 295524 178764 295576 178770
rect 295524 178706 295576 178712
rect 295708 178764 295760 178770
rect 295708 178706 295760 178712
rect 295720 161498 295748 178706
rect 295616 161492 295668 161498
rect 295616 161434 295668 161440
rect 295708 161492 295760 161498
rect 295708 161434 295760 161440
rect 295628 143562 295656 161434
rect 296628 150408 296680 150414
rect 296628 150350 296680 150356
rect 295536 143534 295656 143562
rect 295536 132530 295564 143534
rect 296640 140865 296668 150350
rect 296626 140856 296682 140865
rect 296626 140791 296682 140800
rect 295524 132524 295576 132530
rect 295524 132466 295576 132472
rect 295616 132524 295668 132530
rect 295616 132466 295668 132472
rect 295628 132410 295656 132466
rect 295536 132382 295656 132410
rect 295536 124114 295564 132382
rect 295536 124086 295748 124114
rect 295720 122806 295748 124086
rect 296534 123312 296590 123321
rect 296534 123247 296590 123256
rect 296548 123049 296576 123247
rect 296534 123040 296590 123049
rect 296534 122975 296590 122984
rect 295708 122800 295760 122806
rect 295708 122742 295760 122748
rect 295800 116612 295852 116618
rect 295800 116554 295852 116560
rect 295812 111874 295840 116554
rect 295720 111846 295840 111874
rect 295720 111790 295748 111846
rect 295708 111784 295760 111790
rect 295708 111726 295760 111732
rect 295892 102196 295944 102202
rect 295892 102138 295944 102144
rect 295904 82890 295932 102138
rect 295708 82884 295760 82890
rect 295708 82826 295760 82832
rect 295892 82884 295944 82890
rect 295892 82826 295944 82832
rect 295720 64938 295748 82826
rect 295616 64932 295668 64938
rect 295616 64874 295668 64880
rect 295708 64932 295760 64938
rect 295708 64874 295760 64880
rect 295628 61470 295656 64874
rect 295616 61464 295668 61470
rect 295616 61406 295668 61412
rect 295524 48340 295576 48346
rect 295524 48282 295576 48288
rect 295536 38434 295564 48282
rect 295536 38406 295656 38434
rect 295628 27742 295656 38406
rect 295616 27736 295668 27742
rect 295616 27678 295668 27684
rect 295524 27668 295576 27674
rect 295524 27610 295576 27616
rect 295536 19310 295564 27610
rect 295524 19304 295576 19310
rect 295524 19246 295576 19252
rect 295432 9716 295484 9722
rect 295432 9658 295484 9664
rect 295340 7064 295392 7070
rect 295340 7006 295392 7012
rect 296732 6730 296760 340054
rect 297284 332194 297312 340054
rect 297916 337476 297968 337482
rect 297916 337418 297968 337424
rect 296824 332166 297312 332194
rect 296824 328438 296852 332166
rect 296812 328432 296864 328438
rect 296812 328374 296864 328380
rect 296996 328432 297048 328438
rect 296996 328374 297048 328380
rect 297008 323490 297036 328374
rect 296916 323462 297036 323490
rect 296916 317422 296944 323462
rect 296904 317416 296956 317422
rect 296904 317358 296956 317364
rect 296996 317416 297048 317422
rect 296996 317358 297048 317364
rect 297008 301170 297036 317358
rect 296812 301164 296864 301170
rect 296812 301106 296864 301112
rect 296996 301164 297048 301170
rect 296996 301106 297048 301112
rect 296824 289626 296852 301106
rect 296824 289598 297036 289626
rect 297008 287042 297036 289598
rect 296916 287014 297036 287042
rect 296916 277438 296944 287014
rect 296812 277432 296864 277438
rect 296810 277400 296812 277409
rect 296904 277432 296956 277438
rect 296864 277400 296866 277409
rect 296904 277374 296956 277380
rect 297086 277400 297142 277409
rect 296810 277335 296866 277344
rect 297086 277335 297142 277344
rect 297100 276010 297128 277335
rect 297088 276004 297140 276010
rect 297088 275946 297140 275952
rect 296996 266416 297048 266422
rect 296996 266358 297048 266364
rect 297008 262954 297036 266358
rect 296812 262948 296864 262954
rect 296812 262890 296864 262896
rect 296996 262948 297048 262954
rect 296996 262890 297048 262896
rect 296824 258097 296852 262890
rect 296810 258088 296866 258097
rect 296810 258023 296866 258032
rect 296994 258088 297050 258097
rect 296994 258023 297050 258032
rect 297008 257990 297036 258023
rect 296996 257984 297048 257990
rect 296996 257926 297048 257932
rect 296812 249484 296864 249490
rect 296812 249426 296864 249432
rect 296824 241482 296852 249426
rect 296824 241454 296944 241482
rect 296824 222222 296852 222253
rect 296916 222222 296944 241454
rect 296812 222216 296864 222222
rect 296904 222216 296956 222222
rect 296864 222164 296904 222170
rect 296812 222158 296956 222164
rect 296824 222142 296944 222158
rect 296824 202910 296852 202941
rect 296916 202910 296944 222142
rect 296812 202904 296864 202910
rect 296904 202904 296956 202910
rect 296864 202852 296904 202858
rect 296812 202846 296956 202852
rect 296824 202830 296944 202846
rect 296916 186454 296944 202830
rect 296904 186448 296956 186454
rect 296904 186390 296956 186396
rect 296812 186312 296864 186318
rect 296812 186254 296864 186260
rect 296824 178770 296852 186254
rect 296812 178764 296864 178770
rect 296812 178706 296864 178712
rect 296996 178764 297048 178770
rect 296996 178706 297048 178712
rect 297008 161498 297036 178706
rect 296904 161492 296956 161498
rect 296904 161434 296956 161440
rect 296996 161492 297048 161498
rect 296996 161434 297048 161440
rect 296916 150414 296944 161434
rect 296904 150408 296956 150414
rect 296904 150350 296956 150356
rect 296810 140856 296866 140865
rect 296810 140791 296866 140800
rect 296824 140758 296852 140791
rect 296812 140752 296864 140758
rect 296812 140694 296864 140700
rect 296996 140752 297048 140758
rect 296996 140694 297048 140700
rect 297008 139398 297036 140694
rect 296996 139392 297048 139398
rect 296996 139334 297048 139340
rect 296996 122732 297048 122738
rect 296996 122674 297048 122680
rect 297008 112878 297036 122674
rect 296996 112872 297048 112878
rect 296996 112814 297048 112820
rect 296996 112736 297048 112742
rect 296996 112678 297048 112684
rect 297008 103562 297036 112678
rect 296904 103556 296956 103562
rect 296904 103498 296956 103504
rect 296996 103556 297048 103562
rect 296996 103498 297048 103504
rect 296916 95198 296944 103498
rect 296904 95192 296956 95198
rect 296904 95134 296956 95140
rect 296996 95192 297048 95198
rect 296996 95134 297048 95140
rect 297008 77382 297036 95134
rect 296996 77376 297048 77382
rect 296996 77318 297048 77324
rect 296812 77240 296864 77246
rect 296812 77182 296864 77188
rect 296824 46866 296852 77182
rect 296824 46838 296944 46866
rect 296916 13394 296944 46838
rect 296904 13388 296956 13394
rect 296904 13330 296956 13336
rect 296720 6724 296772 6730
rect 296720 6666 296772 6672
rect 297364 6724 297416 6730
rect 297364 6666 297416 6672
rect 295892 6656 295944 6662
rect 295892 6598 295944 6604
rect 294328 6316 294380 6322
rect 294328 6258 294380 6264
rect 290740 5432 290792 5438
rect 290740 5374 290792 5380
rect 290464 3188 290516 3194
rect 290464 3130 290516 3136
rect 290752 480 290780 5374
rect 291936 3256 291988 3262
rect 291936 3198 291988 3204
rect 291948 480 291976 3198
rect 293132 3052 293184 3058
rect 293132 2994 293184 3000
rect 293144 480 293172 2994
rect 294340 480 294368 6258
rect 295904 4146 295932 6598
rect 295892 4140 295944 4146
rect 295892 4082 295944 4088
rect 296720 4140 296772 4146
rect 296720 4082 296772 4088
rect 295524 3120 295576 3126
rect 295524 3062 295576 3068
rect 295536 480 295564 3062
rect 296732 480 296760 4082
rect 297376 4010 297404 6666
rect 297824 5500 297876 5506
rect 297824 5442 297876 5448
rect 297836 4026 297864 5442
rect 297928 4146 297956 337418
rect 298204 12306 298232 340054
rect 298388 340054 298586 340082
rect 298664 340054 299046 340082
rect 298284 335640 298336 335646
rect 298284 335582 298336 335588
rect 298296 13462 298324 335582
rect 298284 13456 298336 13462
rect 298284 13398 298336 13404
rect 298192 12300 298244 12306
rect 298192 12242 298244 12248
rect 298388 6798 298416 340054
rect 298664 335646 298692 340054
rect 298652 335640 298704 335646
rect 298652 335582 298704 335588
rect 299584 331294 299612 340068
rect 299768 340054 300058 340082
rect 300412 340054 300518 340082
rect 300964 340054 301070 340082
rect 301240 340054 301530 340082
rect 301700 340054 301990 340082
rect 302344 340054 302542 340082
rect 302712 340054 303002 340082
rect 303080 340054 303462 340082
rect 303724 340054 303922 340082
rect 304184 340054 304474 340082
rect 304644 340054 304934 340082
rect 305104 340054 305394 340082
rect 305656 340054 305946 340082
rect 299572 331288 299624 331294
rect 299768 331242 299796 340054
rect 300412 339130 300440 340054
rect 299572 331230 299624 331236
rect 299676 331214 299796 331242
rect 300320 339102 300440 339130
rect 299572 331152 299624 331158
rect 299572 331094 299624 331100
rect 299480 331084 299532 331090
rect 299480 331026 299532 331032
rect 299492 241466 299520 331026
rect 299480 241460 299532 241466
rect 299480 241402 299532 241408
rect 299480 231872 299532 231878
rect 299480 231814 299532 231820
rect 299388 16992 299440 16998
rect 299388 16934 299440 16940
rect 299400 16833 299428 16934
rect 299386 16824 299442 16833
rect 299386 16759 299442 16768
rect 299492 6866 299520 231814
rect 299584 12374 299612 331094
rect 299676 331090 299704 331214
rect 300320 331158 300348 339102
rect 300860 335640 300912 335646
rect 300860 335582 300912 335588
rect 299756 331152 299808 331158
rect 299756 331094 299808 331100
rect 300308 331152 300360 331158
rect 300308 331094 300360 331100
rect 299664 331084 299716 331090
rect 299664 331026 299716 331032
rect 299768 318850 299796 331094
rect 299756 318844 299808 318850
rect 299756 318786 299808 318792
rect 299848 318844 299900 318850
rect 299848 318786 299900 318792
rect 299860 311982 299888 318786
rect 299848 311976 299900 311982
rect 299848 311918 299900 311924
rect 299756 311840 299808 311846
rect 299756 311782 299808 311788
rect 299768 299538 299796 311782
rect 299756 299532 299808 299538
rect 299756 299474 299808 299480
rect 299848 299532 299900 299538
rect 299848 299474 299900 299480
rect 299860 292670 299888 299474
rect 299848 292664 299900 292670
rect 299848 292606 299900 292612
rect 299848 292528 299900 292534
rect 299848 292470 299900 292476
rect 299860 270638 299888 292470
rect 299848 270632 299900 270638
rect 299848 270574 299900 270580
rect 299756 270564 299808 270570
rect 299756 270506 299808 270512
rect 299768 266914 299796 270506
rect 299768 266886 299980 266914
rect 299952 263514 299980 266886
rect 299860 263486 299980 263514
rect 299860 254674 299888 263486
rect 299860 254646 299980 254674
rect 299952 249830 299980 254646
rect 299756 249824 299808 249830
rect 299756 249766 299808 249772
rect 299940 249824 299992 249830
rect 299940 249766 299992 249772
rect 299768 240174 299796 249766
rect 299756 240168 299808 240174
rect 299756 240110 299808 240116
rect 299940 240168 299992 240174
rect 299940 240110 299992 240116
rect 299952 231962 299980 240110
rect 299952 231934 300072 231962
rect 300044 231690 300072 231934
rect 299860 231662 300072 231690
rect 299860 220810 299888 231662
rect 299860 220782 299980 220810
rect 299952 213722 299980 220782
rect 299756 213716 299808 213722
rect 299756 213658 299808 213664
rect 299940 213716 299992 213722
rect 299940 213658 299992 213664
rect 299768 202910 299796 213658
rect 299756 202904 299808 202910
rect 299756 202846 299808 202852
rect 299848 202904 299900 202910
rect 299848 202846 299900 202852
rect 299860 196110 299888 202846
rect 299848 196104 299900 196110
rect 299848 196046 299900 196052
rect 299756 195968 299808 195974
rect 299756 195910 299808 195916
rect 299768 183598 299796 195910
rect 299756 183592 299808 183598
rect 299756 183534 299808 183540
rect 299848 183592 299900 183598
rect 299848 183534 299900 183540
rect 299860 176798 299888 183534
rect 299848 176792 299900 176798
rect 299848 176734 299900 176740
rect 299756 171148 299808 171154
rect 299756 171090 299808 171096
rect 299768 156670 299796 171090
rect 299756 156664 299808 156670
rect 299756 156606 299808 156612
rect 299940 156664 299992 156670
rect 299940 156606 299992 156612
rect 299952 137426 299980 156606
rect 299756 137420 299808 137426
rect 299756 137362 299808 137368
rect 299940 137420 299992 137426
rect 299940 137362 299992 137368
rect 299768 133890 299796 137362
rect 299756 133884 299808 133890
rect 299756 133826 299808 133832
rect 299848 124228 299900 124234
rect 299848 124170 299900 124176
rect 299860 115954 299888 124170
rect 299676 115926 299888 115954
rect 299676 104922 299704 115926
rect 299664 104916 299716 104922
rect 299664 104858 299716 104864
rect 299756 104916 299808 104922
rect 299756 104858 299808 104864
rect 299768 95334 299796 104858
rect 299756 95328 299808 95334
rect 299756 95270 299808 95276
rect 299848 95260 299900 95266
rect 299848 95202 299900 95208
rect 299860 77382 299888 95202
rect 299848 77376 299900 77382
rect 299848 77318 299900 77324
rect 299848 77240 299900 77246
rect 299848 77182 299900 77188
rect 299860 67658 299888 77182
rect 299756 67652 299808 67658
rect 299756 67594 299808 67600
rect 299848 67652 299900 67658
rect 299848 67594 299900 67600
rect 299768 48346 299796 67594
rect 299756 48340 299808 48346
rect 299756 48282 299808 48288
rect 299848 48204 299900 48210
rect 299848 48146 299900 48152
rect 299860 45558 299888 48146
rect 299848 45552 299900 45558
rect 299848 45494 299900 45500
rect 299756 35964 299808 35970
rect 299756 35906 299808 35912
rect 299768 29050 299796 35906
rect 299676 29022 299796 29050
rect 299676 28914 299704 29022
rect 299676 28886 299796 28914
rect 299768 13530 299796 28886
rect 299756 13524 299808 13530
rect 299756 13466 299808 13472
rect 299572 12368 299624 12374
rect 299572 12310 299624 12316
rect 299480 6860 299532 6866
rect 299480 6802 299532 6808
rect 298376 6792 298428 6798
rect 298376 6734 298428 6740
rect 298100 6588 298152 6594
rect 298100 6530 298152 6536
rect 297916 4140 297968 4146
rect 297916 4082 297968 4088
rect 298112 4078 298140 6530
rect 300872 6118 300900 335582
rect 300964 12442 300992 340054
rect 301240 335646 301268 340054
rect 301228 335640 301280 335646
rect 301228 335582 301280 335588
rect 301700 328506 301728 340054
rect 302240 335708 302292 335714
rect 302240 335650 302292 335656
rect 301136 328500 301188 328506
rect 301136 328442 301188 328448
rect 301688 328500 301740 328506
rect 301688 328442 301740 328448
rect 301148 327078 301176 328442
rect 301136 327072 301188 327078
rect 301136 327014 301188 327020
rect 301044 317484 301096 317490
rect 301044 317426 301096 317432
rect 301056 307986 301084 317426
rect 301056 307958 301176 307986
rect 301148 307850 301176 307958
rect 301056 307822 301176 307850
rect 301056 298110 301084 307822
rect 301044 298104 301096 298110
rect 301044 298046 301096 298052
rect 301044 292528 301096 292534
rect 301044 292470 301096 292476
rect 301056 273290 301084 292470
rect 301044 273284 301096 273290
rect 301044 273226 301096 273232
rect 301136 273216 301188 273222
rect 301136 273158 301188 273164
rect 301148 269090 301176 273158
rect 301148 269062 301360 269090
rect 301332 260658 301360 269062
rect 301240 260630 301360 260658
rect 301240 259434 301268 260630
rect 301148 259406 301268 259434
rect 301148 249898 301176 259406
rect 301136 249892 301188 249898
rect 301136 249834 301188 249840
rect 301044 248464 301096 248470
rect 301044 248406 301096 248412
rect 301056 240174 301084 248406
rect 301044 240168 301096 240174
rect 301044 240110 301096 240116
rect 301136 240168 301188 240174
rect 301136 240110 301188 240116
rect 301148 231878 301176 240110
rect 301136 231872 301188 231878
rect 301136 231814 301188 231820
rect 301228 231804 301280 231810
rect 301228 231746 301280 231752
rect 301240 222222 301268 231746
rect 301044 222216 301096 222222
rect 301044 222158 301096 222164
rect 301228 222216 301280 222222
rect 301228 222158 301280 222164
rect 301056 215354 301084 222158
rect 301044 215348 301096 215354
rect 301044 215290 301096 215296
rect 301136 215212 301188 215218
rect 301136 215154 301188 215160
rect 301148 202910 301176 215154
rect 301044 202904 301096 202910
rect 301044 202846 301096 202852
rect 301136 202904 301188 202910
rect 301136 202846 301188 202852
rect 301056 196042 301084 202846
rect 301044 196036 301096 196042
rect 301044 195978 301096 195984
rect 301136 195900 301188 195906
rect 301136 195842 301188 195848
rect 301148 183598 301176 195842
rect 301044 183592 301096 183598
rect 301044 183534 301096 183540
rect 301136 183592 301188 183598
rect 301136 183534 301188 183540
rect 301056 180810 301084 183534
rect 301044 180804 301096 180810
rect 301044 180746 301096 180752
rect 301044 171148 301096 171154
rect 301044 171090 301096 171096
rect 301056 154578 301084 171090
rect 301056 154550 301176 154578
rect 301148 135266 301176 154550
rect 301056 135238 301176 135266
rect 301056 133890 301084 135238
rect 301044 133884 301096 133890
rect 301044 133826 301096 133832
rect 301136 124228 301188 124234
rect 301136 124170 301188 124176
rect 301148 113286 301176 124170
rect 301136 113280 301188 113286
rect 301136 113222 301188 113228
rect 301044 113212 301096 113218
rect 301044 113154 301096 113160
rect 301056 100042 301084 113154
rect 301056 100014 301268 100042
rect 301240 67658 301268 100014
rect 301044 67652 301096 67658
rect 301044 67594 301096 67600
rect 301228 67652 301280 67658
rect 301228 67594 301280 67600
rect 301056 48346 301084 67594
rect 301044 48340 301096 48346
rect 301044 48282 301096 48288
rect 301136 48204 301188 48210
rect 301136 48146 301188 48152
rect 301148 45506 301176 48146
rect 301148 45478 301268 45506
rect 301240 29034 301268 45478
rect 301136 29028 301188 29034
rect 301136 28970 301188 28976
rect 301228 29028 301280 29034
rect 301228 28970 301280 28976
rect 301148 22250 301176 28970
rect 301148 22222 301268 22250
rect 301240 21978 301268 22222
rect 301056 21950 301268 21978
rect 301056 13598 301084 21950
rect 301044 13592 301096 13598
rect 301044 13534 301096 13540
rect 300952 12436 301004 12442
rect 300952 12378 301004 12384
rect 300860 6112 300912 6118
rect 300860 6054 300912 6060
rect 302252 6050 302280 335650
rect 302344 11694 302372 340054
rect 302712 335714 302740 340054
rect 302700 335708 302752 335714
rect 302700 335650 302752 335656
rect 303080 334762 303108 340054
rect 303160 337952 303212 337958
rect 303160 337894 303212 337900
rect 302516 334756 302568 334762
rect 302516 334698 302568 334704
rect 303068 334756 303120 334762
rect 303068 334698 303120 334704
rect 302528 318850 302556 334698
rect 303172 334642 303200 337894
rect 303620 335640 303672 335646
rect 303620 335582 303672 335588
rect 302896 334614 303200 334642
rect 302516 318844 302568 318850
rect 302516 318786 302568 318792
rect 302608 318844 302660 318850
rect 302608 318786 302660 318792
rect 302620 311982 302648 318786
rect 302608 311976 302660 311982
rect 302608 311918 302660 311924
rect 302516 311840 302568 311846
rect 302516 311782 302568 311788
rect 302528 299538 302556 311782
rect 302516 299532 302568 299538
rect 302516 299474 302568 299480
rect 302608 299532 302660 299538
rect 302608 299474 302660 299480
rect 302620 293298 302648 299474
rect 302528 293270 302648 293298
rect 302528 285002 302556 293270
rect 302528 284974 302740 285002
rect 302712 270570 302740 284974
rect 302516 270564 302568 270570
rect 302516 270506 302568 270512
rect 302700 270564 302752 270570
rect 302700 270506 302752 270512
rect 302528 264330 302556 270506
rect 302528 264302 302740 264330
rect 302712 263514 302740 264302
rect 302620 263486 302740 263514
rect 302620 249830 302648 263486
rect 302516 249824 302568 249830
rect 302516 249766 302568 249772
rect 302608 249824 302660 249830
rect 302608 249766 302660 249772
rect 302528 240174 302556 249766
rect 302516 240168 302568 240174
rect 302516 240110 302568 240116
rect 302700 240168 302752 240174
rect 302700 240110 302752 240116
rect 302712 231946 302740 240110
rect 302700 231940 302752 231946
rect 302700 231882 302752 231888
rect 302608 231804 302660 231810
rect 302608 231746 302660 231752
rect 302620 220833 302648 231746
rect 302606 220824 302662 220833
rect 302606 220759 302662 220768
rect 302514 220688 302570 220697
rect 302514 220623 302570 220632
rect 302528 202910 302556 220623
rect 302516 202904 302568 202910
rect 302516 202846 302568 202852
rect 302608 202904 302660 202910
rect 302608 202846 302660 202852
rect 302620 196110 302648 202846
rect 302608 196104 302660 196110
rect 302608 196046 302660 196052
rect 302516 195968 302568 195974
rect 302516 195910 302568 195916
rect 302528 183598 302556 195910
rect 302516 183592 302568 183598
rect 302516 183534 302568 183540
rect 302608 183592 302660 183598
rect 302608 183534 302660 183540
rect 302620 176798 302648 183534
rect 302608 176792 302660 176798
rect 302608 176734 302660 176740
rect 302608 176656 302660 176662
rect 302608 176598 302660 176604
rect 302620 154578 302648 176598
rect 302528 154550 302648 154578
rect 302528 149818 302556 154550
rect 302528 149790 302740 149818
rect 302712 138582 302740 149790
rect 302516 138576 302568 138582
rect 302516 138518 302568 138524
rect 302700 138576 302752 138582
rect 302700 138518 302752 138524
rect 302528 128330 302556 138518
rect 302528 128302 302648 128330
rect 302620 99498 302648 128302
rect 302528 99470 302648 99498
rect 302528 89570 302556 99470
rect 302528 89542 302648 89570
rect 302620 77314 302648 89542
rect 302516 77308 302568 77314
rect 302516 77250 302568 77256
rect 302608 77308 302660 77314
rect 302608 77250 302660 77256
rect 302528 66230 302556 77250
rect 302516 66224 302568 66230
rect 302516 66166 302568 66172
rect 302700 66224 302752 66230
rect 302700 66166 302752 66172
rect 302712 38672 302740 66166
rect 302528 38644 302740 38672
rect 302528 38570 302556 38644
rect 302528 38542 302648 38570
rect 302620 27606 302648 38542
rect 302516 27600 302568 27606
rect 302516 27542 302568 27548
rect 302608 27600 302660 27606
rect 302608 27542 302660 27548
rect 302528 13666 302556 27542
rect 302516 13660 302568 13666
rect 302516 13602 302568 13608
rect 302332 11688 302384 11694
rect 302332 11630 302384 11636
rect 302240 6044 302292 6050
rect 302240 5986 302292 5992
rect 301412 4412 301464 4418
rect 301412 4354 301464 4360
rect 300308 4140 300360 4146
rect 300308 4082 300360 4088
rect 298100 4072 298152 4078
rect 297364 4004 297416 4010
rect 297836 3998 297956 4026
rect 298100 4014 298152 4020
rect 297364 3946 297416 3952
rect 297928 480 297956 3998
rect 299112 3392 299164 3398
rect 299112 3334 299164 3340
rect 299124 480 299152 3334
rect 300320 480 300348 4082
rect 301424 480 301452 4354
rect 302608 4072 302660 4078
rect 302608 4014 302660 4020
rect 302620 480 302648 4014
rect 302896 3398 302924 334614
rect 303632 5982 303660 335582
rect 303724 11626 303752 340054
rect 304184 335646 304212 340054
rect 304172 335640 304224 335646
rect 304172 335582 304224 335588
rect 304644 331226 304672 340054
rect 305000 335640 305052 335646
rect 305000 335582 305052 335588
rect 303896 331220 303948 331226
rect 303896 331162 303948 331168
rect 304632 331220 304684 331226
rect 304632 331162 304684 331168
rect 303908 311930 303936 331162
rect 303816 311902 303936 311930
rect 303816 311794 303844 311902
rect 303816 311766 303936 311794
rect 303908 292618 303936 311766
rect 303816 292590 303936 292618
rect 303816 292482 303844 292590
rect 303816 292454 303936 292482
rect 303908 215370 303936 292454
rect 303816 215342 303936 215370
rect 303816 215234 303844 215342
rect 303816 215206 303936 215234
rect 303908 196058 303936 215206
rect 303816 196030 303936 196058
rect 303816 195922 303844 196030
rect 303816 195894 303936 195922
rect 303908 176746 303936 195894
rect 303816 176718 303936 176746
rect 303816 176610 303844 176718
rect 303816 176582 303936 176610
rect 303908 144922 303936 176582
rect 303908 144894 304028 144922
rect 304000 132546 304028 144894
rect 303908 132518 304028 132546
rect 303908 122806 303936 132518
rect 303896 122800 303948 122806
rect 303896 122742 303948 122748
rect 303896 113212 303948 113218
rect 303896 113154 303948 113160
rect 303908 85762 303936 113154
rect 303816 85734 303936 85762
rect 303816 85626 303844 85734
rect 303816 85598 303936 85626
rect 303908 74730 303936 85598
rect 303896 74724 303948 74730
rect 303896 74666 303948 74672
rect 303896 74588 303948 74594
rect 303896 74530 303948 74536
rect 303908 63510 303936 74530
rect 303896 63504 303948 63510
rect 303896 63446 303948 63452
rect 303988 53848 304040 53854
rect 303988 53790 304040 53796
rect 304000 45801 304028 53790
rect 303986 45792 304042 45801
rect 303986 45727 304042 45736
rect 303802 45656 303858 45665
rect 303802 45591 303858 45600
rect 303816 42430 303844 45591
rect 303804 42424 303856 42430
rect 303804 42366 303856 42372
rect 304080 42424 304132 42430
rect 304080 42366 304132 42372
rect 304092 34490 304120 42366
rect 304000 34462 304120 34490
rect 304000 26314 304028 34462
rect 303988 26308 304040 26314
rect 303988 26250 304040 26256
rect 303988 24880 304040 24886
rect 303988 24822 304040 24828
rect 304000 13802 304028 24822
rect 303988 13796 304040 13802
rect 303988 13738 304040 13744
rect 303712 11620 303764 11626
rect 303712 11562 303764 11568
rect 303620 5976 303672 5982
rect 303620 5918 303672 5924
rect 305012 5914 305040 335582
rect 305104 11558 305132 340054
rect 305656 335646 305684 340054
rect 306196 338020 306248 338026
rect 306196 337962 306248 337968
rect 305644 335640 305696 335646
rect 305644 335582 305696 335588
rect 306012 123072 306064 123078
rect 306010 123040 306012 123049
rect 306064 123040 306066 123049
rect 306010 122975 306066 122984
rect 305092 11552 305144 11558
rect 305092 11494 305144 11500
rect 305000 5908 305052 5914
rect 305000 5850 305052 5856
rect 305000 4344 305052 4350
rect 305000 4286 305052 4292
rect 302884 3392 302936 3398
rect 302884 3334 302936 3340
rect 303804 3324 303856 3330
rect 303804 3266 303856 3272
rect 303816 480 303844 3266
rect 305012 480 305040 4286
rect 306208 480 306236 337962
rect 306392 333418 306420 340068
rect 306668 340054 306866 340082
rect 307036 340054 307418 340082
rect 307878 340054 307984 340082
rect 306392 333390 306604 333418
rect 306472 333328 306524 333334
rect 306472 333270 306524 333276
rect 306378 157584 306434 157593
rect 306378 157519 306380 157528
rect 306432 157519 306434 157528
rect 306380 157490 306432 157496
rect 306288 110832 306340 110838
rect 306286 110800 306288 110809
rect 306340 110800 306342 110809
rect 306286 110735 306342 110744
rect 306288 28960 306340 28966
rect 306286 28928 306288 28937
rect 306340 28928 306342 28937
rect 306286 28863 306342 28872
rect 306484 11490 306512 333270
rect 306576 13734 306604 333390
rect 306668 333334 306696 340054
rect 306656 333328 306708 333334
rect 306656 333270 306708 333276
rect 307036 331242 307064 340054
rect 307760 335640 307812 335646
rect 307760 335582 307812 335588
rect 306760 331214 307064 331242
rect 306760 318850 306788 331214
rect 306748 318844 306800 318850
rect 306748 318786 306800 318792
rect 306840 318844 306892 318850
rect 306840 318786 306892 318792
rect 306852 317422 306880 318786
rect 306840 317416 306892 317422
rect 306840 317358 306892 317364
rect 306840 299532 306892 299538
rect 306840 299474 306892 299480
rect 306852 292670 306880 299474
rect 306840 292664 306892 292670
rect 306840 292606 306892 292612
rect 306840 292528 306892 292534
rect 306840 292470 306892 292476
rect 306852 275346 306880 292470
rect 306760 275318 306880 275346
rect 306760 264466 306788 275318
rect 306760 264438 306972 264466
rect 306944 263514 306972 264438
rect 306852 263486 306972 263514
rect 306852 254674 306880 263486
rect 306852 254646 306972 254674
rect 306944 249830 306972 254646
rect 306748 249824 306800 249830
rect 306748 249766 306800 249772
rect 306932 249824 306984 249830
rect 306932 249766 306984 249772
rect 306760 248402 306788 249766
rect 306748 248396 306800 248402
rect 306748 248338 306800 248344
rect 306840 240100 306892 240106
rect 306840 240042 306892 240048
rect 306852 238762 306880 240042
rect 306852 238734 306972 238762
rect 306944 231946 306972 238734
rect 306932 231940 306984 231946
rect 306932 231882 306984 231888
rect 306840 231804 306892 231810
rect 306840 231746 306892 231752
rect 306852 220810 306880 231746
rect 306852 220782 306972 220810
rect 306944 213722 306972 220782
rect 306748 213716 306800 213722
rect 306748 213658 306800 213664
rect 306932 213716 306984 213722
rect 306932 213658 306984 213664
rect 306760 202910 306788 213658
rect 306748 202904 306800 202910
rect 306748 202846 306800 202852
rect 306840 202904 306892 202910
rect 306840 202846 306892 202852
rect 306852 201482 306880 202846
rect 306840 201476 306892 201482
rect 306840 201418 306892 201424
rect 306932 201476 306984 201482
rect 306932 201418 306984 201424
rect 306944 183598 306972 201418
rect 306840 183592 306892 183598
rect 306840 183534 306892 183540
rect 306932 183592 306984 183598
rect 306932 183534 306984 183540
rect 306852 180810 306880 183534
rect 306840 180804 306892 180810
rect 306840 180746 306892 180752
rect 306840 171148 306892 171154
rect 306840 171090 306892 171096
rect 306852 161378 306880 171090
rect 306852 161350 306972 161378
rect 306944 154578 306972 161350
rect 306760 154550 306972 154578
rect 306760 149682 306788 154550
rect 306760 149654 306880 149682
rect 306852 135266 306880 149654
rect 306760 135238 306880 135266
rect 306760 128382 306788 135238
rect 306748 128376 306800 128382
rect 306748 128318 306800 128324
rect 306840 128308 306892 128314
rect 306840 128250 306892 128256
rect 306852 115954 306880 128250
rect 306760 115926 306880 115954
rect 306760 109834 306788 115926
rect 306760 109806 306880 109834
rect 306852 99498 306880 109806
rect 306852 99470 306972 99498
rect 306944 85610 306972 99470
rect 306840 85604 306892 85610
rect 306840 85546 306892 85552
rect 306932 85604 306984 85610
rect 306932 85546 306984 85552
rect 306852 77314 306880 85546
rect 306748 77308 306800 77314
rect 306748 77250 306800 77256
rect 306840 77308 306892 77314
rect 306840 77250 306892 77256
rect 306760 66230 306788 77250
rect 306748 66224 306800 66230
rect 306748 66166 306800 66172
rect 306932 66224 306984 66230
rect 306932 66166 306984 66172
rect 306944 40798 306972 66166
rect 306932 40792 306984 40798
rect 306932 40734 306984 40740
rect 306748 35964 306800 35970
rect 306748 35906 306800 35912
rect 306760 31142 306788 35906
rect 306748 31136 306800 31142
rect 306748 31078 306800 31084
rect 306656 26376 306708 26382
rect 306656 26318 306708 26324
rect 306668 24857 306696 26318
rect 306654 24848 306710 24857
rect 306654 24783 306710 24792
rect 307022 24848 307078 24857
rect 307022 24783 307078 24792
rect 307036 15230 307064 24783
rect 306840 15224 306892 15230
rect 306840 15166 306892 15172
rect 307024 15224 307076 15230
rect 307024 15166 307076 15172
rect 306564 13728 306616 13734
rect 306564 13670 306616 13676
rect 306472 11484 306524 11490
rect 306472 11426 306524 11432
rect 306852 6934 306880 15166
rect 306656 6928 306708 6934
rect 306656 6870 306708 6876
rect 306840 6928 306892 6934
rect 306840 6870 306892 6876
rect 306668 5846 306696 6870
rect 306656 5840 306708 5846
rect 306656 5782 306708 5788
rect 307772 5778 307800 335582
rect 307956 13054 307984 340054
rect 308048 340054 308338 340082
rect 308600 340054 308890 340082
rect 309244 340054 309350 340082
rect 309428 340054 309810 340082
rect 310072 340054 310362 340082
rect 310624 340054 310822 340082
rect 311084 340054 311282 340082
rect 311544 340054 311834 340082
rect 312004 340054 312294 340082
rect 312464 340054 312754 340082
rect 307944 13048 307996 13054
rect 307944 12990 307996 12996
rect 308048 11422 308076 340054
rect 308600 335646 308628 340054
rect 308588 335640 308640 335646
rect 308588 335582 308640 335588
rect 309140 335640 309192 335646
rect 309140 335582 309192 335588
rect 309048 134088 309100 134094
rect 309046 134056 309048 134065
rect 309100 134056 309102 134065
rect 309046 133991 309102 134000
rect 308036 11416 308088 11422
rect 308036 11358 308088 11364
rect 307760 5772 307812 5778
rect 307760 5714 307812 5720
rect 309152 5710 309180 335582
rect 309244 9450 309272 340054
rect 309428 11354 309456 340054
rect 309784 338088 309836 338094
rect 309784 338030 309836 338036
rect 309416 11348 309468 11354
rect 309416 11290 309468 11296
rect 309232 9444 309284 9450
rect 309232 9386 309284 9392
rect 309140 5704 309192 5710
rect 309140 5646 309192 5652
rect 308588 4276 308640 4282
rect 308588 4218 308640 4224
rect 307390 3360 307446 3369
rect 307390 3295 307446 3304
rect 307404 480 307432 3295
rect 308600 480 308628 4218
rect 309796 4078 309824 338030
rect 310072 335646 310100 340054
rect 310060 335640 310112 335646
rect 310060 335582 310112 335588
rect 310520 335640 310572 335646
rect 310520 335582 310572 335588
rect 310426 75848 310482 75857
rect 310426 75783 310482 75792
rect 310440 66337 310468 75783
rect 310426 66328 310482 66337
rect 310426 66263 310482 66272
rect 310532 5574 310560 335582
rect 310624 9518 310652 340054
rect 311084 331242 311112 340054
rect 311544 335646 311572 340054
rect 311532 335640 311584 335646
rect 311532 335582 311584 335588
rect 310808 331214 311112 331242
rect 310808 321638 310836 331214
rect 310796 321632 310848 321638
rect 310796 321574 310848 321580
rect 310888 321496 310940 321502
rect 310888 321438 310940 321444
rect 310900 311982 310928 321438
rect 310888 311976 310940 311982
rect 310888 311918 310940 311924
rect 310704 307896 310756 307902
rect 310704 307838 310756 307844
rect 310716 307766 310744 307838
rect 310704 307760 310756 307766
rect 310704 307702 310756 307708
rect 310888 298172 310940 298178
rect 310888 298114 310940 298120
rect 310900 293078 310928 298114
rect 310888 293072 310940 293078
rect 310888 293014 310940 293020
rect 310888 282804 310940 282810
rect 310888 282746 310940 282752
rect 310900 278730 310928 282746
rect 310888 278724 310940 278730
rect 310888 278666 310940 278672
rect 310888 263492 310940 263498
rect 310888 263434 310940 263440
rect 310900 256086 310928 263434
rect 310888 256080 310940 256086
rect 310888 256022 310940 256028
rect 310704 251320 310756 251326
rect 310704 251262 310756 251268
rect 310716 251190 310744 251262
rect 310704 251184 310756 251190
rect 310704 251126 310756 251132
rect 310888 241528 310940 241534
rect 310888 241470 310940 241476
rect 310900 234734 310928 241470
rect 310888 234728 310940 234734
rect 310888 234670 310940 234676
rect 310796 234592 310848 234598
rect 310796 234534 310848 234540
rect 310808 231810 310836 234534
rect 310796 231804 310848 231810
rect 310796 231746 310848 231752
rect 310888 222216 310940 222222
rect 310888 222158 310940 222164
rect 310900 215422 310928 222158
rect 310888 215416 310940 215422
rect 310888 215358 310940 215364
rect 310796 215280 310848 215286
rect 310796 215222 310848 215228
rect 310808 212498 310836 215222
rect 310796 212492 310848 212498
rect 310796 212434 310848 212440
rect 310888 202904 310940 202910
rect 310888 202846 310940 202852
rect 310900 196110 310928 202846
rect 310888 196104 310940 196110
rect 310888 196046 310940 196052
rect 310796 195968 310848 195974
rect 310796 195910 310848 195916
rect 310808 193225 310836 195910
rect 310794 193216 310850 193225
rect 310794 193151 310850 193160
rect 311070 193216 311126 193225
rect 311070 193151 311126 193160
rect 311084 183598 311112 193151
rect 310888 183592 310940 183598
rect 310888 183534 310940 183540
rect 311072 183592 311124 183598
rect 311072 183534 311124 183540
rect 310900 176798 310928 183534
rect 310888 176792 310940 176798
rect 310888 176734 310940 176740
rect 310796 176656 310848 176662
rect 310796 176598 310848 176604
rect 310808 167074 310836 176598
rect 310796 167068 310848 167074
rect 310796 167010 310848 167016
rect 310888 166932 310940 166938
rect 310888 166874 310940 166880
rect 310900 153377 310928 166874
rect 310886 153368 310942 153377
rect 310886 153303 310942 153312
rect 310794 153232 310850 153241
rect 310794 153167 310796 153176
rect 310848 153167 310850 153176
rect 310796 153138 310848 153144
rect 310796 147620 310848 147626
rect 310796 147562 310848 147568
rect 310808 143562 310836 147562
rect 310808 143534 310928 143562
rect 310900 138106 310928 143534
rect 310888 138100 310940 138106
rect 310888 138042 310940 138048
rect 310796 137964 310848 137970
rect 310796 137906 310848 137912
rect 310808 125798 310836 137906
rect 310796 125792 310848 125798
rect 310796 125734 310848 125740
rect 310796 121508 310848 121514
rect 310796 121450 310848 121456
rect 310808 111858 310836 121450
rect 310796 111852 310848 111858
rect 310796 111794 310848 111800
rect 310980 111852 311032 111858
rect 310980 111794 311032 111800
rect 310992 102270 311020 111794
rect 310980 102264 311032 102270
rect 310980 102206 311032 102212
rect 310888 102196 310940 102202
rect 310888 102138 310940 102144
rect 310900 98734 310928 102138
rect 310888 98728 310940 98734
rect 310888 98670 310940 98676
rect 310796 89684 310848 89690
rect 310796 89626 310848 89632
rect 310808 85542 310836 89626
rect 310796 85536 310848 85542
rect 310796 85478 310848 85484
rect 310796 75948 310848 75954
rect 310796 75890 310848 75896
rect 310808 75857 310836 75890
rect 310794 75848 310850 75857
rect 310794 75783 310850 75792
rect 310794 66328 310850 66337
rect 310794 66263 310850 66272
rect 310808 66230 310836 66263
rect 310796 66224 310848 66230
rect 310796 66166 310848 66172
rect 310796 60716 310848 60722
rect 310796 60658 310848 60664
rect 310808 56574 310836 60658
rect 310796 56568 310848 56574
rect 310796 56510 310848 56516
rect 310888 56568 310940 56574
rect 310888 56510 310940 56516
rect 310900 45558 310928 56510
rect 310888 45552 310940 45558
rect 310888 45494 310940 45500
rect 311072 45552 311124 45558
rect 311072 45494 311124 45500
rect 311084 27690 311112 45494
rect 310900 27662 311112 27690
rect 310900 26246 310928 27662
rect 310888 26240 310940 26246
rect 310888 26182 310940 26188
rect 311162 17096 311218 17105
rect 311162 17031 311218 17040
rect 311176 16998 311204 17031
rect 311164 16992 311216 16998
rect 311164 16934 311216 16940
rect 310888 16652 310940 16658
rect 310888 16594 310940 16600
rect 310900 11286 310928 16594
rect 310888 11280 310940 11286
rect 310888 11222 310940 11228
rect 312004 9586 312032 340054
rect 312464 337278 312492 340054
rect 312452 337272 312504 337278
rect 312452 337214 312504 337220
rect 312544 337272 312596 337278
rect 312544 337214 312596 337220
rect 311992 9580 312044 9586
rect 311992 9522 312044 9528
rect 310612 9512 310664 9518
rect 310612 9454 310664 9460
rect 310520 5568 310572 5574
rect 310520 5510 310572 5516
rect 312176 4208 312228 4214
rect 312176 4150 312228 4156
rect 309784 4072 309836 4078
rect 309784 4014 309836 4020
rect 310980 3392 311032 3398
rect 310980 3334 311032 3340
rect 309784 3188 309836 3194
rect 309784 3130 309836 3136
rect 309796 480 309824 3130
rect 310992 480 311020 3334
rect 312188 480 312216 4150
rect 312556 3058 312584 337214
rect 313292 5642 313320 340068
rect 313384 340054 313766 340082
rect 313384 9654 313412 340054
rect 314212 337346 314240 340068
rect 314778 340054 314884 340082
rect 314660 337476 314712 337482
rect 314660 337418 314712 337424
rect 314200 337340 314252 337346
rect 314200 337282 314252 337288
rect 314566 123312 314622 123321
rect 314566 123247 314622 123256
rect 314580 123078 314608 123247
rect 314568 123072 314620 123078
rect 314568 123014 314620 123020
rect 314568 28960 314620 28966
rect 314566 28928 314568 28937
rect 314620 28928 314622 28937
rect 314566 28863 314622 28872
rect 313372 9648 313424 9654
rect 313372 9590 313424 9596
rect 313280 5636 313332 5642
rect 313280 5578 313332 5584
rect 314672 4865 314700 337418
rect 314856 12986 314884 340054
rect 314948 340054 315238 340082
rect 315408 340054 315698 340082
rect 314844 12980 314896 12986
rect 314844 12922 314896 12928
rect 314948 8906 314976 340054
rect 315408 337482 315436 340054
rect 315396 337476 315448 337482
rect 315396 337418 315448 337424
rect 316132 337476 316184 337482
rect 316132 337418 316184 337424
rect 316040 337340 316092 337346
rect 316040 337282 316092 337288
rect 315948 157548 316000 157554
rect 315948 157490 316000 157496
rect 315960 157457 315988 157490
rect 315946 157448 316002 157457
rect 315946 157383 316002 157392
rect 315946 134192 316002 134201
rect 315946 134127 316002 134136
rect 315960 134094 315988 134127
rect 315948 134088 316000 134094
rect 315948 134030 316000 134036
rect 315948 110832 316000 110838
rect 315946 110800 315948 110809
rect 316000 110800 316002 110809
rect 315946 110735 316002 110744
rect 314936 8900 314988 8906
rect 314936 8842 314988 8848
rect 314658 4856 314714 4865
rect 314658 4791 314714 4800
rect 316052 4758 316080 337282
rect 316144 8838 316172 337418
rect 316236 12918 316264 340068
rect 316328 340054 316710 340082
rect 316880 340054 317170 340082
rect 317616 340054 317722 340082
rect 317892 340054 318182 340082
rect 318352 340054 318642 340082
rect 318996 340054 319194 340082
rect 319272 340054 319654 340082
rect 319824 340054 320114 340082
rect 320284 340054 320666 340082
rect 320744 340054 321126 340082
rect 316328 337482 316356 340054
rect 316316 337476 316368 337482
rect 316316 337418 316368 337424
rect 316880 337346 316908 340054
rect 317420 337884 317472 337890
rect 317420 337826 317472 337832
rect 317432 337793 317460 337826
rect 317418 337784 317474 337793
rect 317418 337719 317474 337728
rect 317420 337476 317472 337482
rect 317420 337418 317472 337424
rect 316868 337340 316920 337346
rect 316868 337282 316920 337288
rect 316684 337136 316736 337142
rect 316684 337078 316736 337084
rect 316224 12912 316276 12918
rect 316224 12854 316276 12860
rect 316132 8832 316184 8838
rect 316132 8774 316184 8780
rect 316040 4752 316092 4758
rect 316040 4694 316092 4700
rect 314568 4072 314620 4078
rect 314568 4014 314620 4020
rect 313372 4004 313424 4010
rect 313372 3946 313424 3952
rect 312544 3052 312596 3058
rect 312544 2994 312596 3000
rect 313384 480 313412 3946
rect 314580 480 314608 4014
rect 316696 3262 316724 337078
rect 317326 157720 317382 157729
rect 317326 157655 317382 157664
rect 317340 157457 317368 157655
rect 317326 157448 317382 157457
rect 317326 157383 317382 157392
rect 317326 17096 317382 17105
rect 317326 17031 317382 17040
rect 317340 16697 317368 17031
rect 317326 16688 317382 16697
rect 317326 16623 317382 16632
rect 317432 4690 317460 337418
rect 317512 306400 317564 306406
rect 317512 306342 317564 306348
rect 317524 219434 317552 306342
rect 317512 219428 317564 219434
rect 317512 219370 317564 219376
rect 317512 209840 317564 209846
rect 317512 209782 317564 209788
rect 317524 200122 317552 209782
rect 317512 200116 317564 200122
rect 317512 200058 317564 200064
rect 317512 190528 317564 190534
rect 317512 190470 317564 190476
rect 317524 180810 317552 190470
rect 317512 180804 317564 180810
rect 317512 180746 317564 180752
rect 317512 55276 317564 55282
rect 317512 55218 317564 55224
rect 317524 45558 317552 55218
rect 317512 45552 317564 45558
rect 317512 45494 317564 45500
rect 317512 31816 317564 31822
rect 317512 31758 317564 31764
rect 317524 8770 317552 31758
rect 317616 12850 317644 340054
rect 317892 337770 317920 340054
rect 317708 337742 317920 337770
rect 317708 306406 317736 337742
rect 318352 337482 318380 340054
rect 318340 337476 318392 337482
rect 318340 337418 318392 337424
rect 318892 337476 318944 337482
rect 318892 337418 318944 337424
rect 318800 337340 318852 337346
rect 318800 337282 318852 337288
rect 317696 306400 317748 306406
rect 317696 306342 317748 306348
rect 317696 219428 317748 219434
rect 317696 219370 317748 219376
rect 317708 209846 317736 219370
rect 317696 209840 317748 209846
rect 317696 209782 317748 209788
rect 317696 200116 317748 200122
rect 317696 200058 317748 200064
rect 317708 190534 317736 200058
rect 317696 190528 317748 190534
rect 317696 190470 317748 190476
rect 317696 180804 317748 180810
rect 317696 180746 317748 180752
rect 317708 103426 317736 180746
rect 317696 103420 317748 103426
rect 317696 103362 317748 103368
rect 317788 95260 317840 95266
rect 317788 95202 317840 95208
rect 317800 89758 317828 95202
rect 317788 89752 317840 89758
rect 317788 89694 317840 89700
rect 317880 89616 317932 89622
rect 317880 89558 317932 89564
rect 317892 85490 317920 89558
rect 317892 85462 318012 85490
rect 317984 75954 318012 85462
rect 317696 75948 317748 75954
rect 317696 75890 317748 75896
rect 317972 75948 318024 75954
rect 317972 75890 318024 75896
rect 317708 55282 317736 75890
rect 317696 55276 317748 55282
rect 317696 55218 317748 55224
rect 317696 45552 317748 45558
rect 317696 45494 317748 45500
rect 317708 31822 317736 45494
rect 317696 31816 317748 31822
rect 317696 31758 317748 31764
rect 317604 12844 317656 12850
rect 317604 12786 317656 12792
rect 317512 8764 317564 8770
rect 317512 8706 317564 8712
rect 318708 4752 318760 4758
rect 318708 4694 318760 4700
rect 317420 4684 317472 4690
rect 317420 4626 317472 4632
rect 318720 3466 318748 4694
rect 318812 4622 318840 337282
rect 318904 8702 318932 337418
rect 318996 12782 319024 340054
rect 319272 337482 319300 340054
rect 319260 337476 319312 337482
rect 319260 337418 319312 337424
rect 319824 337346 319852 340054
rect 320180 337476 320232 337482
rect 320180 337418 320232 337424
rect 319812 337340 319864 337346
rect 319812 337282 319864 337288
rect 319444 337000 319496 337006
rect 319444 336942 319496 336948
rect 318984 12776 319036 12782
rect 318984 12718 319036 12724
rect 318892 8696 318944 8702
rect 318892 8638 318944 8644
rect 318800 4616 318852 4622
rect 318800 4558 318852 4564
rect 318708 3460 318760 3466
rect 318708 3402 318760 3408
rect 316684 3256 316736 3262
rect 316684 3198 316736 3204
rect 318064 3256 318116 3262
rect 318064 3198 318116 3204
rect 315764 3052 315816 3058
rect 315764 2994 315816 3000
rect 315776 480 315804 2994
rect 316960 2984 317012 2990
rect 316960 2926 317012 2932
rect 316972 480 317000 2926
rect 318076 480 318104 3198
rect 319456 3126 319484 336942
rect 320192 8634 320220 337418
rect 320284 12714 320312 340054
rect 320744 337482 320772 340054
rect 320732 337476 320784 337482
rect 320732 337418 320784 337424
rect 321468 337340 321520 337346
rect 321468 337282 321520 337288
rect 320272 12708 320324 12714
rect 320272 12650 320324 12656
rect 320180 8628 320232 8634
rect 320180 8570 320232 8576
rect 321480 4808 321508 337282
rect 321204 4780 321508 4808
rect 320364 4548 320416 4554
rect 320364 4490 320416 4496
rect 320376 3534 320404 4490
rect 321204 3534 321232 4780
rect 321572 4706 321600 340068
rect 321756 340054 322138 340082
rect 322216 340054 322598 340082
rect 322952 340054 323058 340082
rect 323136 340054 323518 340082
rect 323688 340054 324070 340082
rect 324332 340054 324530 340082
rect 324700 340054 324990 340082
rect 321652 335640 321704 335646
rect 321652 335582 321704 335588
rect 321664 8566 321692 335582
rect 321756 12646 321784 340054
rect 322216 335646 322244 340054
rect 322204 335640 322256 335646
rect 322204 335582 322256 335588
rect 322202 16824 322258 16833
rect 322202 16759 322258 16768
rect 322216 16425 322244 16759
rect 322202 16416 322258 16425
rect 322202 16351 322258 16360
rect 321744 12640 321796 12646
rect 321744 12582 321796 12588
rect 321652 8560 321704 8566
rect 321652 8502 321704 8508
rect 321652 5092 321704 5098
rect 321652 5034 321704 5040
rect 321664 4962 321692 5034
rect 321652 4956 321704 4962
rect 321652 4898 321704 4904
rect 321388 4678 321600 4706
rect 321388 4622 321416 4678
rect 321376 4616 321428 4622
rect 321376 4558 321428 4564
rect 322756 4616 322808 4622
rect 322756 4558 322808 4564
rect 320364 3528 320416 3534
rect 320364 3470 320416 3476
rect 320456 3528 320508 3534
rect 320456 3470 320508 3476
rect 321192 3528 321244 3534
rect 321192 3470 321244 3476
rect 321652 3528 321704 3534
rect 321652 3470 321704 3476
rect 319444 3120 319496 3126
rect 319444 3062 319496 3068
rect 319260 2916 319312 2922
rect 319260 2858 319312 2864
rect 319272 480 319300 2858
rect 320468 480 320496 3470
rect 321664 480 321692 3470
rect 322768 3466 322796 4558
rect 322952 4486 322980 340054
rect 323136 12578 323164 340054
rect 323688 336734 323716 340054
rect 323676 336728 323728 336734
rect 323676 336670 323728 336676
rect 323308 327140 323360 327146
rect 323308 327082 323360 327088
rect 323320 311982 323348 327082
rect 323308 311976 323360 311982
rect 323308 311918 323360 311924
rect 323216 311908 323268 311914
rect 323216 311850 323268 311856
rect 323228 304298 323256 311850
rect 323216 304292 323268 304298
rect 323216 304234 323268 304240
rect 323308 299532 323360 299538
rect 323308 299474 323360 299480
rect 323320 296721 323348 299474
rect 323306 296712 323362 296721
rect 323306 296647 323362 296656
rect 323490 296712 323546 296721
rect 323490 296647 323546 296656
rect 323504 287094 323532 296647
rect 323308 287088 323360 287094
rect 323492 287088 323544 287094
rect 323360 287036 323440 287042
rect 323308 287030 323440 287036
rect 323492 287030 323544 287036
rect 323320 287014 323440 287030
rect 323412 280242 323440 287014
rect 323412 280214 323532 280242
rect 323504 279970 323532 280214
rect 323320 279942 323532 279970
rect 323320 273358 323348 279942
rect 323308 273352 323360 273358
rect 323308 273294 323360 273300
rect 323308 267776 323360 267782
rect 323308 267718 323360 267724
rect 323320 260930 323348 267718
rect 323320 260902 323440 260930
rect 323412 259434 323440 260902
rect 323320 259406 323440 259434
rect 323320 253978 323348 259406
rect 323308 253972 323360 253978
rect 323308 253914 323360 253920
rect 323400 249824 323452 249830
rect 323400 249766 323452 249772
rect 323412 233918 323440 249766
rect 323400 233912 323452 233918
rect 323400 233854 323452 233860
rect 323584 233912 323636 233918
rect 323584 233854 323636 233860
rect 323596 229129 323624 233854
rect 323398 229120 323454 229129
rect 323398 229055 323454 229064
rect 323582 229120 323638 229129
rect 323582 229055 323638 229064
rect 323412 200127 323440 229055
rect 323398 200118 323454 200127
rect 323398 200053 323454 200062
rect 323398 199880 323454 199889
rect 323398 199815 323454 199824
rect 323412 190482 323440 199815
rect 323412 190454 323532 190482
rect 323504 173942 323532 190454
rect 323308 173936 323360 173942
rect 323308 173878 323360 173884
rect 323492 173936 323544 173942
rect 323492 173878 323544 173884
rect 323320 164234 323348 173878
rect 323320 164206 323440 164234
rect 323412 157434 323440 164206
rect 323412 157406 323532 157434
rect 323504 155258 323532 157406
rect 323412 155230 323532 155258
rect 323412 144906 323440 155230
rect 323400 144900 323452 144906
rect 323400 144842 323452 144848
rect 323492 144900 323544 144906
rect 323492 144842 323544 144848
rect 323504 135289 323532 144842
rect 323306 135280 323362 135289
rect 323306 135215 323362 135224
rect 323490 135280 323546 135289
rect 323490 135215 323546 135224
rect 323320 125610 323348 135215
rect 323320 125582 323440 125610
rect 323412 118810 323440 125582
rect 323412 118782 323532 118810
rect 323504 118130 323532 118782
rect 323412 118102 323532 118130
rect 323412 108050 323440 118102
rect 323400 108044 323452 108050
rect 323400 107986 323452 107992
rect 323400 95260 323452 95266
rect 323400 95202 323452 95208
rect 323412 86970 323440 95202
rect 323308 86964 323360 86970
rect 323308 86906 323360 86912
rect 323400 86964 323452 86970
rect 323400 86906 323452 86912
rect 323320 72434 323348 86906
rect 323320 72406 323440 72434
rect 323412 66230 323440 72406
rect 323400 66224 323452 66230
rect 323400 66166 323452 66172
rect 323400 56636 323452 56642
rect 323400 56578 323452 56584
rect 323412 48278 323440 56578
rect 323308 48272 323360 48278
rect 323308 48214 323360 48220
rect 323400 48272 323452 48278
rect 323400 48214 323452 48220
rect 323320 46918 323348 48214
rect 323308 46912 323360 46918
rect 323308 46854 323360 46860
rect 323308 37324 323360 37330
rect 323308 37266 323360 37272
rect 323320 33810 323348 37266
rect 323320 33782 323532 33810
rect 323504 31634 323532 33782
rect 323412 31606 323532 31634
rect 323412 28966 323440 31606
rect 323308 28960 323360 28966
rect 323308 28902 323360 28908
rect 323400 28960 323452 28966
rect 323400 28902 323452 28908
rect 323124 12572 323176 12578
rect 323124 12514 323176 12520
rect 323320 8498 323348 28902
rect 323308 8492 323360 8498
rect 323308 8434 323360 8440
rect 324332 4894 324360 340054
rect 324700 335730 324728 340054
rect 324424 335702 324728 335730
rect 324424 7614 324452 335702
rect 325068 327146 325096 340190
rect 325712 340054 326002 340082
rect 326080 340054 326462 340082
rect 326632 340054 327014 340082
rect 327092 340054 327474 340082
rect 324688 327140 324740 327146
rect 324688 327082 324740 327088
rect 325056 327140 325108 327146
rect 325056 327082 325108 327088
rect 324700 311930 324728 327082
rect 324608 311902 324728 311930
rect 324608 302138 324636 311902
rect 324608 302110 324728 302138
rect 324700 299470 324728 302110
rect 324688 299464 324740 299470
rect 324688 299406 324740 299412
rect 324688 289876 324740 289882
rect 324688 289818 324740 289824
rect 324700 285274 324728 289818
rect 324700 285246 324820 285274
rect 324792 277409 324820 285246
rect 324502 277400 324558 277409
rect 324502 277335 324558 277344
rect 324778 277400 324834 277409
rect 324778 277335 324834 277344
rect 324516 267850 324544 277335
rect 324504 267844 324556 267850
rect 324504 267786 324556 267792
rect 324688 267844 324740 267850
rect 324688 267786 324740 267792
rect 324700 267730 324728 267786
rect 324608 267702 324728 267730
rect 324608 260914 324636 267702
rect 324596 260908 324648 260914
rect 324596 260850 324648 260856
rect 324596 258120 324648 258126
rect 324596 258062 324648 258068
rect 324608 238785 324636 258062
rect 324594 238776 324650 238785
rect 324594 238711 324650 238720
rect 324778 238776 324834 238785
rect 324778 238711 324834 238720
rect 324792 231878 324820 238711
rect 324688 231872 324740 231878
rect 324686 231840 324688 231849
rect 324780 231872 324832 231878
rect 324740 231840 324742 231849
rect 324780 231814 324832 231820
rect 324686 231775 324742 231784
rect 324778 231704 324834 231713
rect 324778 231639 324834 231648
rect 324792 212566 324820 231639
rect 324688 212560 324740 212566
rect 324608 212508 324688 212514
rect 324608 212502 324740 212508
rect 324780 212560 324832 212566
rect 324780 212502 324832 212508
rect 324608 212486 324728 212502
rect 324608 201482 324636 212486
rect 324596 201476 324648 201482
rect 324596 201418 324648 201424
rect 324688 193180 324740 193186
rect 324688 193122 324740 193128
rect 324700 191842 324728 193122
rect 324700 191814 324820 191842
rect 324792 183598 324820 191814
rect 324596 183592 324648 183598
rect 324596 183534 324648 183540
rect 324780 183592 324832 183598
rect 324780 183534 324832 183540
rect 324608 173942 324636 183534
rect 324596 173936 324648 173942
rect 324596 173878 324648 173884
rect 324688 173936 324740 173942
rect 324688 173878 324740 173884
rect 324700 164234 324728 173878
rect 324608 164206 324728 164234
rect 324608 157434 324636 164206
rect 324516 157406 324636 157434
rect 324516 157298 324544 157406
rect 324516 157270 324636 157298
rect 324608 144906 324636 157270
rect 324596 144900 324648 144906
rect 324596 144842 324648 144848
rect 324780 144900 324832 144906
rect 324780 144842 324832 144848
rect 324792 139942 324820 144842
rect 324780 139936 324832 139942
rect 324780 139878 324832 139884
rect 324780 133952 324832 133958
rect 324780 133894 324832 133900
rect 324792 125633 324820 133894
rect 324594 125624 324650 125633
rect 324594 125559 324650 125568
rect 324778 125624 324834 125633
rect 324778 125559 324834 125568
rect 324608 122806 324636 125559
rect 325606 123584 325662 123593
rect 325606 123519 325662 123528
rect 325620 123049 325648 123519
rect 325606 123040 325662 123049
rect 325606 122975 325662 122984
rect 324596 122800 324648 122806
rect 324596 122742 324648 122748
rect 324596 113212 324648 113218
rect 324596 113154 324648 113160
rect 324608 104854 324636 113154
rect 325606 111072 325662 111081
rect 325606 111007 325662 111016
rect 325620 110809 325648 111007
rect 325606 110800 325662 110809
rect 325606 110735 325662 110744
rect 324596 104848 324648 104854
rect 324596 104790 324648 104796
rect 324596 95260 324648 95266
rect 324596 95202 324648 95208
rect 324608 86970 324636 95202
rect 324596 86964 324648 86970
rect 324596 86906 324648 86912
rect 324688 86896 324740 86902
rect 324688 86838 324740 86844
rect 324700 67674 324728 86838
rect 324608 67646 324728 67674
rect 324608 60858 324636 67646
rect 324596 60852 324648 60858
rect 324596 60794 324648 60800
rect 324596 60716 324648 60722
rect 324596 60658 324648 60664
rect 324608 38690 324636 60658
rect 324596 38684 324648 38690
rect 324596 38626 324648 38632
rect 324688 38684 324740 38690
rect 324688 38626 324740 38632
rect 324700 28966 324728 38626
rect 325606 29200 325662 29209
rect 325606 29135 325662 29144
rect 324596 28960 324648 28966
rect 324596 28902 324648 28908
rect 324688 28960 324740 28966
rect 325620 28937 325648 29135
rect 324688 28902 324740 28908
rect 325606 28928 325662 28937
rect 324608 8430 324636 28902
rect 325606 28863 325662 28872
rect 324596 8424 324648 8430
rect 324596 8366 324648 8372
rect 324412 7608 324464 7614
rect 324412 7550 324464 7556
rect 324320 4888 324372 4894
rect 324320 4830 324372 4836
rect 325712 4826 325740 340054
rect 326080 335594 326108 340054
rect 325804 335566 326108 335594
rect 325804 7682 325832 335566
rect 326632 327146 326660 340054
rect 326988 337884 327040 337890
rect 326988 337826 327040 337832
rect 327000 337793 327028 337826
rect 326986 337784 327042 337793
rect 326986 337719 327042 337728
rect 325976 327140 326028 327146
rect 325976 327082 326028 327088
rect 326620 327140 326672 327146
rect 326620 327082 326672 327088
rect 325988 302274 326016 327082
rect 325896 302246 326016 302274
rect 325896 299470 325924 302246
rect 325884 299464 325936 299470
rect 325884 299406 325936 299412
rect 325976 299396 326028 299402
rect 325976 299338 326028 299344
rect 325988 287026 326016 299338
rect 325976 287020 326028 287026
rect 325976 286962 326028 286968
rect 326068 287020 326120 287026
rect 326068 286962 326120 286968
rect 326080 267782 326108 286962
rect 325976 267776 326028 267782
rect 325976 267718 326028 267724
rect 326068 267776 326120 267782
rect 326068 267718 326120 267724
rect 325988 262970 326016 267718
rect 325988 262942 326108 262970
rect 326080 231878 326108 262942
rect 325976 231872 326028 231878
rect 325976 231814 326028 231820
rect 326068 231872 326120 231878
rect 326068 231814 326120 231820
rect 325988 222290 326016 231814
rect 325976 222284 326028 222290
rect 325976 222226 326028 222232
rect 325884 222216 325936 222222
rect 325884 222158 325936 222164
rect 325896 212566 325924 222158
rect 325884 212560 325936 212566
rect 325884 212502 325936 212508
rect 325976 212560 326028 212566
rect 325976 212502 326028 212508
rect 325988 202978 326016 212502
rect 325976 202972 326028 202978
rect 325976 202914 326028 202920
rect 325884 202904 325936 202910
rect 325882 202872 325884 202881
rect 325936 202872 325938 202881
rect 325882 202807 325938 202816
rect 325974 202736 326030 202745
rect 325974 202671 326030 202680
rect 325988 188442 326016 202671
rect 325896 188414 326016 188442
rect 325896 173942 325924 188414
rect 325884 173936 325936 173942
rect 325884 173878 325936 173884
rect 325976 173936 326028 173942
rect 325976 173878 326028 173884
rect 325988 164234 326016 173878
rect 325896 164206 326016 164234
rect 325896 157978 325924 164206
rect 325896 157950 326016 157978
rect 325988 157282 326016 157950
rect 325976 157276 326028 157282
rect 325976 157218 326028 157224
rect 325976 157140 326028 157146
rect 325976 157082 326028 157088
rect 325988 149818 326016 157082
rect 325988 149790 326108 149818
rect 326080 144945 326108 149790
rect 325882 144936 325938 144945
rect 325882 144871 325884 144880
rect 325936 144871 325938 144880
rect 326066 144936 326122 144945
rect 326066 144871 326068 144880
rect 325884 144842 325936 144848
rect 326120 144871 326122 144880
rect 326068 144842 326120 144848
rect 326080 137766 326108 144842
rect 326068 137760 326120 137766
rect 326068 137702 326120 137708
rect 326068 133952 326120 133958
rect 326068 133894 326120 133900
rect 326080 125633 326108 133894
rect 325882 125624 325938 125633
rect 325882 125559 325938 125568
rect 326066 125624 326122 125633
rect 326066 125559 326122 125568
rect 325896 122806 325924 125559
rect 325884 122800 325936 122806
rect 325884 122742 325936 122748
rect 326068 114436 326120 114442
rect 326068 114378 326120 114384
rect 326080 104922 326108 114378
rect 325976 104916 326028 104922
rect 325976 104858 326028 104864
rect 326068 104916 326120 104922
rect 326068 104858 326120 104864
rect 325988 67674 326016 104858
rect 325896 67646 326016 67674
rect 325896 60790 325924 67646
rect 325884 60784 325936 60790
rect 325884 60726 325936 60732
rect 325976 60648 326028 60654
rect 325976 60590 326028 60596
rect 325988 53258 326016 60590
rect 325988 53230 326108 53258
rect 326080 48346 326108 53230
rect 325884 48340 325936 48346
rect 325884 48282 325936 48288
rect 326068 48340 326120 48346
rect 326068 48282 326120 48288
rect 325896 38758 325924 48282
rect 325884 38752 325936 38758
rect 325884 38694 325936 38700
rect 325884 38616 325936 38622
rect 325884 38558 325936 38564
rect 325896 28966 325924 38558
rect 326986 29336 327042 29345
rect 326986 29271 327042 29280
rect 325884 28960 325936 28966
rect 325884 28902 325936 28908
rect 325976 28960 326028 28966
rect 327000 28937 327028 29271
rect 325976 28902 326028 28908
rect 326986 28928 327042 28937
rect 325988 8974 326016 28902
rect 326986 28863 327042 28872
rect 325976 8968 326028 8974
rect 325976 8910 326028 8916
rect 325792 7676 325844 7682
rect 325792 7618 325844 7624
rect 327092 5098 327120 340054
rect 327920 338434 327948 340068
rect 328486 340054 328684 340082
rect 327356 338428 327408 338434
rect 327356 338370 327408 338376
rect 327908 338428 327960 338434
rect 327908 338370 327960 338376
rect 327170 337784 327226 337793
rect 327170 337719 327172 337728
rect 327224 337719 327226 337728
rect 327172 337690 327224 337696
rect 327368 331106 327396 338370
rect 327724 336932 327776 336938
rect 327724 336874 327776 336880
rect 327276 331078 327396 331106
rect 327276 327078 327304 331078
rect 327264 327072 327316 327078
rect 327264 327014 327316 327020
rect 327264 317484 327316 317490
rect 327264 317426 327316 317432
rect 327276 317370 327304 317426
rect 327184 317342 327304 317370
rect 327184 309194 327212 317342
rect 327172 309188 327224 309194
rect 327172 309130 327224 309136
rect 327172 309052 327224 309058
rect 327172 308994 327224 309000
rect 327184 280226 327212 308994
rect 327172 280220 327224 280226
rect 327172 280162 327224 280168
rect 327172 278792 327224 278798
rect 327172 278734 327224 278740
rect 327184 270570 327212 278734
rect 327172 270564 327224 270570
rect 327172 270506 327224 270512
rect 327264 270564 327316 270570
rect 327264 270506 327316 270512
rect 327276 260982 327304 270506
rect 327264 260976 327316 260982
rect 327264 260918 327316 260924
rect 327172 260772 327224 260778
rect 327172 260714 327224 260720
rect 327184 259457 327212 260714
rect 327170 259448 327226 259457
rect 327170 259383 327226 259392
rect 327354 259312 327410 259321
rect 327354 259247 327410 259256
rect 327368 231878 327396 259247
rect 327264 231872 327316 231878
rect 327264 231814 327316 231820
rect 327356 231872 327408 231878
rect 327356 231814 327408 231820
rect 327276 222290 327304 231814
rect 327264 222284 327316 222290
rect 327264 222226 327316 222232
rect 327172 222216 327224 222222
rect 327172 222158 327224 222164
rect 327184 212566 327212 222158
rect 327172 212560 327224 212566
rect 327172 212502 327224 212508
rect 327264 212560 327316 212566
rect 327264 212502 327316 212508
rect 327276 202978 327304 212502
rect 327264 202972 327316 202978
rect 327264 202914 327316 202920
rect 327172 202904 327224 202910
rect 327172 202846 327224 202852
rect 327184 201482 327212 202846
rect 327172 201476 327224 201482
rect 327172 201418 327224 201424
rect 327264 193180 327316 193186
rect 327264 193122 327316 193128
rect 327276 191842 327304 193122
rect 327276 191814 327396 191842
rect 327368 183598 327396 191814
rect 327172 183592 327224 183598
rect 327172 183534 327224 183540
rect 327356 183592 327408 183598
rect 327356 183534 327408 183540
rect 327184 173942 327212 183534
rect 327172 173936 327224 173942
rect 327172 173878 327224 173884
rect 327264 173936 327316 173942
rect 327264 173878 327316 173884
rect 327276 166138 327304 173878
rect 327276 166110 327488 166138
rect 327460 162897 327488 166110
rect 327262 162888 327318 162897
rect 327262 162823 327318 162832
rect 327446 162888 327502 162897
rect 327446 162823 327502 162832
rect 327276 148458 327304 162823
rect 327276 148430 327396 148458
rect 327368 137714 327396 148430
rect 327276 137686 327396 137714
rect 327276 130370 327304 137686
rect 327184 130342 327304 130370
rect 327184 113393 327212 130342
rect 327170 113384 327226 113393
rect 327170 113319 327226 113328
rect 327170 113248 327226 113257
rect 327170 113183 327226 113192
rect 327184 103494 327212 113183
rect 327172 103488 327224 103494
rect 327172 103430 327224 103436
rect 327172 96620 327224 96626
rect 327172 96562 327224 96568
rect 327184 86970 327212 96562
rect 327172 86964 327224 86970
rect 327172 86906 327224 86912
rect 327264 86896 327316 86902
rect 327264 86838 327316 86844
rect 327276 70514 327304 86838
rect 327264 70508 327316 70514
rect 327264 70450 327316 70456
rect 327172 70372 327224 70378
rect 327172 70314 327224 70320
rect 327184 66230 327212 70314
rect 327172 66224 327224 66230
rect 327172 66166 327224 66172
rect 327448 56636 327500 56642
rect 327448 56578 327500 56584
rect 327460 56522 327488 56578
rect 327368 56494 327488 56522
rect 327368 48346 327396 56494
rect 327356 48340 327408 48346
rect 327356 48282 327408 48288
rect 327356 46980 327408 46986
rect 327356 46922 327408 46928
rect 327368 38690 327396 46922
rect 327264 38684 327316 38690
rect 327264 38626 327316 38632
rect 327356 38684 327408 38690
rect 327356 38626 327408 38632
rect 327276 7002 327304 38626
rect 327264 6996 327316 7002
rect 327264 6938 327316 6944
rect 327080 5092 327132 5098
rect 327080 5034 327132 5040
rect 327080 4956 327132 4962
rect 327080 4898 327132 4904
rect 326344 4888 326396 4894
rect 326344 4830 326396 4836
rect 325700 4820 325752 4826
rect 325700 4762 325752 4768
rect 323308 4752 323360 4758
rect 323308 4694 323360 4700
rect 322940 4480 322992 4486
rect 322940 4422 322992 4428
rect 322848 3596 322900 3602
rect 322848 3538 322900 3544
rect 322756 3460 322808 3466
rect 322756 3402 322808 3408
rect 322860 480 322888 3538
rect 323320 3058 323348 4694
rect 325148 4480 325200 4486
rect 325148 4422 325200 4428
rect 325160 3670 325188 4422
rect 325148 3664 325200 3670
rect 325148 3606 325200 3612
rect 325240 3664 325292 3670
rect 325240 3606 325292 3612
rect 324044 3460 324096 3466
rect 324044 3402 324096 3408
rect 323308 3052 323360 3058
rect 323308 2994 323360 3000
rect 324056 480 324084 3402
rect 325252 480 325280 3606
rect 326356 2922 326384 4830
rect 326436 3732 326488 3738
rect 326436 3674 326488 3680
rect 326344 2916 326396 2922
rect 326344 2858 326396 2864
rect 326448 480 326476 3674
rect 327092 3602 327120 4898
rect 327080 3596 327132 3602
rect 327080 3538 327132 3544
rect 327736 3126 327764 336874
rect 328552 331696 328604 331702
rect 328552 331638 328604 331644
rect 328458 134192 328514 134201
rect 328458 134127 328514 134136
rect 328472 133929 328500 134127
rect 328458 133920 328514 133929
rect 328458 133855 328514 133864
rect 328458 123176 328514 123185
rect 328458 123111 328514 123120
rect 328472 123049 328500 123111
rect 328458 123040 328514 123049
rect 328458 122975 328514 122984
rect 328564 7750 328592 331638
rect 328656 9042 328684 340054
rect 328748 340054 328946 340082
rect 329024 340054 329406 340082
rect 329958 340054 330064 340082
rect 328644 9036 328696 9042
rect 328644 8978 328696 8984
rect 328552 7744 328604 7750
rect 328552 7686 328604 7692
rect 328748 5030 328776 340054
rect 329024 331702 329052 340054
rect 329840 335640 329892 335646
rect 329840 335582 329892 335588
rect 329012 331696 329064 331702
rect 329012 331638 329064 331644
rect 329852 5098 329880 335582
rect 329932 278928 329984 278934
rect 329932 278870 329984 278876
rect 329944 267782 329972 278870
rect 329932 267776 329984 267782
rect 329932 267718 329984 267724
rect 330036 249898 330064 340054
rect 330128 340054 330418 340082
rect 330588 340054 330878 340082
rect 330128 335646 330156 340054
rect 330116 335640 330168 335646
rect 330116 335582 330168 335588
rect 330588 331786 330616 340054
rect 331312 335708 331364 335714
rect 331312 335650 331364 335656
rect 331220 335640 331272 335646
rect 331220 335582 331272 335588
rect 330220 331758 330616 331786
rect 330220 317422 330248 331758
rect 330208 317416 330260 317422
rect 330208 317358 330260 317364
rect 330208 307828 330260 307834
rect 330208 307770 330260 307776
rect 330220 299554 330248 307770
rect 330128 299526 330248 299554
rect 330128 288454 330156 299526
rect 330116 288448 330168 288454
rect 330116 288390 330168 288396
rect 330208 288448 330260 288454
rect 330208 288390 330260 288396
rect 330220 278934 330248 288390
rect 330208 278928 330260 278934
rect 330208 278870 330260 278876
rect 330116 267776 330168 267782
rect 330116 267718 330168 267724
rect 330128 258058 330156 267718
rect 330116 258052 330168 258058
rect 330116 257994 330168 258000
rect 330300 258052 330352 258058
rect 330300 257994 330352 258000
rect 330024 249892 330076 249898
rect 330024 249834 330076 249840
rect 330024 249756 330076 249762
rect 330024 249698 330076 249704
rect 329930 248432 329986 248441
rect 329930 248367 329986 248376
rect 329944 245002 329972 248367
rect 329932 244996 329984 245002
rect 329932 244938 329984 244944
rect 329932 182096 329984 182102
rect 329932 182038 329984 182044
rect 329944 172553 329972 182038
rect 329930 172544 329986 172553
rect 329930 172479 329932 172488
rect 329984 172479 329986 172488
rect 329932 172450 329984 172456
rect 329944 162897 329972 172450
rect 329930 162888 329986 162897
rect 329930 162823 329986 162832
rect 329932 143540 329984 143546
rect 329932 143482 329984 143488
rect 329944 125633 329972 143482
rect 329930 125624 329986 125633
rect 329930 125559 329986 125568
rect 329932 84244 329984 84250
rect 329932 84186 329984 84192
rect 329944 67658 329972 84186
rect 330036 77382 330064 249698
rect 330312 248441 330340 257994
rect 330298 248432 330354 248441
rect 330298 248367 330354 248376
rect 330208 244996 330260 245002
rect 330208 244938 330260 244944
rect 330220 240145 330248 244938
rect 330206 240136 330262 240145
rect 330206 240071 330262 240080
rect 330390 240136 330446 240145
rect 330390 240071 330446 240080
rect 330404 230518 330432 240071
rect 330208 230512 330260 230518
rect 330208 230454 330260 230460
rect 330392 230512 330444 230518
rect 330392 230454 330444 230460
rect 330128 222222 330156 222253
rect 330220 222222 330248 230454
rect 330116 222216 330168 222222
rect 330208 222216 330260 222222
rect 330168 222164 330208 222170
rect 330116 222158 330260 222164
rect 330128 222142 330248 222158
rect 330220 212634 330248 222142
rect 330208 212628 330260 212634
rect 330208 212570 330260 212576
rect 330208 212492 330260 212498
rect 330208 212434 330260 212440
rect 330220 211154 330248 212434
rect 330220 211138 330340 211154
rect 330220 211132 330352 211138
rect 330220 211126 330300 211132
rect 330300 211074 330352 211080
rect 330312 211043 330340 211074
rect 330116 202836 330168 202842
rect 330116 202778 330168 202784
rect 330128 201482 330156 202778
rect 330116 201476 330168 201482
rect 330116 201418 330168 201424
rect 330300 201476 330352 201482
rect 330300 201418 330352 201424
rect 330312 200122 330340 201418
rect 330300 200116 330352 200122
rect 330300 200058 330352 200064
rect 330484 200116 330536 200122
rect 330484 200058 330536 200064
rect 330496 190505 330524 200058
rect 330298 190496 330354 190505
rect 330298 190431 330354 190440
rect 330482 190496 330538 190505
rect 330482 190431 330538 190440
rect 330312 182209 330340 190431
rect 330114 182200 330170 182209
rect 330114 182135 330170 182144
rect 330298 182200 330354 182209
rect 330298 182135 330354 182144
rect 330128 182102 330156 182135
rect 330116 182096 330168 182102
rect 330116 182038 330168 182044
rect 330206 172544 330262 172553
rect 330206 172479 330208 172488
rect 330260 172479 330262 172488
rect 330208 172450 330260 172456
rect 330114 162888 330170 162897
rect 330114 162823 330170 162832
rect 330128 162790 330156 162823
rect 330116 162784 330168 162790
rect 330116 162726 330168 162732
rect 330208 144968 330260 144974
rect 330208 144910 330260 144916
rect 330220 143546 330248 144910
rect 330208 143540 330260 143546
rect 330208 143482 330260 143488
rect 330114 125624 330170 125633
rect 330114 125559 330116 125568
rect 330168 125559 330170 125568
rect 330300 125588 330352 125594
rect 330116 125530 330168 125536
rect 330300 125530 330352 125536
rect 330312 114492 330340 125530
rect 330128 114464 330340 114492
rect 330128 103426 330156 114464
rect 330116 103420 330168 103426
rect 330116 103362 330168 103368
rect 330208 98728 330260 98734
rect 330208 98670 330260 98676
rect 330220 93922 330248 98670
rect 330128 93894 330248 93922
rect 330128 93838 330156 93894
rect 330116 93832 330168 93838
rect 330116 93774 330168 93780
rect 330024 77376 330076 77382
rect 330024 77318 330076 77324
rect 330024 77240 330076 77246
rect 330024 77182 330076 77188
rect 329932 67652 329984 67658
rect 329932 67594 329984 67600
rect 329930 48240 329986 48249
rect 329930 48175 329986 48184
rect 329944 38690 329972 48175
rect 329932 38684 329984 38690
rect 329932 38626 329984 38632
rect 329932 26308 329984 26314
rect 329932 26250 329984 26256
rect 329944 25906 329972 26250
rect 329932 25900 329984 25906
rect 329932 25842 329984 25848
rect 330036 9110 330064 77182
rect 330116 67652 330168 67658
rect 330116 67594 330168 67600
rect 330128 61470 330156 67594
rect 330116 61464 330168 61470
rect 330116 61406 330168 61412
rect 330300 57860 330352 57866
rect 330300 57802 330352 57808
rect 330312 48385 330340 57802
rect 330298 48376 330354 48385
rect 330298 48311 330354 48320
rect 331126 48240 331182 48249
rect 331126 48175 331182 48184
rect 331140 38690 331168 48175
rect 330208 38684 330260 38690
rect 330208 38626 330260 38632
rect 331128 38684 331180 38690
rect 331128 38626 331180 38632
rect 330220 26314 330248 38626
rect 330208 26308 330260 26314
rect 330208 26250 330260 26256
rect 330208 9716 330260 9722
rect 330208 9658 330260 9664
rect 330024 9104 330076 9110
rect 330024 9046 330076 9052
rect 330220 7818 330248 9658
rect 330208 7812 330260 7818
rect 330208 7754 330260 7760
rect 331232 5166 331260 335582
rect 331324 7886 331352 335650
rect 331416 331906 331444 340068
rect 331600 340054 331890 340082
rect 331968 340054 332350 340082
rect 332796 340054 332902 340082
rect 333072 340054 333362 340082
rect 333440 340054 333822 340082
rect 334176 340054 334374 340082
rect 334544 340054 334834 340082
rect 334912 340054 335294 340082
rect 335464 340054 335846 340082
rect 336016 340054 336306 340082
rect 331600 335646 331628 340054
rect 331968 335714 331996 340054
rect 331956 335708 332008 335714
rect 331956 335650 332008 335656
rect 331588 335640 331640 335646
rect 331588 335582 331640 335588
rect 332600 335640 332652 335646
rect 332600 335582 332652 335588
rect 331404 331900 331456 331906
rect 331404 331842 331456 331848
rect 331404 318912 331456 318918
rect 331404 318854 331456 318860
rect 331416 317422 331444 318854
rect 331404 317416 331456 317422
rect 331404 317358 331456 317364
rect 331404 299600 331456 299606
rect 331404 299542 331456 299548
rect 331416 288454 331444 299542
rect 331404 288448 331456 288454
rect 331404 288390 331456 288396
rect 331496 288448 331548 288454
rect 331496 288390 331548 288396
rect 331508 278866 331536 288390
rect 331496 278860 331548 278866
rect 331496 278802 331548 278808
rect 331404 278724 331456 278730
rect 331404 278666 331456 278672
rect 331416 277370 331444 278666
rect 331404 277364 331456 277370
rect 331404 277306 331456 277312
rect 331404 267776 331456 267782
rect 331404 267718 331456 267724
rect 331416 259418 331444 267718
rect 331404 259412 331456 259418
rect 331404 259354 331456 259360
rect 331404 236700 331456 236706
rect 331404 236642 331456 236648
rect 331416 222222 331444 236642
rect 331404 222216 331456 222222
rect 331404 222158 331456 222164
rect 331416 220862 331444 220893
rect 331404 220856 331456 220862
rect 331456 220804 331536 220810
rect 331404 220798 331536 220804
rect 331416 220782 331536 220798
rect 331508 211154 331536 220782
rect 331416 211126 331536 211154
rect 331416 203046 331444 211126
rect 331404 203040 331456 203046
rect 331404 202982 331456 202988
rect 331404 202904 331456 202910
rect 331404 202846 331456 202852
rect 331416 200122 331444 202846
rect 331404 200116 331456 200122
rect 331404 200058 331456 200064
rect 331588 191820 331640 191826
rect 331588 191762 331640 191768
rect 331600 190482 331628 191762
rect 331600 190466 331720 190482
rect 331404 190460 331456 190466
rect 331600 190460 331732 190466
rect 331600 190454 331680 190460
rect 331404 190402 331456 190408
rect 331680 190402 331732 190408
rect 331416 180849 331444 190402
rect 331692 190371 331720 190402
rect 331402 180840 331458 180849
rect 331402 180775 331458 180784
rect 331586 180840 331642 180849
rect 331586 180775 331642 180784
rect 331600 172582 331628 180775
rect 331588 172576 331640 172582
rect 331588 172518 331640 172524
rect 331588 172440 331640 172446
rect 331588 172382 331640 172388
rect 331600 171086 331628 172382
rect 331588 171080 331640 171086
rect 331588 171022 331640 171028
rect 331680 161492 331732 161498
rect 331680 161434 331732 161440
rect 331692 151881 331720 161434
rect 331494 151872 331550 151881
rect 331416 151830 331494 151858
rect 331416 146062 331444 151830
rect 331494 151807 331550 151816
rect 331678 151872 331734 151881
rect 331678 151807 331734 151816
rect 331404 146056 331456 146062
rect 331404 145998 331456 146004
rect 331404 133952 331456 133958
rect 331404 133894 331456 133900
rect 331416 125594 331444 133894
rect 331404 125588 331456 125594
rect 331404 125530 331456 125536
rect 331588 125588 331640 125594
rect 331588 125530 331640 125536
rect 331600 118402 331628 125530
rect 331508 118374 331628 118402
rect 331508 104938 331536 118374
rect 331416 104910 331536 104938
rect 331416 103494 331444 104910
rect 331404 103488 331456 103494
rect 331404 103430 331456 103436
rect 331404 93900 331456 93906
rect 331404 93842 331456 93848
rect 331416 85610 331444 93842
rect 331862 87408 331918 87417
rect 331862 87343 331918 87352
rect 331876 87145 331904 87343
rect 331862 87136 331918 87145
rect 331862 87071 331918 87080
rect 331404 85604 331456 85610
rect 331404 85546 331456 85552
rect 331680 85604 331732 85610
rect 331680 85546 331732 85552
rect 331692 75954 331720 85546
rect 331404 75948 331456 75954
rect 331404 75890 331456 75896
rect 331680 75948 331732 75954
rect 331680 75890 331732 75896
rect 331416 66201 331444 75890
rect 331402 66192 331458 66201
rect 331402 66127 331458 66136
rect 331586 66056 331642 66065
rect 331586 65991 331642 66000
rect 331600 48385 331628 65991
rect 331586 48376 331642 48385
rect 331586 48311 331642 48320
rect 331496 38684 331548 38690
rect 331496 38626 331548 38632
rect 331508 27849 331536 38626
rect 331494 27840 331550 27849
rect 331494 27775 331550 27784
rect 331402 27704 331458 27713
rect 331402 27639 331458 27648
rect 331416 26246 331444 27639
rect 331404 26240 331456 26246
rect 331404 26182 331456 26188
rect 331404 9716 331456 9722
rect 331404 9658 331456 9664
rect 331416 8362 331444 9658
rect 331404 8356 331456 8362
rect 331404 8298 331456 8304
rect 331312 7880 331364 7886
rect 331312 7822 331364 7828
rect 332612 5234 332640 335582
rect 332692 335096 332744 335102
rect 332692 335038 332744 335044
rect 332704 7954 332732 335038
rect 332796 9178 332824 340054
rect 333072 335646 333100 340054
rect 333244 337204 333296 337210
rect 333244 337146 333296 337152
rect 333060 335640 333112 335646
rect 333060 335582 333112 335588
rect 332784 9172 332836 9178
rect 332784 9114 332836 9120
rect 332692 7948 332744 7954
rect 332692 7890 332744 7896
rect 332600 5228 332652 5234
rect 332600 5170 332652 5176
rect 331220 5160 331272 5166
rect 331220 5102 331272 5108
rect 329840 5092 329892 5098
rect 329840 5034 329892 5040
rect 328736 5024 328788 5030
rect 328736 4966 328788 4972
rect 328460 4820 328512 4826
rect 328460 4762 328512 4768
rect 328472 3738 328500 4762
rect 333256 4146 333284 337146
rect 333440 335102 333468 340054
rect 334072 335708 334124 335714
rect 334072 335650 334124 335656
rect 333980 335640 334032 335646
rect 333980 335582 334032 335588
rect 333428 335096 333480 335102
rect 333428 335038 333480 335044
rect 333612 5024 333664 5030
rect 333612 4966 333664 4972
rect 332416 4140 332468 4146
rect 332416 4082 332468 4088
rect 333244 4140 333296 4146
rect 333244 4082 333296 4088
rect 328460 3732 328512 3738
rect 328460 3674 328512 3680
rect 331220 3732 331272 3738
rect 331220 3674 331272 3680
rect 327724 3120 327776 3126
rect 327724 3062 327776 3068
rect 328828 3120 328880 3126
rect 328828 3062 328880 3068
rect 327632 3052 327684 3058
rect 327632 2994 327684 3000
rect 327644 480 327672 2994
rect 328840 480 328868 3062
rect 330024 2848 330076 2854
rect 330024 2790 330076 2796
rect 330036 480 330064 2790
rect 331232 480 331260 3674
rect 332428 480 332456 4082
rect 333624 480 333652 4966
rect 333992 4690 334020 335582
rect 334084 8022 334112 335650
rect 334176 9246 334204 340054
rect 334544 335646 334572 340054
rect 334912 335714 334940 340054
rect 335268 337068 335320 337074
rect 335268 337010 335320 337016
rect 334900 335708 334952 335714
rect 334900 335650 334952 335656
rect 334532 335640 334584 335646
rect 334532 335582 334584 335588
rect 335174 110800 335230 110809
rect 335174 110735 335230 110744
rect 335188 110673 335216 110735
rect 335174 110664 335230 110673
rect 335174 110599 335230 110608
rect 334164 9240 334216 9246
rect 334164 9182 334216 9188
rect 334072 8016 334124 8022
rect 334072 7958 334124 7964
rect 333980 4684 334032 4690
rect 333980 4626 334032 4632
rect 335280 4146 335308 337010
rect 335360 333940 335412 333946
rect 335360 333882 335412 333888
rect 335372 4554 335400 333882
rect 335464 6662 335492 340054
rect 336016 333946 336044 340054
rect 336096 337884 336148 337890
rect 336096 337826 336148 337832
rect 336004 333940 336056 333946
rect 336004 333882 336056 333888
rect 336108 333010 336136 337826
rect 336186 337784 336242 337793
rect 336186 337719 336188 337728
rect 336240 337719 336242 337728
rect 336188 337690 336240 337696
rect 336016 332982 336136 333010
rect 335452 6656 335504 6662
rect 335452 6598 335504 6604
rect 335360 4548 335412 4554
rect 335360 4490 335412 4496
rect 334716 4140 334768 4146
rect 334716 4082 334768 4088
rect 335268 4140 335320 4146
rect 335268 4082 335320 4088
rect 334728 480 334756 4082
rect 335544 3800 335596 3806
rect 336016 3754 336044 332982
rect 336752 331906 336780 340068
rect 337028 340054 337318 340082
rect 336740 331900 336792 331906
rect 336740 331842 336792 331848
rect 336924 331900 336976 331906
rect 336924 331842 336976 331848
rect 336832 327140 336884 327146
rect 336832 327082 336884 327088
rect 336738 157584 336794 157593
rect 336738 157519 336740 157528
rect 336792 157519 336794 157528
rect 336740 157490 336792 157496
rect 336738 87136 336794 87145
rect 336738 87071 336740 87080
rect 336792 87071 336794 87080
rect 336740 87042 336792 87048
rect 336646 29336 336702 29345
rect 336646 29271 336702 29280
rect 336660 29073 336688 29271
rect 336646 29064 336702 29073
rect 336646 28999 336702 29008
rect 336646 17096 336702 17105
rect 336646 17031 336702 17040
rect 336660 16697 336688 17031
rect 336646 16688 336702 16697
rect 336646 16623 336702 16632
rect 336844 6730 336872 327082
rect 336936 8090 336964 331842
rect 337028 327214 337056 340054
rect 337396 335594 337424 340190
rect 338238 340054 338344 340082
rect 337120 335566 337424 335594
rect 338120 335640 338172 335646
rect 338120 335582 338172 335588
rect 337120 331208 337148 335566
rect 337120 331180 337240 331208
rect 337016 327208 337068 327214
rect 337016 327150 337068 327156
rect 337212 319025 337240 331180
rect 337198 319016 337254 319025
rect 337198 318951 337254 318960
rect 337106 318880 337162 318889
rect 337106 318815 337162 318824
rect 337120 311982 337148 318815
rect 337108 311976 337160 311982
rect 337108 311918 337160 311924
rect 337200 309120 337252 309126
rect 337200 309062 337252 309068
rect 337212 307850 337240 309062
rect 337120 307822 337240 307850
rect 337120 307766 337148 307822
rect 337108 307760 337160 307766
rect 337108 307702 337160 307708
rect 337292 298172 337344 298178
rect 337292 298114 337344 298120
rect 337304 290426 337332 298114
rect 337108 290420 337160 290426
rect 337108 290362 337160 290368
rect 337292 290420 337344 290426
rect 337292 290362 337344 290368
rect 337120 288386 337148 290362
rect 337108 288380 337160 288386
rect 337108 288322 337160 288328
rect 337200 278792 337252 278798
rect 337200 278734 337252 278740
rect 337212 273358 337240 278734
rect 337200 273352 337252 273358
rect 337200 273294 337252 273300
rect 337108 273216 337160 273222
rect 337108 273158 337160 273164
rect 337120 269113 337148 273158
rect 337106 269104 337162 269113
rect 337106 269039 337162 269048
rect 337290 269104 337346 269113
rect 337290 269039 337346 269048
rect 337304 259486 337332 269039
rect 337108 259480 337160 259486
rect 337108 259422 337160 259428
rect 337292 259480 337344 259486
rect 337292 259422 337344 259428
rect 337120 253978 337148 259422
rect 337108 253972 337160 253978
rect 337108 253914 337160 253920
rect 337292 253836 337344 253842
rect 337292 253778 337344 253784
rect 337304 240145 337332 253778
rect 337106 240136 337162 240145
rect 337106 240071 337162 240080
rect 337290 240136 337346 240145
rect 337290 240071 337346 240080
rect 337120 231554 337148 240071
rect 337120 231526 337332 231554
rect 337304 225350 337332 231526
rect 337292 225344 337344 225350
rect 337292 225286 337344 225292
rect 337292 222216 337344 222222
rect 337292 222158 337344 222164
rect 337304 220833 337332 222158
rect 337106 220824 337162 220833
rect 337106 220759 337162 220768
rect 337290 220824 337346 220833
rect 337290 220759 337346 220768
rect 337120 212242 337148 220759
rect 337120 212214 337332 212242
rect 337304 202910 337332 212214
rect 337200 202904 337252 202910
rect 337200 202846 337252 202852
rect 337292 202904 337344 202910
rect 337292 202846 337344 202852
rect 337212 196110 337240 202846
rect 337200 196104 337252 196110
rect 337200 196046 337252 196052
rect 337108 195968 337160 195974
rect 337108 195910 337160 195916
rect 337120 191826 337148 195910
rect 337108 191820 337160 191826
rect 337108 191762 337160 191768
rect 337108 186312 337160 186318
rect 337108 186254 337160 186260
rect 337120 172582 337148 186254
rect 337108 172576 337160 172582
rect 337108 172518 337160 172524
rect 337108 172440 337160 172446
rect 337108 172382 337160 172388
rect 337120 171086 337148 172382
rect 337108 171080 337160 171086
rect 337108 171022 337160 171028
rect 337292 161492 337344 161498
rect 337292 161434 337344 161440
rect 337304 153270 337332 161434
rect 337292 153264 337344 153270
rect 337292 153206 337344 153212
rect 337200 153196 337252 153202
rect 337200 153138 337252 153144
rect 337212 135425 337240 153138
rect 337198 135416 337254 135425
rect 337198 135351 337254 135360
rect 337198 135280 337254 135289
rect 337108 135244 337160 135250
rect 337198 135215 337200 135224
rect 337108 135186 337160 135192
rect 337252 135215 337254 135224
rect 337200 135186 337252 135192
rect 337120 125594 337148 135186
rect 337108 125588 337160 125594
rect 337108 125530 337160 125536
rect 337292 125588 337344 125594
rect 337292 125530 337344 125536
rect 337304 120578 337332 125530
rect 337212 120550 337332 120578
rect 337212 114510 337240 120550
rect 337200 114504 337252 114510
rect 337200 114446 337252 114452
rect 337016 104916 337068 104922
rect 337016 104858 337068 104864
rect 337028 104786 337056 104858
rect 337016 104780 337068 104786
rect 337016 104722 337068 104728
rect 337200 95260 337252 95266
rect 337200 95202 337252 95208
rect 337212 80458 337240 95202
rect 337212 80430 337332 80458
rect 337304 80186 337332 80430
rect 337212 80158 337332 80186
rect 337212 60858 337240 80158
rect 337200 60852 337252 60858
rect 337200 60794 337252 60800
rect 337200 60648 337252 60654
rect 337200 60590 337252 60596
rect 337212 51134 337240 60590
rect 337200 51128 337252 51134
rect 337200 51070 337252 51076
rect 337108 48340 337160 48346
rect 337108 48282 337160 48288
rect 337120 43466 337148 48282
rect 337120 43438 337240 43466
rect 337212 22114 337240 43438
rect 337120 22086 337240 22114
rect 337120 14498 337148 22086
rect 337120 14470 337240 14498
rect 336924 8084 336976 8090
rect 336924 8026 336976 8032
rect 336832 6724 336884 6730
rect 336832 6666 336884 6672
rect 337108 5092 337160 5098
rect 337108 5034 337160 5040
rect 335596 3748 336044 3754
rect 335544 3742 336044 3748
rect 335556 3726 336044 3742
rect 335556 3194 335952 3210
rect 335556 3188 335964 3194
rect 335556 3182 335912 3188
rect 335556 2854 335584 3182
rect 335912 3130 335964 3136
rect 335912 3052 335964 3058
rect 335912 2994 335964 3000
rect 335544 2848 335596 2854
rect 335544 2790 335596 2796
rect 335924 480 335952 2994
rect 337120 480 337148 5034
rect 337212 4622 337240 14470
rect 337200 4616 337252 4622
rect 337200 4558 337252 4564
rect 338132 4486 338160 335582
rect 338316 8158 338344 340054
rect 338408 340054 338790 340082
rect 338960 340054 339250 340082
rect 339604 340054 339710 340082
rect 338304 8152 338356 8158
rect 338304 8094 338356 8100
rect 338408 6594 338436 340054
rect 338764 337476 338816 337482
rect 338764 337418 338816 337424
rect 338396 6588 338448 6594
rect 338396 6530 338448 6536
rect 338120 4480 338172 4486
rect 338120 4422 338172 4428
rect 338776 4146 338804 337418
rect 338960 335646 338988 340054
rect 338948 335640 339000 335646
rect 338948 335582 339000 335588
rect 339604 8226 339632 340054
rect 340248 337414 340276 340068
rect 340236 337408 340288 337414
rect 340236 337350 340288 337356
rect 340340 328506 340368 340190
rect 340984 340054 341182 340082
rect 340788 337408 340840 337414
rect 340788 337350 340840 337356
rect 339776 328500 339828 328506
rect 339776 328442 339828 328448
rect 340328 328500 340380 328506
rect 340328 328442 340380 328448
rect 339788 311930 339816 328442
rect 339696 311902 339816 311930
rect 339696 311794 339724 311902
rect 339696 311766 339816 311794
rect 339788 282962 339816 311766
rect 339696 282934 339816 282962
rect 339696 282826 339724 282934
rect 339696 282798 339816 282826
rect 339788 263650 339816 282798
rect 339696 263622 339816 263650
rect 339696 263514 339724 263622
rect 339696 263486 339816 263514
rect 339788 244338 339816 263486
rect 339696 244310 339816 244338
rect 339696 244202 339724 244310
rect 339696 244174 339816 244202
rect 339788 225026 339816 244174
rect 339696 224998 339816 225026
rect 339696 224890 339724 224998
rect 339696 224862 339816 224890
rect 339788 205714 339816 224862
rect 339696 205686 339816 205714
rect 339696 205578 339724 205686
rect 339696 205550 339816 205578
rect 339788 186998 339816 205550
rect 339776 186992 339828 186998
rect 339776 186934 339828 186940
rect 339960 186992 340012 186998
rect 339960 186934 340012 186940
rect 339972 182209 340000 186934
rect 339774 182200 339830 182209
rect 339774 182135 339830 182144
rect 339958 182200 340014 182209
rect 339958 182135 340014 182144
rect 339788 172530 339816 182135
rect 339696 172502 339816 172530
rect 339696 169130 339724 172502
rect 339696 169102 339908 169130
rect 339880 157298 339908 169102
rect 339788 157270 339908 157298
rect 339788 138122 339816 157270
rect 339696 138094 339816 138122
rect 339696 137986 339724 138094
rect 339696 137958 339816 137986
rect 339788 135250 339816 137958
rect 339776 135244 339828 135250
rect 339776 135186 339828 135192
rect 339684 124296 339736 124302
rect 339736 124244 339816 124250
rect 339684 124238 339816 124244
rect 339696 124222 339816 124238
rect 339788 122806 339816 124222
rect 339776 122800 339828 122806
rect 339776 122742 339828 122748
rect 339776 118040 339828 118046
rect 339776 117982 339828 117988
rect 339788 80170 339816 117982
rect 339776 80164 339828 80170
rect 339776 80106 339828 80112
rect 339776 80028 339828 80034
rect 339776 79970 339828 79976
rect 339788 60858 339816 79970
rect 339776 60852 339828 60858
rect 339776 60794 339828 60800
rect 339776 56636 339828 56642
rect 339776 56578 339828 56584
rect 339788 46918 339816 56578
rect 339776 46912 339828 46918
rect 339776 46854 339828 46860
rect 339776 42084 339828 42090
rect 339776 42026 339828 42032
rect 339788 31822 339816 42026
rect 339776 31816 339828 31822
rect 339776 31758 339828 31764
rect 339684 29028 339736 29034
rect 339684 28970 339736 28976
rect 339696 19378 339724 28970
rect 339684 19372 339736 19378
rect 339684 19314 339736 19320
rect 339776 19372 339828 19378
rect 339776 19314 339828 19320
rect 339788 19242 339816 19314
rect 339776 19236 339828 19242
rect 339776 19178 339828 19184
rect 339684 9716 339736 9722
rect 339684 9658 339736 9664
rect 339592 8220 339644 8226
rect 339592 8162 339644 8168
rect 339696 6526 339724 9658
rect 339684 6520 339736 6526
rect 339684 6462 339736 6468
rect 340800 4146 340828 337350
rect 340880 164212 340932 164218
rect 340880 164154 340932 164160
rect 340892 154601 340920 164154
rect 340878 154592 340934 154601
rect 340878 154527 340934 154536
rect 340984 8294 341012 340054
rect 341628 338842 341656 340068
rect 341720 340054 342194 340082
rect 342364 340054 342654 340082
rect 341616 338836 341668 338842
rect 341616 338778 341668 338784
rect 341720 331362 341748 340054
rect 341892 337136 341944 337142
rect 341892 337078 341944 337084
rect 341432 331356 341484 331362
rect 341432 331298 341484 331304
rect 341708 331356 341760 331362
rect 341708 331298 341760 331304
rect 341444 328522 341472 331298
rect 341904 331242 341932 337078
rect 341352 328494 341472 328522
rect 341536 331214 341932 331242
rect 341352 328438 341380 328494
rect 341340 328432 341392 328438
rect 341340 328374 341392 328380
rect 341432 318844 341484 318850
rect 341432 318786 341484 318792
rect 341444 311914 341472 318786
rect 341248 311908 341300 311914
rect 341248 311850 341300 311856
rect 341432 311908 341484 311914
rect 341432 311850 341484 311856
rect 341260 309126 341288 311850
rect 341248 309120 341300 309126
rect 341248 309062 341300 309068
rect 341156 299532 341208 299538
rect 341156 299474 341208 299480
rect 341168 299418 341196 299474
rect 341246 299432 341302 299441
rect 341168 299390 341246 299418
rect 341246 299367 341302 299376
rect 341246 289912 341302 289921
rect 341246 289847 341302 289856
rect 341260 289814 341288 289847
rect 341248 289808 341300 289814
rect 341248 289750 341300 289756
rect 341156 280220 341208 280226
rect 341156 280162 341208 280168
rect 341168 280106 341196 280162
rect 341246 280120 341302 280129
rect 341168 280078 341246 280106
rect 341246 280055 341302 280064
rect 341246 270600 341302 270609
rect 341246 270535 341302 270544
rect 341260 270502 341288 270535
rect 341248 270496 341300 270502
rect 341248 270438 341300 270444
rect 341156 260908 341208 260914
rect 341156 260850 341208 260856
rect 341168 260794 341196 260850
rect 341246 260808 341302 260817
rect 341168 260766 341246 260794
rect 341246 260743 341302 260752
rect 341246 251288 341302 251297
rect 341246 251223 341302 251232
rect 341260 244390 341288 251223
rect 341248 244384 341300 244390
rect 341248 244326 341300 244332
rect 341156 244248 341208 244254
rect 341156 244190 341208 244196
rect 341168 240145 341196 244190
rect 341154 240136 341210 240145
rect 341154 240071 341210 240080
rect 341430 240136 341486 240145
rect 341430 240071 341486 240080
rect 341444 230518 341472 240071
rect 341248 230512 341300 230518
rect 341248 230454 341300 230460
rect 341432 230512 341484 230518
rect 341432 230454 341484 230460
rect 341260 225078 341288 230454
rect 341248 225072 341300 225078
rect 341248 225014 341300 225020
rect 341156 224936 341208 224942
rect 341156 224878 341208 224884
rect 341168 220794 341196 224878
rect 341156 220788 341208 220794
rect 341156 220730 341208 220736
rect 341156 215280 341208 215286
rect 341156 215222 341208 215228
rect 341168 211154 341196 215222
rect 341168 211126 341288 211154
rect 341260 202910 341288 211126
rect 341156 202904 341208 202910
rect 341154 202872 341156 202881
rect 341248 202904 341300 202910
rect 341208 202872 341210 202881
rect 341248 202846 341300 202852
rect 341430 202872 341486 202881
rect 341154 202807 341210 202816
rect 341430 202807 341486 202816
rect 341444 193254 341472 202807
rect 341248 193248 341300 193254
rect 341248 193190 341300 193196
rect 341432 193248 341484 193254
rect 341432 193190 341484 193196
rect 341260 186266 341288 193190
rect 341168 186238 341288 186266
rect 341168 182170 341196 186238
rect 341156 182164 341208 182170
rect 341156 182106 341208 182112
rect 341248 182164 341300 182170
rect 341248 182106 341300 182112
rect 341260 164966 341288 182106
rect 341064 164960 341116 164966
rect 341064 164902 341116 164908
rect 341248 164960 341300 164966
rect 341248 164902 341300 164908
rect 341076 164218 341104 164902
rect 341064 164212 341116 164218
rect 341064 164154 341116 164160
rect 341338 154592 341394 154601
rect 341338 154527 341394 154536
rect 341352 147642 341380 154527
rect 341260 147614 341380 147642
rect 341260 138718 341288 147614
rect 341248 138712 341300 138718
rect 341248 138654 341300 138660
rect 341340 128308 341392 128314
rect 341340 128250 341392 128256
rect 341352 125610 341380 128250
rect 341352 125582 341472 125610
rect 341444 118726 341472 125582
rect 341248 118720 341300 118726
rect 341248 118662 341300 118668
rect 341432 118720 341484 118726
rect 341432 118662 341484 118668
rect 341260 115938 341288 118662
rect 341248 115932 341300 115938
rect 341248 115874 341300 115880
rect 341156 106344 341208 106350
rect 341156 106286 341208 106292
rect 341168 99414 341196 106286
rect 341156 99408 341208 99414
rect 341156 99350 341208 99356
rect 341248 99340 341300 99346
rect 341248 99282 341300 99288
rect 341260 89706 341288 99282
rect 341168 89678 341288 89706
rect 341168 86970 341196 89678
rect 341156 86964 341208 86970
rect 341156 86906 341208 86912
rect 341064 77308 341116 77314
rect 341064 77250 341116 77256
rect 341076 77178 341104 77250
rect 341064 77172 341116 77178
rect 341064 77114 341116 77120
rect 341156 70304 341208 70310
rect 341156 70246 341208 70252
rect 341168 61554 341196 70246
rect 341168 61526 341472 61554
rect 341444 56658 341472 61526
rect 341352 56630 341472 56658
rect 341352 56574 341380 56630
rect 341340 56568 341392 56574
rect 341340 56510 341392 56516
rect 341340 50652 341392 50658
rect 341340 50594 341392 50600
rect 341352 38570 341380 50594
rect 341168 38542 341380 38570
rect 341168 31822 341196 38542
rect 341156 31816 341208 31822
rect 341156 31758 341208 31764
rect 341156 31680 341208 31686
rect 341156 31622 341208 31628
rect 341168 28937 341196 31622
rect 341154 28928 341210 28937
rect 341154 28863 341210 28872
rect 341338 28928 341394 28937
rect 341338 28863 341394 28872
rect 341352 19378 341380 28863
rect 341248 19372 341300 19378
rect 341248 19314 341300 19320
rect 341340 19372 341392 19378
rect 341340 19314 341392 19320
rect 340972 8288 341024 8294
rect 340972 8230 341024 8236
rect 341260 6458 341288 19314
rect 341248 6452 341300 6458
rect 341248 6394 341300 6400
rect 338764 4140 338816 4146
rect 338764 4082 338816 4088
rect 339500 4140 339552 4146
rect 339500 4082 339552 4088
rect 340788 4140 340840 4146
rect 340788 4082 340840 4088
rect 338304 3732 338356 3738
rect 338304 3674 338356 3680
rect 338316 480 338344 3674
rect 339512 480 339540 4082
rect 341536 3806 341564 331214
rect 342364 6186 342392 340054
rect 342904 337544 342956 337550
rect 342904 337486 342956 337492
rect 342352 6180 342404 6186
rect 342352 6122 342404 6128
rect 342916 3874 342944 337486
rect 343100 336870 343128 340068
rect 343088 336864 343140 336870
rect 343088 336806 343140 336812
rect 343652 6390 343680 340068
rect 344112 336802 344140 340068
rect 344572 337890 344600 340068
rect 345138 340054 345244 340082
rect 344560 337884 344612 337890
rect 344560 337826 344612 337832
rect 344284 336864 344336 336870
rect 344284 336806 344336 336812
rect 344100 336796 344152 336802
rect 344100 336738 344152 336744
rect 343640 6384 343692 6390
rect 343640 6326 343692 6332
rect 342904 3868 342956 3874
rect 342904 3810 342956 3816
rect 343088 3868 343140 3874
rect 343088 3810 343140 3816
rect 341524 3800 341576 3806
rect 341524 3742 341576 3748
rect 341892 3800 341944 3806
rect 341892 3742 341944 3748
rect 340696 3188 340748 3194
rect 340696 3130 340748 3136
rect 340708 480 340736 3130
rect 340878 3088 340934 3097
rect 340878 3023 340934 3032
rect 340892 2922 340920 3023
rect 340880 2916 340932 2922
rect 340880 2858 340932 2864
rect 341904 480 341932 3742
rect 343100 480 343128 3810
rect 344296 3074 344324 336806
rect 344376 336796 344428 336802
rect 344376 336738 344428 336744
rect 344388 3330 344416 336738
rect 345216 6254 345244 340054
rect 345308 340054 345598 340082
rect 345676 340054 346058 340082
rect 345308 337618 345336 340054
rect 345296 337612 345348 337618
rect 345296 337554 345348 337560
rect 345676 337090 345704 340054
rect 345492 337062 345704 337090
rect 345492 336938 345520 337062
rect 345480 336932 345532 336938
rect 345480 336874 345532 336880
rect 345664 336932 345716 336938
rect 345664 336874 345716 336880
rect 345204 6248 345256 6254
rect 345204 6190 345256 6196
rect 345676 4146 345704 336874
rect 346308 157548 346360 157554
rect 346308 157490 346360 157496
rect 346320 157457 346348 157490
rect 346306 157448 346362 157457
rect 346306 157383 346362 157392
rect 346308 87100 346360 87106
rect 346308 87042 346360 87048
rect 346320 87009 346348 87042
rect 346306 87000 346362 87009
rect 346306 86935 346362 86944
rect 346596 5302 346624 340068
rect 347056 337686 347084 340068
rect 347044 337680 347096 337686
rect 347044 337622 347096 337628
rect 347516 337482 347544 340068
rect 347976 340054 348082 340082
rect 347504 337476 347556 337482
rect 347504 337418 347556 337424
rect 347976 5370 348004 340054
rect 348528 338706 348556 340068
rect 348516 338700 348568 338706
rect 348516 338642 348568 338648
rect 348424 337680 348476 337686
rect 348424 337622 348476 337628
rect 347964 5364 348016 5370
rect 347964 5306 348016 5312
rect 346584 5296 346636 5302
rect 346584 5238 346636 5244
rect 345664 4140 345716 4146
rect 345664 4082 345716 4088
rect 347872 4140 347924 4146
rect 347872 4082 347924 4088
rect 344376 3324 344428 3330
rect 344376 3266 344428 3272
rect 345756 3324 345808 3330
rect 345756 3266 345808 3272
rect 345768 3097 345796 3266
rect 346676 3188 346728 3194
rect 346676 3130 346728 3136
rect 345754 3088 345810 3097
rect 344296 3046 344416 3074
rect 344388 2990 344416 3046
rect 345754 3023 345810 3032
rect 344376 2984 344428 2990
rect 344376 2926 344428 2932
rect 345480 2984 345532 2990
rect 345480 2926 345532 2932
rect 344284 2916 344336 2922
rect 344284 2858 344336 2864
rect 344296 480 344324 2858
rect 345492 480 345520 2926
rect 346688 480 346716 3130
rect 347884 480 347912 4082
rect 348436 3330 348464 337622
rect 348988 337142 349016 340068
rect 349356 340054 349554 340082
rect 349068 337476 349120 337482
rect 349068 337418 349120 337424
rect 348976 337136 349028 337142
rect 348976 337078 349028 337084
rect 349080 4146 349108 337418
rect 349356 5438 349384 340054
rect 350000 337890 350028 340068
rect 349988 337884 350040 337890
rect 349988 337826 350040 337832
rect 350460 337278 350488 340068
rect 350644 340054 351026 340082
rect 350448 337272 350500 337278
rect 350448 337214 350500 337220
rect 350644 6322 350672 340054
rect 351472 337618 351500 340068
rect 351932 337822 351960 340068
rect 352116 340054 352498 340082
rect 351920 337816 351972 337822
rect 351920 337758 351972 337764
rect 351460 337612 351512 337618
rect 351460 337554 351512 337560
rect 351644 337612 351696 337618
rect 351644 337554 351696 337560
rect 351656 336870 351684 337554
rect 351828 337136 351880 337142
rect 351828 337078 351880 337084
rect 351184 336864 351236 336870
rect 351184 336806 351236 336812
rect 351644 336864 351696 336870
rect 351644 336806 351696 336812
rect 350632 6316 350684 6322
rect 350632 6258 350684 6264
rect 349344 5432 349396 5438
rect 349344 5374 349396 5380
rect 351196 4146 351224 336806
rect 351840 4146 351868 337078
rect 352116 5506 352144 340054
rect 352944 337958 352972 340068
rect 352932 337952 352984 337958
rect 352932 337894 352984 337900
rect 353404 337550 353432 340068
rect 353496 340054 353970 340082
rect 353392 337544 353444 337550
rect 353392 337486 353444 337492
rect 352564 336796 352616 336802
rect 352564 336738 352616 336744
rect 352104 5500 352156 5506
rect 352104 5442 352156 5448
rect 352576 4486 352604 336738
rect 353496 4554 353524 340054
rect 354416 338094 354444 340068
rect 354404 338088 354456 338094
rect 354404 338030 354456 338036
rect 354876 336870 354904 340068
rect 354968 340054 355442 340082
rect 354864 336864 354916 336870
rect 354864 336806 354916 336812
rect 353484 4548 353536 4554
rect 353484 4490 353536 4496
rect 352564 4480 352616 4486
rect 352564 4422 352616 4428
rect 354968 4350 354996 340054
rect 355888 338026 355916 340068
rect 356256 340054 356362 340082
rect 356624 340054 356914 340082
rect 355876 338020 355928 338026
rect 355876 337962 355928 337968
rect 355324 337952 355376 337958
rect 355324 337894 355376 337900
rect 354956 4344 355008 4350
rect 354956 4286 355008 4292
rect 349068 4140 349120 4146
rect 349068 4082 349120 4088
rect 351184 4140 351236 4146
rect 351184 4082 351236 4088
rect 351368 4140 351420 4146
rect 351368 4082 351420 4088
rect 351828 4140 351880 4146
rect 351828 4082 351880 4088
rect 348424 3324 348476 3330
rect 348424 3266 348476 3272
rect 349068 3324 349120 3330
rect 349068 3266 349120 3272
rect 349080 480 349108 3266
rect 350264 3256 350316 3262
rect 350264 3198 350316 3204
rect 350276 480 350304 3198
rect 351380 480 351408 4082
rect 355336 4010 355364 337894
rect 355968 337272 356020 337278
rect 355968 337214 356020 337220
rect 355324 4004 355376 4010
rect 355324 3946 355376 3952
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 352564 3256 352616 3262
rect 352564 3198 352616 3204
rect 352576 480 352604 3198
rect 353772 480 353800 3334
rect 355980 2990 356008 337214
rect 356152 335640 356204 335646
rect 356152 335582 356204 335588
rect 356164 4282 356192 335582
rect 356152 4276 356204 4282
rect 356152 4218 356204 4224
rect 356256 3369 356284 340054
rect 356624 335646 356652 340054
rect 356704 337680 356756 337686
rect 356704 337622 356756 337628
rect 356612 335640 356664 335646
rect 356612 335582 356664 335588
rect 356242 3360 356298 3369
rect 356242 3295 356298 3304
rect 354956 2984 355008 2990
rect 354956 2926 355008 2932
rect 355968 2984 356020 2990
rect 355968 2926 356020 2932
rect 354968 480 354996 2926
rect 356716 2854 356744 337622
rect 357360 337550 357388 340068
rect 357348 337544 357400 337550
rect 357348 337486 357400 337492
rect 357820 336802 357848 340068
rect 357808 336796 357860 336802
rect 357808 336738 357860 336744
rect 357912 335594 357940 340190
rect 358846 340054 358952 340082
rect 358084 338088 358136 338094
rect 358084 338030 358136 338036
rect 357728 335566 357940 335594
rect 357728 318850 357756 335566
rect 357624 318844 357676 318850
rect 357624 318786 357676 318792
rect 357716 318844 357768 318850
rect 357716 318786 357768 318792
rect 357636 311930 357664 318786
rect 357636 311902 357756 311930
rect 357728 302258 357756 311902
rect 357532 302252 357584 302258
rect 357532 302194 357584 302200
rect 357716 302252 357768 302258
rect 357716 302194 357768 302200
rect 357544 302138 357572 302194
rect 357544 302110 357664 302138
rect 357636 292618 357664 302110
rect 357636 292590 357756 292618
rect 357728 282946 357756 292590
rect 357532 282940 357584 282946
rect 357532 282882 357584 282888
rect 357716 282940 357768 282946
rect 357716 282882 357768 282888
rect 357544 282826 357572 282882
rect 357544 282798 357664 282826
rect 357636 273306 357664 282798
rect 357636 273278 357756 273306
rect 357728 263634 357756 273278
rect 357532 263628 357584 263634
rect 357532 263570 357584 263576
rect 357716 263628 357768 263634
rect 357716 263570 357768 263576
rect 357544 263514 357572 263570
rect 357544 263486 357664 263514
rect 357636 253994 357664 263486
rect 357636 253966 357756 253994
rect 357728 244322 357756 253966
rect 357532 244316 357584 244322
rect 357532 244258 357584 244264
rect 357716 244316 357768 244322
rect 357716 244258 357768 244264
rect 357544 244202 357572 244258
rect 357544 244174 357664 244202
rect 357636 234682 357664 244174
rect 357636 234654 357756 234682
rect 357728 225010 357756 234654
rect 357532 225004 357584 225010
rect 357532 224946 357584 224952
rect 357716 225004 357768 225010
rect 357716 224946 357768 224952
rect 357544 224890 357572 224946
rect 357544 224862 357664 224890
rect 357636 215370 357664 224862
rect 357636 215342 357756 215370
rect 357728 205698 357756 215342
rect 357532 205692 357584 205698
rect 357532 205634 357584 205640
rect 357716 205692 357768 205698
rect 357716 205634 357768 205640
rect 357544 205578 357572 205634
rect 357544 205550 357664 205578
rect 357636 196058 357664 205550
rect 357636 196030 357756 196058
rect 357728 186386 357756 196030
rect 357532 186380 357584 186386
rect 357532 186322 357584 186328
rect 357716 186380 357768 186386
rect 357716 186322 357768 186328
rect 357544 186266 357572 186322
rect 357544 186238 357664 186266
rect 357636 183569 357664 186238
rect 357438 183560 357494 183569
rect 357438 183495 357494 183504
rect 357622 183560 357678 183569
rect 357622 183495 357678 183504
rect 357452 173942 357480 183495
rect 357440 173936 357492 173942
rect 357440 173878 357492 173884
rect 357716 173936 357768 173942
rect 357716 173878 357768 173884
rect 357728 167074 357756 173878
rect 357532 167068 357584 167074
rect 357532 167010 357584 167016
rect 357716 167068 357768 167074
rect 357716 167010 357768 167016
rect 357544 166954 357572 167010
rect 357544 166926 357664 166954
rect 357636 157418 357664 166926
rect 357624 157412 357676 157418
rect 357624 157354 357676 157360
rect 357716 157276 357768 157282
rect 357716 157218 357768 157224
rect 357728 147694 357756 157218
rect 357532 147688 357584 147694
rect 357716 147688 357768 147694
rect 357584 147636 357664 147642
rect 357532 147630 357664 147636
rect 357716 147630 357768 147636
rect 357544 147614 357664 147630
rect 357636 144906 357664 147614
rect 357624 144900 357676 144906
rect 357624 144842 357676 144848
rect 357624 137964 357676 137970
rect 357624 137906 357676 137912
rect 357636 135266 357664 137906
rect 357636 135250 357756 135266
rect 357532 135244 357584 135250
rect 357636 135244 357768 135250
rect 357636 135238 357716 135244
rect 357532 135186 357584 135192
rect 357716 135186 357768 135192
rect 357544 133890 357572 135186
rect 357728 135155 357756 135186
rect 357532 133884 357584 133890
rect 357532 133826 357584 133832
rect 357624 124228 357676 124234
rect 357624 124170 357676 124176
rect 357636 124137 357664 124170
rect 357622 124128 357678 124137
rect 357622 124063 357678 124072
rect 357806 124128 357862 124137
rect 357806 124063 357862 124072
rect 357820 118674 357848 124063
rect 357728 118646 357848 118674
rect 357728 109750 357756 118646
rect 357716 109744 357768 109750
rect 357716 109686 357768 109692
rect 357624 99340 357676 99346
rect 357624 99282 357676 99288
rect 357636 96642 357664 99282
rect 357636 96614 357756 96642
rect 357728 89758 357756 96614
rect 357532 89752 357584 89758
rect 357716 89752 357768 89758
rect 357584 89700 357664 89706
rect 357532 89694 357664 89700
rect 357716 89694 357768 89700
rect 357544 89678 357664 89694
rect 357636 86970 357664 89678
rect 357624 86964 357676 86970
rect 357624 86906 357676 86912
rect 357716 77308 357768 77314
rect 357716 77250 357768 77256
rect 357728 67726 357756 77250
rect 357716 67720 357768 67726
rect 357716 67662 357768 67668
rect 357624 67652 357676 67658
rect 357624 67594 357676 67600
rect 357636 60738 357664 67594
rect 357636 60710 357756 60738
rect 357728 57934 357756 60710
rect 357716 57928 357768 57934
rect 357716 57870 357768 57876
rect 357624 48340 357676 48346
rect 357624 48282 357676 48288
rect 357636 41426 357664 48282
rect 357636 41398 357756 41426
rect 357728 29102 357756 41398
rect 357716 29096 357768 29102
rect 357716 29038 357768 29044
rect 357624 29028 357676 29034
rect 357624 28970 357676 28976
rect 357636 22114 357664 28970
rect 357636 22086 357756 22114
rect 357728 12458 357756 22086
rect 357544 12430 357756 12458
rect 357544 4214 357572 12430
rect 357532 4208 357584 4214
rect 357532 4150 357584 4156
rect 358096 3670 358124 338030
rect 358728 337816 358780 337822
rect 358728 337758 358780 337764
rect 358084 3664 358136 3670
rect 358084 3606 358136 3612
rect 357348 3256 357400 3262
rect 357348 3198 357400 3204
rect 356704 2848 356756 2854
rect 356704 2790 356756 2796
rect 356152 2712 356204 2718
rect 356152 2654 356204 2660
rect 356164 480 356192 2654
rect 357360 480 357388 3198
rect 358740 610 358768 337758
rect 358924 4146 358952 340054
rect 359108 340054 359306 340082
rect 359384 340054 359766 340082
rect 359004 335640 359056 335646
rect 359004 335582 359056 335588
rect 359016 4758 359044 335582
rect 359004 4752 359056 4758
rect 359004 4694 359056 4700
rect 358912 4140 358964 4146
rect 358912 4082 358964 4088
rect 359108 4010 359136 340054
rect 359384 335646 359412 340054
rect 359464 337544 359516 337550
rect 359464 337486 359516 337492
rect 359372 335640 359424 335646
rect 359372 335582 359424 335588
rect 359096 4004 359148 4010
rect 359096 3946 359148 3952
rect 359476 3126 359504 337486
rect 360304 336938 360332 340068
rect 360764 337686 360792 340068
rect 360948 340054 361238 340082
rect 360752 337680 360804 337686
rect 360752 337622 360804 337628
rect 360948 337498 360976 340054
rect 361672 337748 361724 337754
rect 361672 337690 361724 337696
rect 360396 337470 360976 337498
rect 360292 336932 360344 336938
rect 360292 336874 360344 336880
rect 360106 157584 360162 157593
rect 360290 157584 360346 157593
rect 360162 157542 360290 157570
rect 360106 157519 360162 157528
rect 360290 157519 360346 157528
rect 360106 134056 360162 134065
rect 360290 134056 360346 134065
rect 360162 134014 360290 134042
rect 360106 133991 360162 134000
rect 360290 133991 360346 134000
rect 360106 76120 360162 76129
rect 360290 76120 360346 76129
rect 360162 76078 360290 76106
rect 360106 76055 360162 76064
rect 360290 76055 360346 76064
rect 360106 63744 360162 63753
rect 360290 63744 360346 63753
rect 360162 63702 360290 63730
rect 360106 63679 360162 63688
rect 360290 63679 360346 63688
rect 360106 40216 360162 40225
rect 360290 40216 360346 40225
rect 360162 40174 360290 40202
rect 360106 40151 360162 40160
rect 360290 40151 360346 40160
rect 360396 4894 360424 337470
rect 361684 4962 361712 337690
rect 361776 337346 361804 340068
rect 361868 340054 362250 340082
rect 362328 340054 362710 340082
rect 363156 340054 363262 340082
rect 361764 337340 361816 337346
rect 361764 337282 361816 337288
rect 361672 4956 361724 4962
rect 361672 4898 361724 4904
rect 360384 4888 360436 4894
rect 360384 4830 360436 4836
rect 359740 4004 359792 4010
rect 359740 3946 359792 3952
rect 359464 3120 359516 3126
rect 359464 3062 359516 3068
rect 358544 604 358596 610
rect 358544 546 358596 552
rect 358728 604 358780 610
rect 358728 546 358780 552
rect 358556 480 358584 546
rect 359752 480 359780 3946
rect 360936 3664 360988 3670
rect 360936 3606 360988 3612
rect 360948 480 360976 3606
rect 361868 3602 361896 340054
rect 362328 337754 362356 340054
rect 362868 337816 362920 337822
rect 362868 337758 362920 337764
rect 362316 337748 362368 337754
rect 362316 337690 362368 337696
rect 362224 336864 362276 336870
rect 362224 336806 362276 336812
rect 362132 4140 362184 4146
rect 362132 4082 362184 4088
rect 361856 3596 361908 3602
rect 361856 3538 361908 3544
rect 362144 480 362172 4082
rect 362236 2922 362264 336806
rect 362880 4146 362908 337758
rect 363052 337748 363104 337754
rect 363052 337690 363104 337696
rect 363064 4826 363092 337690
rect 363052 4820 363104 4826
rect 363052 4762 363104 4768
rect 362868 4140 362920 4146
rect 362868 4082 362920 4088
rect 363156 3534 363184 340054
rect 363708 337550 363736 340068
rect 363800 340054 364182 340082
rect 363800 337754 363828 340054
rect 364248 338020 364300 338026
rect 364248 337962 364300 337968
rect 363788 337748 363840 337754
rect 363788 337690 363840 337696
rect 363696 337544 363748 337550
rect 363696 337486 363748 337492
rect 363604 336796 363656 336802
rect 363604 336738 363656 336744
rect 363328 4140 363380 4146
rect 363328 4082 363380 4088
rect 363144 3528 363196 3534
rect 363144 3470 363196 3476
rect 362224 2916 362276 2922
rect 362224 2858 362276 2864
rect 363340 480 363368 4082
rect 363616 3466 363644 336738
rect 364260 4146 364288 337962
rect 364720 336802 364748 340068
rect 365180 336870 365208 340068
rect 365640 337890 365668 340068
rect 365824 340054 366206 340082
rect 365628 337884 365680 337890
rect 365628 337826 365680 337832
rect 365168 336864 365220 336870
rect 365168 336806 365220 336812
rect 364708 336796 364760 336802
rect 364708 336738 364760 336744
rect 365626 123040 365682 123049
rect 365626 122975 365682 122984
rect 365640 122913 365668 122975
rect 365626 122904 365682 122913
rect 365626 122839 365682 122848
rect 365720 4684 365772 4690
rect 365720 4626 365772 4632
rect 364248 4140 364300 4146
rect 364248 4082 364300 4088
rect 363604 3460 363656 3466
rect 363604 3402 363656 3408
rect 365536 3324 365588 3330
rect 365536 3266 365588 3272
rect 365548 3058 365576 3266
rect 364524 3052 364576 3058
rect 364524 2994 364576 3000
rect 365536 3052 365588 3058
rect 365536 2994 365588 3000
rect 364536 480 364564 2994
rect 365732 480 365760 4626
rect 365824 3942 365852 340054
rect 366652 337210 366680 340068
rect 367126 340054 367232 340082
rect 366916 337340 366968 337346
rect 366916 337282 366968 337288
rect 366640 337204 366692 337210
rect 366640 337146 366692 337152
rect 366928 251546 366956 337282
rect 367008 328500 367060 328506
rect 367008 328442 367060 328448
rect 367020 328370 367048 328442
rect 367008 328364 367060 328370
rect 367008 328306 367060 328312
rect 367008 318844 367060 318850
rect 367008 318786 367060 318792
rect 367020 309126 367048 318786
rect 367008 309120 367060 309126
rect 367008 309062 367060 309068
rect 367008 299532 367060 299538
rect 367008 299474 367060 299480
rect 367020 289814 367048 299474
rect 367008 289808 367060 289814
rect 367008 289750 367060 289756
rect 367008 280220 367060 280226
rect 367008 280162 367060 280168
rect 367020 270502 367048 280162
rect 367008 270496 367060 270502
rect 367008 270438 367060 270444
rect 367008 260908 367060 260914
rect 367008 260850 367060 260856
rect 366836 251518 366956 251546
rect 366836 251326 366864 251518
rect 367020 251462 367048 260850
rect 367008 251456 367060 251462
rect 367008 251398 367060 251404
rect 366824 251320 366876 251326
rect 366824 251262 366876 251268
rect 366916 251252 366968 251258
rect 366916 251194 366968 251200
rect 367008 251252 367060 251258
rect 367008 251194 367060 251200
rect 366822 183560 366878 183569
rect 366822 183495 366878 183504
rect 366836 174078 366864 183495
rect 366824 174072 366876 174078
rect 366824 174014 366876 174020
rect 366732 154556 366784 154562
rect 366732 154498 366784 154504
rect 366744 144945 366772 154498
rect 366730 144936 366786 144945
rect 366730 144871 366786 144880
rect 366732 115932 366784 115938
rect 366732 115874 366784 115880
rect 366744 106321 366772 115874
rect 366730 106312 366786 106321
rect 366730 106247 366786 106256
rect 366928 87242 366956 251194
rect 367020 251122 367048 251194
rect 367008 251116 367060 251122
rect 367008 251058 367060 251064
rect 367008 241528 367060 241534
rect 367008 241470 367060 241476
rect 367020 231810 367048 241470
rect 367008 231804 367060 231810
rect 367008 231746 367060 231752
rect 367008 222216 367060 222222
rect 367008 222158 367060 222164
rect 367020 212498 367048 222158
rect 367008 212492 367060 212498
rect 367008 212434 367060 212440
rect 367008 202904 367060 202910
rect 367008 202846 367060 202852
rect 367020 193186 367048 202846
rect 367008 193180 367060 193186
rect 367008 193122 367060 193128
rect 367008 183592 367060 183598
rect 367006 183560 367008 183569
rect 367060 183560 367062 183569
rect 367006 183495 367062 183504
rect 367008 174072 367060 174078
rect 367008 174014 367060 174020
rect 367020 173913 367048 174014
rect 367006 173904 367062 173913
rect 367006 173839 367062 173848
rect 367006 164248 367062 164257
rect 367006 164183 367008 164192
rect 367060 164183 367062 164192
rect 367008 164154 367060 164160
rect 367008 154692 367060 154698
rect 367008 154634 367060 154640
rect 367020 154562 367048 154634
rect 367008 154556 367060 154562
rect 367008 154498 367060 154504
rect 367006 144936 367062 144945
rect 367006 144871 367008 144880
rect 367060 144871 367062 144880
rect 367008 144842 367060 144848
rect 367008 135380 367060 135386
rect 367008 135322 367060 135328
rect 367020 135250 367048 135322
rect 367008 135244 367060 135250
rect 367008 135186 367060 135192
rect 367008 125656 367060 125662
rect 367008 125598 367060 125604
rect 367020 115938 367048 125598
rect 367008 115932 367060 115938
rect 367008 115874 367060 115880
rect 367006 106312 367062 106321
rect 367006 106247 367008 106256
rect 367060 106247 367062 106256
rect 367008 106218 367060 106224
rect 367008 96756 367060 96762
rect 367008 96698 367060 96704
rect 367020 87281 367048 96698
rect 367006 87272 367062 87281
rect 366916 87236 366968 87242
rect 367006 87207 367062 87216
rect 366916 87178 366968 87184
rect 367006 87136 367062 87145
rect 366916 87100 366968 87106
rect 367006 87071 367062 87080
rect 366916 87042 366968 87048
rect 366928 48521 366956 87042
rect 367020 85542 367048 87071
rect 367008 85536 367060 85542
rect 367008 85478 367060 85484
rect 367008 75948 367060 75954
rect 367008 75890 367060 75896
rect 367020 66230 367048 75890
rect 367008 66224 367060 66230
rect 367008 66166 367060 66172
rect 366914 48512 366970 48521
rect 366914 48447 366970 48456
rect 367008 48408 367060 48414
rect 366914 48376 366970 48385
rect 367008 48350 367060 48356
rect 366914 48311 366970 48320
rect 366928 38758 366956 48311
rect 367020 46918 367048 48350
rect 367008 46912 367060 46918
rect 367008 46854 367060 46860
rect 366916 38752 366968 38758
rect 366916 38694 366968 38700
rect 366916 38616 366968 38622
rect 366916 38558 366968 38564
rect 366824 37324 366876 37330
rect 366824 37266 366876 37272
rect 366836 29238 366864 37266
rect 366824 29232 366876 29238
rect 366824 29174 366876 29180
rect 366928 12510 366956 38558
rect 367098 29200 367154 29209
rect 367008 29164 367060 29170
rect 367098 29135 367154 29144
rect 367008 29106 367060 29112
rect 367020 27606 367048 29106
rect 367112 29073 367140 29135
rect 367098 29064 367154 29073
rect 367098 28999 367154 29008
rect 367008 27600 367060 27606
rect 367008 27542 367060 27548
rect 366916 12504 366968 12510
rect 366916 12446 366968 12452
rect 366916 12368 366968 12374
rect 366916 12310 366968 12316
rect 366824 9716 366876 9722
rect 366824 9658 366876 9664
rect 366836 9602 366864 9658
rect 366744 9574 366864 9602
rect 366744 4434 366772 9574
rect 366928 4690 366956 12310
rect 367204 5030 367232 340054
rect 367664 337074 367692 340068
rect 367940 340054 368138 340082
rect 367652 337068 367704 337074
rect 367652 337010 367704 337016
rect 367940 335374 367968 340054
rect 367284 335368 367336 335374
rect 367284 335310 367336 335316
rect 367928 335368 367980 335374
rect 367928 335310 367980 335316
rect 367192 5024 367244 5030
rect 367192 4966 367244 4972
rect 366916 4684 366968 4690
rect 366916 4626 366968 4632
rect 366744 4406 366956 4434
rect 365812 3936 365864 3942
rect 365812 3878 365864 3884
rect 366928 480 366956 4406
rect 367296 2922 367324 335310
rect 368584 5098 368612 340068
rect 368676 340054 369150 340082
rect 368572 5092 368624 5098
rect 368572 5034 368624 5040
rect 368676 3738 368704 340054
rect 369124 337612 369176 337618
rect 369124 337554 369176 337560
rect 369136 3874 369164 337554
rect 369596 337414 369624 340068
rect 370056 337958 370084 340068
rect 370148 340054 370622 340082
rect 370044 337952 370096 337958
rect 370044 337894 370096 337900
rect 369584 337408 369636 337414
rect 369584 337350 369636 337356
rect 369768 337408 369820 337414
rect 369768 337350 369820 337356
rect 369676 123072 369728 123078
rect 369676 123014 369728 123020
rect 369688 122913 369716 123014
rect 369674 122904 369730 122913
rect 369674 122839 369730 122848
rect 369780 4146 369808 337350
rect 369216 4140 369268 4146
rect 369216 4082 369268 4088
rect 369768 4140 369820 4146
rect 369768 4082 369820 4088
rect 369124 3868 369176 3874
rect 369124 3810 369176 3816
rect 368664 3732 368716 3738
rect 368664 3674 368716 3680
rect 368020 3460 368072 3466
rect 368020 3402 368072 3408
rect 367284 2916 367336 2922
rect 367284 2858 367336 2864
rect 368032 480 368060 3402
rect 369228 480 369256 4082
rect 370148 3806 370176 340054
rect 371068 337618 371096 340068
rect 371528 338094 371556 340068
rect 371516 338088 371568 338094
rect 371516 338030 371568 338036
rect 371148 337952 371200 337958
rect 371148 337894 371200 337900
rect 371056 337612 371108 337618
rect 371056 337554 371108 337560
rect 370504 336796 370556 336802
rect 370504 336738 370556 336744
rect 370412 4140 370464 4146
rect 370412 4082 370464 4088
rect 370136 3800 370188 3806
rect 370136 3742 370188 3748
rect 370424 480 370452 4082
rect 370516 3194 370544 336738
rect 371160 4146 371188 337894
rect 372080 337210 372108 340068
rect 372068 337204 372120 337210
rect 372068 337146 372120 337152
rect 372540 336802 372568 340068
rect 373000 337482 373028 340068
rect 372988 337476 373040 337482
rect 372988 337418 373040 337424
rect 372528 336796 372580 336802
rect 372528 336738 372580 336744
rect 373092 328506 373120 340190
rect 373908 337612 373960 337618
rect 373908 337554 373960 337560
rect 372712 328500 372764 328506
rect 372712 328442 372764 328448
rect 373080 328500 373132 328506
rect 373080 328442 373132 328448
rect 372724 318782 372752 328442
rect 372712 318776 372764 318782
rect 372712 318718 372764 318724
rect 372712 309188 372764 309194
rect 372712 309130 372764 309136
rect 372724 299470 372752 309130
rect 372712 299464 372764 299470
rect 372712 299406 372764 299412
rect 372712 289876 372764 289882
rect 372712 289818 372764 289824
rect 372724 280158 372752 289818
rect 372712 280152 372764 280158
rect 372712 280094 372764 280100
rect 372712 270564 372764 270570
rect 372712 270506 372764 270512
rect 372724 260846 372752 270506
rect 372712 260840 372764 260846
rect 372712 260782 372764 260788
rect 372712 251252 372764 251258
rect 372712 251194 372764 251200
rect 372724 241505 372752 251194
rect 372526 241496 372582 241505
rect 372526 241431 372582 241440
rect 372710 241496 372766 241505
rect 372710 241431 372766 241440
rect 372540 231878 372568 241431
rect 372528 231872 372580 231878
rect 372528 231814 372580 231820
rect 372712 231872 372764 231878
rect 372712 231814 372764 231820
rect 372724 222193 372752 231814
rect 372526 222184 372582 222193
rect 372526 222119 372582 222128
rect 372710 222184 372766 222193
rect 372710 222119 372766 222128
rect 372540 212566 372568 222119
rect 372528 212560 372580 212566
rect 372528 212502 372580 212508
rect 372712 212560 372764 212566
rect 372712 212502 372764 212508
rect 372724 202881 372752 212502
rect 372526 202872 372582 202881
rect 372526 202807 372582 202816
rect 372710 202872 372766 202881
rect 372710 202807 372766 202816
rect 372540 193254 372568 202807
rect 372528 193248 372580 193254
rect 372528 193190 372580 193196
rect 372712 193248 372764 193254
rect 372712 193190 372764 193196
rect 372724 176458 372752 193190
rect 372712 176452 372764 176458
rect 372712 176394 372764 176400
rect 372804 176452 372856 176458
rect 372804 176394 372856 176400
rect 372816 164218 372844 176394
rect 372528 164212 372580 164218
rect 372528 164154 372580 164160
rect 372804 164212 372856 164218
rect 372804 164154 372856 164160
rect 372540 154601 372568 164154
rect 372526 154592 372582 154601
rect 372526 154527 372582 154536
rect 372710 154592 372766 154601
rect 372710 154527 372766 154536
rect 372724 147778 372752 154527
rect 372632 147750 372752 147778
rect 372632 147642 372660 147750
rect 372632 147614 372752 147642
rect 372724 128058 372752 147614
rect 372724 128030 372844 128058
rect 372816 122806 372844 128030
rect 372804 122800 372856 122806
rect 372804 122742 372856 122748
rect 372804 113212 372856 113218
rect 372804 113154 372856 113160
rect 372816 103494 372844 113154
rect 372804 103488 372856 103494
rect 372804 103430 372856 103436
rect 372712 77308 372764 77314
rect 372712 77250 372764 77256
rect 372724 70394 372752 77250
rect 372632 70366 372752 70394
rect 372632 70258 372660 70366
rect 372632 70230 372752 70258
rect 372724 51082 372752 70230
rect 372632 51054 372752 51082
rect 372632 50946 372660 51054
rect 372632 50918 372752 50946
rect 372724 38622 372752 50918
rect 372712 38616 372764 38622
rect 372712 38558 372764 38564
rect 372804 38616 372856 38622
rect 372804 38558 372856 38564
rect 372816 21978 372844 38558
rect 372816 21950 373028 21978
rect 371148 4140 371200 4146
rect 371148 4082 371200 4088
rect 371608 3936 371660 3942
rect 371608 3878 371660 3884
rect 370504 3188 370556 3194
rect 370504 3130 370556 3136
rect 371620 480 371648 3878
rect 372804 3868 372856 3874
rect 372804 3810 372856 3816
rect 372816 480 372844 3810
rect 373000 3126 373028 21950
rect 373920 3874 373948 337554
rect 374012 4078 374040 340068
rect 374472 337142 374500 340068
rect 374460 337136 374512 337142
rect 374460 337078 374512 337084
rect 374564 331242 374592 340190
rect 375498 340054 375696 340082
rect 375288 337476 375340 337482
rect 375288 337418 375340 337424
rect 374104 331214 374592 331242
rect 374000 4072 374052 4078
rect 374000 4014 374052 4020
rect 373908 3868 373960 3874
rect 373908 3810 373960 3816
rect 374000 3800 374052 3806
rect 374000 3742 374052 3748
rect 372988 3120 373040 3126
rect 372988 3062 373040 3068
rect 374012 480 374040 3742
rect 374104 2990 374132 331214
rect 375300 3806 375328 337418
rect 375288 3800 375340 3806
rect 375288 3742 375340 3748
rect 375196 3732 375248 3738
rect 375196 3674 375248 3680
rect 374092 2984 374144 2990
rect 374092 2926 374144 2932
rect 375208 480 375236 3674
rect 375668 3398 375696 340054
rect 375944 337754 375972 340068
rect 376036 340054 376510 340082
rect 375932 337748 375984 337754
rect 375932 337690 375984 337696
rect 376036 336954 376064 340054
rect 375852 336926 376064 336954
rect 375852 321638 375880 336926
rect 376956 336802 376984 340068
rect 377416 337822 377444 340068
rect 377508 340054 377890 340082
rect 377404 337816 377456 337822
rect 377404 337758 377456 337764
rect 376024 336796 376076 336802
rect 376024 336738 376076 336744
rect 376944 336796 376996 336802
rect 376944 336738 376996 336744
rect 375840 321632 375892 321638
rect 375840 321574 375892 321580
rect 375932 321428 375984 321434
rect 375932 321370 375984 321376
rect 375944 289882 375972 321370
rect 375840 289876 375892 289882
rect 375840 289818 375892 289824
rect 375932 289876 375984 289882
rect 375932 289818 375984 289824
rect 375852 280158 375880 289818
rect 375840 280152 375892 280158
rect 375840 280094 375892 280100
rect 375840 270564 375892 270570
rect 375840 270506 375892 270512
rect 375852 260846 375880 270506
rect 375840 260840 375892 260846
rect 375840 260782 375892 260788
rect 375840 251252 375892 251258
rect 375840 251194 375892 251200
rect 375852 241466 375880 251194
rect 375840 241460 375892 241466
rect 375840 241402 375892 241408
rect 375840 231872 375892 231878
rect 375840 231814 375892 231820
rect 375852 222154 375880 231814
rect 375840 222148 375892 222154
rect 375840 222090 375892 222096
rect 375840 212560 375892 212566
rect 375840 212502 375892 212508
rect 375852 202842 375880 212502
rect 375840 202836 375892 202842
rect 375840 202778 375892 202784
rect 375840 193248 375892 193254
rect 375840 193190 375892 193196
rect 375852 176458 375880 193190
rect 375840 176452 375892 176458
rect 375840 176394 375892 176400
rect 375932 176452 375984 176458
rect 375932 176394 375984 176400
rect 375944 164218 375972 176394
rect 375932 164212 375984 164218
rect 375932 164154 375984 164160
rect 375840 154624 375892 154630
rect 375840 154566 375892 154572
rect 375852 147778 375880 154566
rect 375760 147750 375880 147778
rect 375760 147642 375788 147750
rect 375760 147614 375880 147642
rect 375852 130422 375880 147614
rect 375840 130416 375892 130422
rect 375840 130358 375892 130364
rect 375838 125624 375894 125633
rect 375838 125559 375840 125568
rect 375892 125559 375894 125568
rect 375840 125530 375892 125536
rect 375748 116000 375800 116006
rect 375748 115942 375800 115948
rect 375760 109070 375788 115942
rect 375748 109064 375800 109070
rect 375748 109006 375800 109012
rect 375840 108996 375892 109002
rect 375840 108938 375892 108944
rect 375852 86970 375880 108938
rect 375840 86964 375892 86970
rect 375840 86906 375892 86912
rect 375840 77308 375892 77314
rect 375840 77250 375892 77256
rect 375852 70514 375880 77250
rect 375840 70508 375892 70514
rect 375840 70450 375892 70456
rect 375840 70372 375892 70378
rect 375840 70314 375892 70320
rect 375852 51202 375880 70314
rect 375840 51196 375892 51202
rect 375840 51138 375892 51144
rect 375840 51060 375892 51066
rect 375840 51002 375892 51008
rect 375852 46918 375880 51002
rect 375748 46912 375800 46918
rect 375748 46854 375800 46860
rect 375840 46912 375892 46918
rect 375840 46854 375892 46860
rect 375760 29034 375788 46854
rect 375748 29028 375800 29034
rect 375748 28970 375800 28976
rect 375840 29028 375892 29034
rect 375840 28970 375892 28976
rect 375852 27606 375880 28970
rect 375840 27600 375892 27606
rect 375840 27542 375892 27548
rect 375840 20868 375892 20874
rect 375840 20810 375892 20816
rect 375656 3392 375708 3398
rect 375656 3334 375708 3340
rect 375852 2854 375880 20810
rect 376036 3262 376064 336738
rect 377508 335594 377536 340054
rect 378048 337000 378100 337006
rect 378048 336942 378100 336948
rect 377680 336796 377732 336802
rect 377680 336738 377732 336744
rect 377140 335566 377536 335594
rect 377140 321638 377168 335566
rect 377692 335458 377720 336738
rect 377416 335430 377720 335458
rect 377128 321632 377180 321638
rect 377128 321574 377180 321580
rect 377220 321428 377272 321434
rect 377220 321370 377272 321376
rect 377232 289882 377260 321370
rect 377128 289876 377180 289882
rect 377128 289818 377180 289824
rect 377220 289876 377272 289882
rect 377220 289818 377272 289824
rect 377140 280158 377168 289818
rect 377128 280152 377180 280158
rect 377128 280094 377180 280100
rect 377128 270564 377180 270570
rect 377128 270506 377180 270512
rect 377140 260846 377168 270506
rect 377128 260840 377180 260846
rect 377128 260782 377180 260788
rect 377128 251252 377180 251258
rect 377128 251194 377180 251200
rect 377140 241505 377168 251194
rect 376942 241496 376998 241505
rect 376942 241431 376998 241440
rect 377126 241496 377182 241505
rect 377126 241431 377182 241440
rect 376956 231878 376984 241431
rect 376944 231872 376996 231878
rect 376944 231814 376996 231820
rect 377128 231872 377180 231878
rect 377128 231814 377180 231820
rect 377140 222193 377168 231814
rect 376942 222184 376998 222193
rect 376942 222119 376998 222128
rect 377126 222184 377182 222193
rect 377126 222119 377182 222128
rect 376956 212566 376984 222119
rect 376944 212560 376996 212566
rect 376944 212502 376996 212508
rect 377128 212560 377180 212566
rect 377128 212502 377180 212508
rect 377140 202881 377168 212502
rect 376942 202872 376998 202881
rect 376942 202807 376998 202816
rect 377126 202872 377182 202881
rect 377126 202807 377182 202816
rect 376956 193254 376984 202807
rect 376944 193248 376996 193254
rect 376944 193190 376996 193196
rect 377128 193248 377180 193254
rect 377128 193190 377180 193196
rect 377140 183569 377168 193190
rect 376942 183560 376998 183569
rect 376942 183495 376998 183504
rect 377126 183560 377182 183569
rect 377126 183495 377182 183504
rect 376956 173942 376984 183495
rect 376944 173936 376996 173942
rect 376944 173878 376996 173884
rect 377036 173936 377088 173942
rect 377036 173878 377088 173884
rect 377048 166954 377076 173878
rect 377048 166926 377168 166954
rect 377140 147778 377168 166926
rect 377048 147750 377168 147778
rect 377048 147642 377076 147750
rect 377048 147614 377168 147642
rect 376116 130416 376168 130422
rect 376116 130358 376168 130364
rect 376128 125633 376156 130358
rect 377140 128602 377168 147614
rect 377140 128574 377260 128602
rect 377232 125662 377260 128574
rect 377128 125656 377180 125662
rect 376114 125624 376170 125633
rect 377128 125598 377180 125604
rect 377220 125656 377272 125662
rect 377220 125598 377272 125604
rect 376114 125559 376170 125568
rect 377140 124166 377168 125598
rect 377128 124160 377180 124166
rect 377128 124102 377180 124108
rect 376666 123176 376722 123185
rect 376666 123111 376722 123120
rect 376680 123078 376708 123111
rect 376668 123072 376720 123078
rect 376668 123014 376720 123020
rect 377036 114572 377088 114578
rect 377036 114514 377088 114520
rect 377048 109070 377076 114514
rect 377036 109064 377088 109070
rect 377036 109006 377088 109012
rect 377128 108996 377180 109002
rect 377128 108938 377180 108944
rect 377140 99482 377168 108938
rect 377128 99476 377180 99482
rect 377128 99418 377180 99424
rect 377128 99340 377180 99346
rect 377128 99282 377180 99288
rect 377140 86970 377168 99282
rect 377128 86964 377180 86970
rect 377128 86906 377180 86912
rect 377128 77308 377180 77314
rect 377128 77250 377180 77256
rect 377140 70514 377168 77250
rect 377128 70508 377180 70514
rect 377128 70450 377180 70456
rect 377128 67652 377180 67658
rect 377128 67594 377180 67600
rect 377140 51218 377168 67594
rect 377140 51190 377260 51218
rect 377232 47002 377260 51190
rect 377140 46974 377260 47002
rect 377140 46918 377168 46974
rect 377036 46912 377088 46918
rect 377036 46854 377088 46860
rect 377128 46912 377180 46918
rect 377128 46854 377180 46860
rect 377048 39930 377076 46854
rect 377048 39902 377168 39930
rect 377140 31822 377168 39902
rect 377128 31816 377180 31822
rect 377128 31758 377180 31764
rect 377128 31680 377180 31686
rect 377128 31622 377180 31628
rect 377140 22166 377168 31622
rect 377128 22160 377180 22166
rect 377128 22102 377180 22108
rect 377128 22024 377180 22030
rect 377128 21966 377180 21972
rect 377140 4010 377168 21966
rect 377128 4004 377180 4010
rect 377128 3946 377180 3952
rect 377416 3670 377444 335430
rect 378060 4146 378088 336942
rect 378428 336802 378456 340068
rect 378888 338094 378916 340068
rect 378876 338088 378928 338094
rect 378876 338030 378928 338036
rect 379348 338026 379376 340068
rect 379716 340054 379914 340082
rect 379336 338020 379388 338026
rect 379336 337962 379388 337968
rect 378416 336796 378468 336802
rect 378416 336738 378468 336744
rect 378232 157752 378284 157758
rect 378230 157720 378232 157729
rect 378284 157720 378286 157729
rect 378230 157655 378286 157664
rect 378232 134224 378284 134230
rect 378230 134192 378232 134201
rect 378284 134192 378286 134201
rect 378230 134127 378286 134136
rect 379058 87136 379114 87145
rect 379058 87071 379060 87080
rect 379112 87071 379114 87080
rect 379060 87042 379112 87048
rect 378232 76288 378284 76294
rect 378230 76256 378232 76265
rect 378284 76256 378286 76265
rect 378230 76191 378286 76200
rect 378232 63912 378284 63918
rect 378230 63880 378232 63889
rect 378284 63880 378286 63889
rect 378230 63815 378286 63824
rect 377588 4140 377640 4146
rect 377588 4082 377640 4088
rect 378048 4140 378100 4146
rect 378048 4082 378100 4088
rect 378784 4140 378836 4146
rect 378784 4082 378836 4088
rect 377404 3664 377456 3670
rect 377404 3606 377456 3612
rect 376024 3256 376076 3262
rect 376024 3198 376076 3204
rect 376392 3052 376444 3058
rect 376392 2994 376444 3000
rect 375840 2848 375892 2854
rect 375840 2790 375892 2796
rect 376404 480 376432 2994
rect 377600 480 377628 4082
rect 378796 480 378824 4082
rect 379716 3466 379744 340054
rect 380164 337748 380216 337754
rect 380164 337690 380216 337696
rect 380176 5030 380204 337690
rect 380360 337346 380388 340068
rect 380820 337890 380848 340068
rect 380808 337884 380860 337890
rect 380808 337826 380860 337832
rect 381372 337754 381400 340068
rect 381360 337748 381412 337754
rect 381360 337690 381412 337696
rect 381544 337748 381596 337754
rect 381544 337690 381596 337696
rect 380348 337340 380400 337346
rect 380348 337282 380400 337288
rect 380808 336932 380860 336938
rect 380808 336874 380860 336880
rect 380164 5024 380216 5030
rect 380164 4966 380216 4972
rect 380820 3534 380848 336874
rect 381556 4962 381584 337690
rect 381832 337686 381860 340068
rect 382292 337958 382320 340068
rect 382280 337952 382332 337958
rect 382280 337894 382332 337900
rect 382844 337754 382872 340068
rect 382832 337748 382884 337754
rect 382832 337690 382884 337696
rect 381820 337680 381872 337686
rect 381820 337622 381872 337628
rect 383304 337618 383332 340068
rect 383292 337612 383344 337618
rect 383292 337554 383344 337560
rect 383764 337482 383792 340068
rect 383856 340054 384330 340082
rect 383752 337476 383804 337482
rect 383752 337418 383804 337424
rect 382188 337408 382240 337414
rect 382188 337350 382240 337356
rect 381636 336864 381688 336870
rect 381636 336806 381688 336812
rect 381544 4956 381596 4962
rect 381544 4898 381596 4904
rect 379980 3528 380032 3534
rect 379980 3470 380032 3476
rect 380808 3528 380860 3534
rect 380808 3470 380860 3476
rect 381176 3528 381228 3534
rect 381176 3470 381228 3476
rect 379704 3460 379756 3466
rect 379704 3402 379756 3408
rect 379992 480 380020 3470
rect 381188 480 381216 3470
rect 381648 3058 381676 336806
rect 382200 3534 382228 337350
rect 383568 4072 383620 4078
rect 383568 4014 383620 4020
rect 382372 3596 382424 3602
rect 382372 3538 382424 3544
rect 382188 3528 382240 3534
rect 382188 3470 382240 3476
rect 381636 3052 381688 3058
rect 381636 2994 381688 3000
rect 382384 480 382412 3538
rect 383580 480 383608 4014
rect 383856 3738 383884 340054
rect 384304 337680 384356 337686
rect 384304 337622 384356 337628
rect 384316 4078 384344 337622
rect 384776 336870 384804 340068
rect 384948 337748 385000 337754
rect 384948 337690 385000 337696
rect 384764 336864 384816 336870
rect 384764 336806 384816 336812
rect 384304 4072 384356 4078
rect 384304 4014 384356 4020
rect 383844 3732 383896 3738
rect 383844 3674 383896 3680
rect 384960 610 384988 337690
rect 385236 337006 385264 340068
rect 385328 340054 385802 340082
rect 385224 337000 385276 337006
rect 385224 336942 385276 336948
rect 385328 4146 385356 340054
rect 386248 336938 386276 340068
rect 386708 337414 386736 340068
rect 386696 337408 386748 337414
rect 386696 337350 386748 337356
rect 386800 337226 386828 340190
rect 387720 337686 387748 340068
rect 388180 337754 388208 340068
rect 388444 337884 388496 337890
rect 388444 337826 388496 337832
rect 388168 337748 388220 337754
rect 388168 337690 388220 337696
rect 387708 337680 387760 337686
rect 387708 337622 387760 337628
rect 387064 337476 387116 337482
rect 387064 337418 387116 337424
rect 386616 337198 386828 337226
rect 386236 336932 386288 336938
rect 386236 336874 386288 336880
rect 386328 157752 386380 157758
rect 386326 157720 386328 157729
rect 386380 157720 386382 157729
rect 386326 157655 386382 157664
rect 386328 134224 386380 134230
rect 386326 134192 386328 134201
rect 386380 134192 386382 134201
rect 386326 134127 386382 134136
rect 386236 87100 386288 87106
rect 386236 87042 386288 87048
rect 386248 86986 386276 87042
rect 386326 87000 386382 87009
rect 386248 86958 386326 86986
rect 386326 86935 386382 86944
rect 386328 76288 386380 76294
rect 386326 76256 386328 76265
rect 386380 76256 386382 76265
rect 386326 76191 386382 76200
rect 386328 63912 386380 63918
rect 386326 63880 386328 63889
rect 386380 63880 386382 63889
rect 386326 63815 386382 63824
rect 385316 4140 385368 4146
rect 385316 4082 385368 4088
rect 386616 3602 386644 337198
rect 386604 3596 386656 3602
rect 386604 3538 386656 3544
rect 387076 2922 387104 337418
rect 388260 3528 388312 3534
rect 388260 3470 388312 3476
rect 385868 2916 385920 2922
rect 385868 2858 385920 2864
rect 387064 2916 387116 2922
rect 387064 2858 387116 2864
rect 384672 604 384724 610
rect 384672 546 384724 552
rect 384948 604 385000 610
rect 384948 546 385000 552
rect 384684 480 384712 546
rect 385880 480 385908 2858
rect 387064 2780 387116 2786
rect 387064 2722 387116 2728
rect 387076 480 387104 2722
rect 388272 480 388300 3470
rect 388456 2854 388484 337826
rect 388732 337482 388760 340068
rect 389192 337890 389220 340068
rect 389284 340054 389666 340082
rect 389180 337884 389232 337890
rect 389180 337826 389232 337832
rect 389284 337770 389312 340054
rect 389100 337742 389312 337770
rect 388720 337476 388772 337482
rect 388720 337418 388772 337424
rect 389100 3534 389128 337742
rect 389744 331242 389772 340190
rect 389284 331226 389772 331242
rect 389272 331220 389772 331226
rect 389324 331214 389456 331220
rect 389272 331162 389324 331168
rect 389508 331214 389772 331220
rect 390572 340054 390678 340082
rect 390848 340054 391138 340082
rect 391690 340054 391888 340082
rect 389456 331162 389508 331168
rect 389468 328438 389496 331162
rect 389456 328432 389508 328438
rect 389456 328374 389508 328380
rect 389548 318844 389600 318850
rect 389548 318786 389600 318792
rect 389560 311914 389588 318786
rect 389364 311908 389416 311914
rect 389364 311850 389416 311856
rect 389548 311908 389600 311914
rect 389548 311850 389600 311856
rect 389376 302258 389404 311850
rect 389180 302252 389232 302258
rect 389180 302194 389232 302200
rect 389364 302252 389416 302258
rect 389364 302194 389416 302200
rect 389192 302138 389220 302194
rect 389192 302110 389312 302138
rect 389284 292618 389312 302110
rect 389284 292590 389496 292618
rect 389468 289814 389496 292590
rect 389456 289808 389508 289814
rect 389456 289750 389508 289756
rect 389364 280220 389416 280226
rect 389364 280162 389416 280168
rect 389376 273306 389404 280162
rect 389376 273278 389496 273306
rect 389468 270502 389496 273278
rect 389456 270496 389508 270502
rect 389456 270438 389508 270444
rect 389364 260908 389416 260914
rect 389364 260850 389416 260856
rect 389376 251258 389404 260850
rect 389180 251252 389232 251258
rect 389180 251194 389232 251200
rect 389364 251252 389416 251258
rect 389364 251194 389416 251200
rect 389192 244202 389220 251194
rect 389192 244174 389312 244202
rect 389284 234682 389312 244174
rect 389284 234654 389496 234682
rect 389468 231849 389496 234654
rect 389270 231840 389326 231849
rect 389270 231775 389326 231784
rect 389454 231840 389510 231849
rect 389454 231775 389510 231784
rect 389284 222222 389312 231775
rect 389272 222216 389324 222222
rect 389272 222158 389324 222164
rect 389548 222216 389600 222222
rect 389548 222158 389600 222164
rect 389560 215422 389588 222158
rect 389548 215416 389600 215422
rect 389548 215358 389600 215364
rect 389456 215280 389508 215286
rect 389456 215222 389508 215228
rect 389468 212537 389496 215222
rect 389270 212528 389326 212537
rect 389270 212463 389326 212472
rect 389454 212528 389510 212537
rect 389454 212463 389510 212472
rect 389284 202910 389312 212463
rect 389272 202904 389324 202910
rect 389272 202846 389324 202852
rect 389548 202904 389600 202910
rect 389548 202846 389600 202852
rect 389560 196110 389588 202846
rect 389548 196104 389600 196110
rect 389548 196046 389600 196052
rect 389456 195968 389508 195974
rect 389456 195910 389508 195916
rect 389468 193225 389496 195910
rect 389270 193216 389326 193225
rect 389270 193151 389326 193160
rect 389454 193216 389510 193225
rect 389454 193151 389510 193160
rect 389284 183598 389312 193151
rect 389272 183592 389324 183598
rect 389272 183534 389324 183540
rect 389548 183592 389600 183598
rect 389548 183534 389600 183540
rect 389560 176798 389588 183534
rect 389548 176792 389600 176798
rect 389548 176734 389600 176740
rect 389456 176656 389508 176662
rect 389456 176598 389508 176604
rect 389468 122890 389496 176598
rect 389376 122862 389496 122890
rect 389376 121446 389404 122862
rect 389364 121440 389416 121446
rect 389364 121382 389416 121388
rect 389364 103556 389416 103562
rect 389364 103498 389416 103504
rect 389376 98734 389404 103498
rect 389364 98728 389416 98734
rect 389364 98670 389416 98676
rect 389272 89684 389324 89690
rect 389272 89626 389324 89632
rect 389284 86986 389312 89626
rect 389284 86958 389404 86986
rect 389376 80102 389404 86958
rect 389364 80096 389416 80102
rect 389364 80038 389416 80044
rect 389456 79960 389508 79966
rect 389456 79902 389508 79908
rect 389468 75886 389496 79902
rect 389456 75880 389508 75886
rect 389456 75822 389508 75828
rect 389364 66292 389416 66298
rect 389364 66234 389416 66240
rect 389376 57594 389404 66234
rect 389364 57588 389416 57594
rect 389364 57530 389416 57536
rect 389272 48340 389324 48346
rect 389272 48282 389324 48288
rect 389284 42106 389312 48282
rect 389192 42078 389312 42106
rect 389192 37330 389220 42078
rect 389180 37324 389232 37330
rect 389180 37266 389232 37272
rect 389364 37324 389416 37330
rect 389364 37266 389416 37272
rect 389376 31634 389404 37266
rect 389284 31606 389404 31634
rect 389284 27742 389312 31606
rect 389272 27736 389324 27742
rect 389272 27678 389324 27684
rect 389364 27736 389416 27742
rect 389364 27678 389416 27684
rect 389376 26246 389404 27678
rect 389364 26240 389416 26246
rect 389364 26182 389416 26188
rect 389364 16652 389416 16658
rect 389364 16594 389416 16600
rect 389376 16561 389404 16594
rect 389362 16552 389418 16561
rect 389362 16487 389418 16496
rect 389546 16552 389602 16561
rect 389546 16487 389602 16496
rect 389376 6934 389404 6965
rect 389560 6934 389588 16487
rect 389364 6928 389416 6934
rect 389284 6876 389364 6882
rect 389284 6870 389416 6876
rect 389548 6928 389600 6934
rect 389548 6870 389600 6876
rect 389284 6854 389404 6870
rect 389284 3534 389312 6854
rect 389088 3528 389140 3534
rect 389088 3470 389140 3476
rect 389272 3528 389324 3534
rect 389272 3470 389324 3476
rect 388444 2848 388496 2854
rect 388444 2790 388496 2796
rect 390572 1442 390600 340054
rect 390848 4146 390876 340054
rect 391860 336818 391888 340054
rect 392136 336938 392164 340068
rect 392124 336932 392176 336938
rect 392124 336874 392176 336880
rect 391860 336790 392164 336818
rect 392596 336802 392624 340068
rect 390836 4140 390888 4146
rect 390836 4082 390888 4088
rect 391848 4140 391900 4146
rect 391848 4082 391900 4088
rect 390572 1414 390692 1442
rect 389456 604 389508 610
rect 389456 546 389508 552
rect 389468 480 389496 546
rect 390664 480 390692 1414
rect 391860 480 391888 4082
rect 392136 1442 392164 336790
rect 392584 336796 392636 336802
rect 392584 336738 392636 336744
rect 393148 4078 393176 340068
rect 393608 337074 393636 340068
rect 393596 337068 393648 337074
rect 393596 337010 393648 337016
rect 393596 336932 393648 336938
rect 393596 336874 393648 336880
rect 393228 336796 393280 336802
rect 393228 336738 393280 336744
rect 393240 4146 393268 336738
rect 393608 328438 393636 336874
rect 394068 336802 394096 340068
rect 394528 340054 394634 340082
rect 394056 336796 394108 336802
rect 394056 336738 394108 336744
rect 393596 328432 393648 328438
rect 393596 328374 393648 328380
rect 393688 328432 393740 328438
rect 393688 328374 393740 328380
rect 393700 318866 393728 328374
rect 393608 318838 393728 318866
rect 393608 317422 393636 318838
rect 393596 317416 393648 317422
rect 393596 317358 393648 317364
rect 393596 307828 393648 307834
rect 393596 307770 393648 307776
rect 393608 298110 393636 307770
rect 393596 298104 393648 298110
rect 393596 298046 393648 298052
rect 393596 280220 393648 280226
rect 393596 280162 393648 280168
rect 393608 278730 393636 280162
rect 393596 278724 393648 278730
rect 393596 278666 393648 278672
rect 393596 260908 393648 260914
rect 393596 260850 393648 260856
rect 393608 259457 393636 260850
rect 393594 259448 393650 259457
rect 393594 259383 393650 259392
rect 393778 259448 393834 259457
rect 393778 259383 393834 259392
rect 393792 249830 393820 259383
rect 393596 249824 393648 249830
rect 393596 249766 393648 249772
rect 393780 249824 393832 249830
rect 393780 249766 393832 249772
rect 393608 240122 393636 249766
rect 393516 240094 393636 240122
rect 393516 238746 393544 240094
rect 393320 238740 393372 238746
rect 393320 238682 393372 238688
rect 393504 238740 393556 238746
rect 393504 238682 393556 238688
rect 393332 229129 393360 238682
rect 393318 229120 393374 229129
rect 393318 229055 393374 229064
rect 393502 229120 393558 229129
rect 393502 229055 393558 229064
rect 393516 224262 393544 229055
rect 393320 224256 393372 224262
rect 393320 224198 393372 224204
rect 393504 224256 393556 224262
rect 393504 224198 393556 224204
rect 393332 219473 393360 224198
rect 393318 219464 393374 219473
rect 393318 219399 393374 219408
rect 393502 219464 393558 219473
rect 393502 219399 393558 219408
rect 393516 204950 393544 219399
rect 393504 204944 393556 204950
rect 393504 204886 393556 204892
rect 393504 193112 393556 193118
rect 393504 193054 393556 193060
rect 393516 191826 393544 193054
rect 393504 191820 393556 191826
rect 393504 191762 393556 191768
rect 393504 183524 393556 183530
rect 393504 183466 393556 183472
rect 393516 182170 393544 183466
rect 393320 182164 393372 182170
rect 393320 182106 393372 182112
rect 393504 182164 393556 182170
rect 393504 182106 393556 182112
rect 393332 172553 393360 182106
rect 393318 172544 393374 172553
rect 393318 172479 393374 172488
rect 393594 172544 393650 172553
rect 393594 172479 393650 172488
rect 393608 163033 393636 172479
rect 393594 163024 393650 163033
rect 393594 162959 393650 162968
rect 393686 162888 393742 162897
rect 393686 162823 393688 162832
rect 393740 162823 393742 162832
rect 393688 162794 393740 162800
rect 393596 153264 393648 153270
rect 393596 153206 393648 153212
rect 393608 148510 393636 153206
rect 393596 148504 393648 148510
rect 393596 148446 393648 148452
rect 393688 142180 393740 142186
rect 393688 142122 393740 142128
rect 393700 133906 393728 142122
rect 393700 133878 393820 133906
rect 393792 131102 393820 133878
rect 393596 131096 393648 131102
rect 393596 131038 393648 131044
rect 393780 131096 393832 131102
rect 393780 131038 393832 131044
rect 393608 121689 393636 131038
rect 393594 121680 393650 121689
rect 393594 121615 393650 121624
rect 393594 121544 393650 121553
rect 393594 121479 393650 121488
rect 393608 120086 393636 121479
rect 393596 120080 393648 120086
rect 393596 120022 393648 120028
rect 393596 110492 393648 110498
rect 393596 110434 393648 110440
rect 393608 104922 393636 110434
rect 393596 104916 393648 104922
rect 393596 104858 393648 104864
rect 393688 104780 393740 104786
rect 393688 104722 393740 104728
rect 393700 100706 393728 104722
rect 393688 100700 393740 100706
rect 393688 100642 393740 100648
rect 393596 86896 393648 86902
rect 393596 86838 393648 86844
rect 393608 75834 393636 86838
rect 393608 75806 393728 75834
rect 393700 74526 393728 75806
rect 393688 74520 393740 74526
rect 393688 74462 393740 74468
rect 393780 64932 393832 64938
rect 393780 64874 393832 64880
rect 393792 55282 393820 64874
rect 393504 55276 393556 55282
rect 393504 55218 393556 55224
rect 393780 55276 393832 55282
rect 393780 55218 393832 55224
rect 393516 55185 393544 55218
rect 393502 55176 393558 55185
rect 393502 55111 393558 55120
rect 393686 55176 393742 55185
rect 393686 55111 393742 55120
rect 393700 45626 393728 55111
rect 393412 45620 393464 45626
rect 393412 45562 393464 45568
rect 393688 45620 393740 45626
rect 393688 45562 393740 45568
rect 393424 37369 393452 45562
rect 393410 37360 393466 37369
rect 393410 37295 393466 37304
rect 393594 37360 393650 37369
rect 393594 37295 393650 37304
rect 393608 37262 393636 37295
rect 393596 37256 393648 37262
rect 393596 37198 393648 37204
rect 393688 27668 393740 27674
rect 393688 27610 393740 27616
rect 393700 18086 393728 27610
rect 393688 18080 393740 18086
rect 393688 18022 393740 18028
rect 393688 17944 393740 17950
rect 393688 17886 393740 17892
rect 393700 6934 393728 17886
rect 393688 6928 393740 6934
rect 393688 6870 393740 6876
rect 394148 6928 394200 6934
rect 394148 6870 394200 6876
rect 393228 4140 393280 4146
rect 393228 4082 393280 4088
rect 393136 4072 393188 4078
rect 393136 4014 393188 4020
rect 392136 1414 393084 1442
rect 393056 480 393084 1414
rect 394160 1086 394188 6870
rect 394528 3330 394556 340054
rect 395080 336802 395108 340068
rect 395554 340054 396028 340082
rect 394608 336796 394660 336802
rect 394608 336738 394660 336744
rect 395068 336796 395120 336802
rect 395068 336738 395120 336744
rect 395896 336796 395948 336802
rect 395896 336738 395948 336744
rect 394620 3534 394648 336738
rect 395436 4140 395488 4146
rect 395436 4082 395488 4088
rect 394608 3528 394660 3534
rect 394608 3470 394660 3476
rect 394516 3324 394568 3330
rect 394516 3266 394568 3272
rect 394148 1080 394200 1086
rect 394148 1022 394200 1028
rect 394240 604 394292 610
rect 394240 546 394292 552
rect 394252 480 394280 546
rect 395448 480 395476 4082
rect 395908 3058 395936 336738
rect 395896 3052 395948 3058
rect 395896 2994 395948 3000
rect 396000 2990 396028 340054
rect 396092 336870 396120 340068
rect 396080 336864 396132 336870
rect 396080 336806 396132 336812
rect 396552 336802 396580 340068
rect 397012 337346 397040 340068
rect 397472 337890 397500 340068
rect 397460 337884 397512 337890
rect 397460 337826 397512 337832
rect 398024 337822 398052 340068
rect 398012 337816 398064 337822
rect 398012 337758 398064 337764
rect 398484 337482 398512 340068
rect 398472 337476 398524 337482
rect 398472 337418 398524 337424
rect 397000 337340 397052 337346
rect 397000 337282 397052 337288
rect 397460 337068 397512 337074
rect 397460 337010 397512 337016
rect 396540 336796 396592 336802
rect 396540 336738 396592 336744
rect 396078 87136 396134 87145
rect 396078 87071 396080 87080
rect 396132 87071 396134 87080
rect 396080 87042 396132 87048
rect 396632 4072 396684 4078
rect 396632 4014 396684 4020
rect 395988 2984 396040 2990
rect 395988 2926 396040 2932
rect 396644 480 396672 4014
rect 397472 1442 397500 337010
rect 398944 337006 398972 340068
rect 399496 338026 399524 340068
rect 399484 338020 399536 338026
rect 399484 337962 399536 337968
rect 399956 337890 399984 340068
rect 400128 338020 400180 338026
rect 400128 337962 400180 337968
rect 399484 337884 399536 337890
rect 399484 337826 399536 337832
rect 399944 337884 399996 337890
rect 399944 337826 399996 337832
rect 398932 337000 398984 337006
rect 398932 336942 398984 336948
rect 398104 336864 398156 336870
rect 398104 336806 398156 336812
rect 398116 4146 398144 336806
rect 398196 336796 398248 336802
rect 398196 336738 398248 336744
rect 398104 4140 398156 4146
rect 398104 4082 398156 4088
rect 398208 3126 398236 336738
rect 399496 3874 399524 337826
rect 399576 337816 399628 337822
rect 399576 337758 399628 337764
rect 399484 3868 399536 3874
rect 399484 3810 399536 3816
rect 399588 3806 399616 337758
rect 399576 3800 399628 3806
rect 399576 3742 399628 3748
rect 400140 3670 400168 337962
rect 400416 337550 400444 340068
rect 400404 337544 400456 337550
rect 400404 337486 400456 337492
rect 400968 337414 400996 340068
rect 400956 337408 401008 337414
rect 400956 337350 401008 337356
rect 401428 337074 401456 340068
rect 401888 337822 401916 340068
rect 402454 340054 402836 340082
rect 401876 337816 401928 337822
rect 401876 337758 401928 337764
rect 402244 337408 402296 337414
rect 402244 337350 402296 337356
rect 401416 337068 401468 337074
rect 401416 337010 401468 337016
rect 400128 3664 400180 3670
rect 400128 3606 400180 3612
rect 402256 3534 402284 337350
rect 402808 3738 402836 340054
rect 402796 3732 402848 3738
rect 402796 3674 402848 3680
rect 402900 3602 402928 340068
rect 403360 338026 403388 340068
rect 403926 340054 404308 340082
rect 403348 338020 403400 338026
rect 403348 337962 403400 337968
rect 403624 337000 403676 337006
rect 403624 336942 403676 336948
rect 402888 3596 402940 3602
rect 402888 3538 402940 3544
rect 399024 3528 399076 3534
rect 399024 3470 399076 3476
rect 402244 3528 402296 3534
rect 402244 3470 402296 3476
rect 398196 3120 398248 3126
rect 398196 3062 398248 3068
rect 397472 1414 397868 1442
rect 397840 480 397868 1414
rect 399036 480 399064 3470
rect 403636 3330 403664 336942
rect 403716 4140 403768 4146
rect 403716 4082 403768 4088
rect 400220 3324 400272 3330
rect 400220 3266 400272 3272
rect 403624 3324 403676 3330
rect 403624 3266 403676 3272
rect 400232 480 400260 3266
rect 401324 3052 401376 3058
rect 401324 2994 401376 3000
rect 401336 480 401364 2994
rect 402520 2984 402572 2990
rect 402520 2926 402572 2932
rect 402532 480 402560 2926
rect 403728 480 403756 4082
rect 404280 3466 404308 340054
rect 404372 337686 404400 340068
rect 404360 337680 404412 337686
rect 404360 337622 404412 337628
rect 404832 337618 404860 340068
rect 405398 340054 405688 340082
rect 404820 337612 404872 337618
rect 404820 337554 404872 337560
rect 405004 337068 405056 337074
rect 405004 337010 405056 337016
rect 405016 3942 405044 337010
rect 405556 87100 405608 87106
rect 405556 87042 405608 87048
rect 405568 87009 405596 87042
rect 405554 87000 405610 87009
rect 405554 86935 405610 86944
rect 405004 3936 405056 3942
rect 405004 3878 405056 3884
rect 404268 3460 404320 3466
rect 404268 3402 404320 3408
rect 405660 3194 405688 340054
rect 405844 337482 405872 340068
rect 405832 337476 405884 337482
rect 405832 337418 405884 337424
rect 405924 337340 405976 337346
rect 405924 337282 405976 337288
rect 405648 3188 405700 3194
rect 405648 3130 405700 3136
rect 404912 3052 404964 3058
rect 404912 2994 404964 3000
rect 404924 480 404952 2994
rect 405936 610 405964 337282
rect 406304 337142 406332 340068
rect 406870 340054 407068 340082
rect 406384 337544 406436 337550
rect 406384 337486 406436 337492
rect 406292 337136 406344 337142
rect 406292 337078 406344 337084
rect 406396 4010 406424 337486
rect 406384 4004 406436 4010
rect 406384 3946 406436 3952
rect 407040 3262 407068 340054
rect 407316 337550 407344 340068
rect 407304 337544 407356 337550
rect 407304 337486 407356 337492
rect 407776 337006 407804 340068
rect 408342 340054 408448 340082
rect 407764 337000 407816 337006
rect 407764 336942 407816 336948
rect 408420 5438 408448 340054
rect 408788 337754 408816 340068
rect 409248 337958 409276 340068
rect 409708 340054 409814 340082
rect 409236 337952 409288 337958
rect 409236 337894 409288 337900
rect 408776 337748 408828 337754
rect 408776 337690 408828 337696
rect 408684 337408 408736 337414
rect 408684 337350 408736 337356
rect 408408 5432 408460 5438
rect 408408 5374 408460 5380
rect 407304 3868 407356 3874
rect 407304 3810 407356 3816
rect 407028 3256 407080 3262
rect 407028 3198 407080 3204
rect 405924 604 405976 610
rect 405924 546 405976 552
rect 406108 604 406160 610
rect 406108 546 406160 552
rect 406120 480 406148 546
rect 407316 480 407344 3810
rect 408500 3800 408552 3806
rect 408500 3742 408552 3748
rect 408512 480 408540 3742
rect 408696 2530 408724 337350
rect 409708 4146 409736 340054
rect 409788 337748 409840 337754
rect 409788 337690 409840 337696
rect 409696 4140 409748 4146
rect 409696 4082 409748 4088
rect 409800 3398 409828 337690
rect 410260 336938 410288 340068
rect 410734 340054 411116 340082
rect 410248 336932 410300 336938
rect 410248 336874 410300 336880
rect 411088 4078 411116 340054
rect 411272 338094 411300 340068
rect 411260 338088 411312 338094
rect 411260 338030 411312 338036
rect 411732 337414 411760 340068
rect 412206 340054 412588 340082
rect 412456 338088 412508 338094
rect 412456 338030 412508 338036
rect 411720 337408 411772 337414
rect 411720 337350 411772 337356
rect 411904 337136 411956 337142
rect 411904 337078 411956 337084
rect 411168 336932 411220 336938
rect 411168 336874 411220 336880
rect 411076 4072 411128 4078
rect 411076 4014 411128 4020
rect 411180 3398 411208 336874
rect 409788 3392 409840 3398
rect 409788 3334 409840 3340
rect 411168 3392 411220 3398
rect 411168 3334 411220 3340
rect 410892 3324 410944 3330
rect 410892 3266 410944 3272
rect 408696 2502 409736 2530
rect 409708 480 409736 2502
rect 410904 480 410932 3266
rect 411916 3126 411944 337078
rect 412468 5370 412496 338030
rect 412456 5364 412508 5370
rect 412456 5306 412508 5312
rect 412560 3874 412588 340054
rect 412744 337346 412772 340068
rect 413218 340054 413600 340082
rect 412824 337884 412876 337890
rect 412824 337826 412876 337832
rect 412732 337340 412784 337346
rect 412732 337282 412784 337288
rect 412548 3868 412600 3874
rect 412548 3810 412600 3816
rect 412088 3664 412140 3670
rect 412088 3606 412140 3612
rect 411904 3120 411956 3126
rect 411904 3062 411956 3068
rect 412100 480 412128 3606
rect 412836 3346 412864 337826
rect 413572 337736 413600 340054
rect 413664 337890 413692 340068
rect 413652 337884 413704 337890
rect 413652 337826 413704 337832
rect 413572 337708 413968 337736
rect 413836 337340 413888 337346
rect 413836 337282 413888 337288
rect 413284 336932 413336 336938
rect 413284 336874 413336 336880
rect 413296 3806 413324 336874
rect 413848 5302 413876 337282
rect 413836 5296 413888 5302
rect 413836 5238 413888 5244
rect 413940 3806 413968 337708
rect 414216 337278 414244 340068
rect 414676 338094 414704 340068
rect 414664 338088 414716 338094
rect 414664 338030 414716 338036
rect 415136 338026 415164 340068
rect 415124 338020 415176 338026
rect 415124 337962 415176 337968
rect 415596 337618 415624 340068
rect 416162 340054 416544 340082
rect 416044 337952 416096 337958
rect 416044 337894 416096 337900
rect 415584 337612 415636 337618
rect 415584 337554 415636 337560
rect 414204 337272 414256 337278
rect 414204 337214 414256 337220
rect 415308 337272 415360 337278
rect 415308 337214 415360 337220
rect 415320 5234 415348 337214
rect 415308 5228 415360 5234
rect 415308 5170 415360 5176
rect 414480 4004 414532 4010
rect 414480 3946 414532 3952
rect 413284 3800 413336 3806
rect 413284 3742 413336 3748
rect 413468 3800 413520 3806
rect 413468 3742 413520 3748
rect 413928 3800 413980 3806
rect 413928 3742 413980 3748
rect 412836 3318 413324 3346
rect 413296 480 413324 3318
rect 413480 2990 413508 3742
rect 413468 2984 413520 2990
rect 413468 2926 413520 2932
rect 414492 480 414520 3946
rect 415676 3528 415728 3534
rect 415676 3470 415728 3476
rect 415688 480 415716 3470
rect 416056 2854 416084 337894
rect 416516 337736 416544 340054
rect 416608 337958 416636 340068
rect 416596 337952 416648 337958
rect 416596 337894 416648 337900
rect 416964 337816 417016 337822
rect 416964 337758 417016 337764
rect 416516 337708 416728 337736
rect 416596 337612 416648 337618
rect 416596 337554 416648 337560
rect 416608 5166 416636 337554
rect 416596 5160 416648 5166
rect 416596 5102 416648 5108
rect 416700 3058 416728 337708
rect 416872 3936 416924 3942
rect 416872 3878 416924 3884
rect 416688 3052 416740 3058
rect 416688 2994 416740 3000
rect 416044 2848 416096 2854
rect 416044 2790 416096 2796
rect 416884 480 416912 3878
rect 416976 3346 417004 337758
rect 417068 337142 417096 340068
rect 417620 337890 417648 340068
rect 417424 337884 417476 337890
rect 417424 337826 417476 337832
rect 417608 337884 417660 337890
rect 417608 337826 417660 337832
rect 417056 337136 417108 337142
rect 417056 337078 417108 337084
rect 417436 3670 417464 337826
rect 417976 337136 418028 337142
rect 417976 337078 418028 337084
rect 417882 157584 417938 157593
rect 417882 157519 417884 157528
rect 417936 157519 417938 157528
rect 417884 157490 417936 157496
rect 417882 134056 417938 134065
rect 417882 133991 417884 134000
rect 417936 133991 417938 134000
rect 417884 133962 417936 133968
rect 417882 123040 417938 123049
rect 417882 122975 417884 122984
rect 417936 122975 417938 122984
rect 417884 122946 417936 122952
rect 417882 110664 417938 110673
rect 417882 110599 417884 110608
rect 417936 110599 417938 110608
rect 417884 110570 417936 110576
rect 417884 87168 417936 87174
rect 417882 87136 417884 87145
rect 417936 87136 417938 87145
rect 417882 87071 417938 87080
rect 417882 76120 417938 76129
rect 417882 76055 417884 76064
rect 417936 76055 417938 76064
rect 417884 76026 417936 76032
rect 417882 63744 417938 63753
rect 417882 63679 417884 63688
rect 417936 63679 417938 63688
rect 417884 63650 417936 63656
rect 417882 40216 417938 40225
rect 417882 40151 417884 40160
rect 417936 40151 417938 40160
rect 417884 40122 417936 40128
rect 417882 29200 417938 29209
rect 417882 29135 417884 29144
rect 417936 29135 417938 29144
rect 417884 29106 417936 29112
rect 417882 16824 417938 16833
rect 417882 16759 417884 16768
rect 417936 16759 417938 16768
rect 417884 16730 417936 16736
rect 417988 5098 418016 337078
rect 417976 5092 418028 5098
rect 417976 5034 418028 5040
rect 417424 3664 417476 3670
rect 417424 3606 417476 3612
rect 418080 3534 418108 340068
rect 418540 337346 418568 340068
rect 418528 337340 418580 337346
rect 418528 337282 418580 337288
rect 419092 337142 419120 340068
rect 419552 337754 419580 340068
rect 420012 337822 420040 340068
rect 420564 338026 420592 340068
rect 420276 338020 420328 338026
rect 420276 337962 420328 337968
rect 420552 338020 420604 338026
rect 420552 337962 420604 337968
rect 420000 337816 420052 337822
rect 420000 337758 420052 337764
rect 419540 337748 419592 337754
rect 419540 337690 419592 337696
rect 420184 337680 420236 337686
rect 420184 337622 420236 337628
rect 419448 337340 419500 337346
rect 419448 337282 419500 337288
rect 419080 337136 419132 337142
rect 419080 337078 419132 337084
rect 418158 157584 418214 157593
rect 418158 157519 418160 157528
rect 418212 157519 418214 157528
rect 418160 157490 418212 157496
rect 418158 134056 418214 134065
rect 418158 133991 418160 134000
rect 418212 133991 418214 134000
rect 418160 133962 418212 133968
rect 419354 123040 419410 123049
rect 419354 122975 419356 122984
rect 419408 122975 419410 122984
rect 419356 122946 419408 122952
rect 418158 110664 418214 110673
rect 418158 110599 418160 110608
rect 418212 110599 418214 110608
rect 418160 110570 418212 110576
rect 418620 87168 418672 87174
rect 418618 87136 418620 87145
rect 418672 87136 418674 87145
rect 418618 87071 418674 87080
rect 419354 76120 419410 76129
rect 419354 76055 419356 76064
rect 419408 76055 419410 76064
rect 419356 76026 419408 76032
rect 418158 63744 418214 63753
rect 418158 63679 418160 63688
rect 418212 63679 418214 63688
rect 418160 63650 418212 63656
rect 418158 40216 418214 40225
rect 418158 40151 418160 40160
rect 418212 40151 418214 40160
rect 418160 40122 418212 40128
rect 418158 29200 418214 29209
rect 418158 29135 418160 29144
rect 418212 29135 418214 29144
rect 418160 29106 418212 29112
rect 418158 16824 418214 16833
rect 418158 16759 418160 16768
rect 418212 16759 418214 16768
rect 418160 16730 418212 16736
rect 419460 5030 419488 337282
rect 419448 5024 419500 5030
rect 419448 4966 419500 4972
rect 420196 4010 420224 337622
rect 420184 4004 420236 4010
rect 420184 3946 420236 3952
rect 420288 3942 420316 337962
rect 420736 337816 420788 337822
rect 420736 337758 420788 337764
rect 420748 4962 420776 337758
rect 420828 337748 420880 337754
rect 420828 337690 420880 337696
rect 420736 4956 420788 4962
rect 420736 4898 420788 4904
rect 420276 3936 420328 3942
rect 420276 3878 420328 3884
rect 419172 3732 419224 3738
rect 419172 3674 419224 3680
rect 418068 3528 418120 3534
rect 418068 3470 418120 3476
rect 416976 3318 418016 3346
rect 417988 480 418016 3318
rect 419184 480 419212 3674
rect 420840 3602 420868 337690
rect 421024 337346 421052 340068
rect 421484 337754 421512 340068
rect 422036 337958 422064 340068
rect 421564 337952 421616 337958
rect 421564 337894 421616 337900
rect 422024 337952 422076 337958
rect 422024 337894 422076 337900
rect 421472 337748 421524 337754
rect 421472 337690 421524 337696
rect 421012 337340 421064 337346
rect 421012 337282 421064 337288
rect 421104 337068 421156 337074
rect 421104 337010 421156 337016
rect 420368 3596 420420 3602
rect 420368 3538 420420 3544
rect 420828 3596 420880 3602
rect 420828 3538 420880 3544
rect 420380 480 420408 3538
rect 421116 3346 421144 337010
rect 421576 3738 421604 337894
rect 422496 337754 422524 340068
rect 422208 337748 422260 337754
rect 422208 337690 422260 337696
rect 422484 337748 422536 337754
rect 422484 337690 422536 337696
rect 422220 4894 422248 337690
rect 423416 337090 423444 340190
rect 423508 337278 423536 340068
rect 423496 337272 423548 337278
rect 423496 337214 423548 337220
rect 423416 337062 423628 337090
rect 422208 4888 422260 4894
rect 422208 4830 422260 4836
rect 423600 4826 423628 337062
rect 423968 336870 423996 340068
rect 424416 337748 424468 337754
rect 424416 337690 424468 337696
rect 424324 337204 424376 337210
rect 424324 337146 424376 337152
rect 423956 336864 424008 336870
rect 423956 336806 424008 336812
rect 423588 4820 423640 4826
rect 423588 4762 423640 4768
rect 423956 4004 424008 4010
rect 423956 3946 424008 3952
rect 421564 3732 421616 3738
rect 421564 3674 421616 3680
rect 422760 3460 422812 3466
rect 422760 3402 422812 3408
rect 421116 3318 421604 3346
rect 421576 480 421604 3318
rect 422772 480 422800 3402
rect 423968 480 423996 3946
rect 424336 3466 424364 337146
rect 424428 4010 424456 337690
rect 424888 337634 424916 340190
rect 424980 337822 425008 340068
rect 424968 337816 425020 337822
rect 424968 337758 425020 337764
rect 425440 337754 425468 340068
rect 425914 340054 426388 340082
rect 426466 340054 426848 340082
rect 426926 340054 427216 340082
rect 427386 340054 427768 340082
rect 425428 337748 425480 337754
rect 425428 337690 425480 337696
rect 424888 337606 425008 337634
rect 424980 4214 425008 337606
rect 426360 5778 426388 340054
rect 426440 337476 426492 337482
rect 426440 337418 426492 337424
rect 426348 5772 426400 5778
rect 426348 5714 426400 5720
rect 424968 4208 425020 4214
rect 424968 4150 425020 4156
rect 424416 4004 424468 4010
rect 424416 3946 424468 3952
rect 424324 3460 424376 3466
rect 424324 3402 424376 3408
rect 425152 3460 425204 3466
rect 425152 3402 425204 3408
rect 425164 480 425192 3402
rect 426452 3346 426480 337418
rect 426820 337006 426848 340054
rect 427188 337550 427216 340054
rect 427176 337544 427228 337550
rect 427176 337486 427228 337492
rect 427084 337136 427136 337142
rect 427084 337078 427136 337084
rect 426808 337000 426860 337006
rect 426808 336942 426860 336948
rect 427096 3670 427124 337078
rect 427740 5846 427768 340054
rect 427924 337686 427952 340068
rect 427912 337680 427964 337686
rect 427912 337622 427964 337628
rect 428384 336870 428412 340068
rect 428858 340054 429148 340082
rect 428464 337748 428516 337754
rect 428464 337690 428516 337696
rect 428372 336864 428424 336870
rect 428372 336806 428424 336812
rect 427728 5840 427780 5846
rect 427728 5782 427780 5788
rect 427084 3664 427136 3670
rect 427084 3606 427136 3612
rect 426452 3318 427584 3346
rect 428476 3330 428504 337690
rect 429120 5914 429148 340054
rect 429396 336802 429424 340068
rect 429870 340054 430160 340082
rect 430330 340054 430528 340082
rect 429844 338088 429896 338094
rect 429844 338030 429896 338036
rect 429384 336796 429436 336802
rect 429384 336738 429436 336744
rect 429856 7698 429884 338030
rect 430132 337618 430160 340054
rect 430120 337612 430172 337618
rect 430120 337554 430172 337560
rect 430396 336796 430448 336802
rect 430396 336738 430448 336744
rect 429856 7670 430160 7698
rect 429108 5908 429160 5914
rect 429108 5850 429160 5856
rect 426348 3188 426400 3194
rect 426348 3130 426400 3136
rect 426360 480 426388 3130
rect 427556 480 427584 3318
rect 428464 3324 428516 3330
rect 428464 3266 428516 3272
rect 430132 3262 430160 7670
rect 430408 5982 430436 336738
rect 430500 6050 430528 340054
rect 430868 336802 430896 340068
rect 431328 336870 431356 340068
rect 431802 340054 431908 340082
rect 431500 337204 431552 337210
rect 431500 337146 431552 337152
rect 431224 336864 431276 336870
rect 431224 336806 431276 336812
rect 431316 336864 431368 336870
rect 431316 336806 431368 336812
rect 430856 336796 430908 336802
rect 430856 336738 430908 336744
rect 430488 6044 430540 6050
rect 430488 5986 430540 5992
rect 430396 5976 430448 5982
rect 430396 5918 430448 5924
rect 431132 3664 431184 3670
rect 431132 3606 431184 3612
rect 429936 3256 429988 3262
rect 429936 3198 429988 3204
rect 430120 3256 430172 3262
rect 430120 3198 430172 3204
rect 428740 3120 428792 3126
rect 428740 3062 428792 3068
rect 428752 480 428780 3062
rect 429948 480 429976 3198
rect 431144 480 431172 3606
rect 431236 3126 431264 336806
rect 431512 318850 431540 337146
rect 431776 336796 431828 336802
rect 431776 336738 431828 336744
rect 431408 318844 431460 318850
rect 431408 318786 431460 318792
rect 431500 318844 431552 318850
rect 431500 318786 431552 318792
rect 431420 311982 431448 318786
rect 431408 311976 431460 311982
rect 431408 311918 431460 311924
rect 431500 311976 431552 311982
rect 431500 311918 431552 311924
rect 431512 302258 431540 311918
rect 431316 302252 431368 302258
rect 431316 302194 431368 302200
rect 431500 302252 431552 302258
rect 431500 302194 431552 302200
rect 431328 302138 431356 302194
rect 431328 302110 431448 302138
rect 431420 292618 431448 302110
rect 431420 292590 431540 292618
rect 431512 282946 431540 292590
rect 431316 282940 431368 282946
rect 431316 282882 431368 282888
rect 431500 282940 431552 282946
rect 431500 282882 431552 282888
rect 431328 282826 431356 282882
rect 431328 282798 431448 282826
rect 431420 273306 431448 282798
rect 431420 273278 431540 273306
rect 431512 263634 431540 273278
rect 431316 263628 431368 263634
rect 431316 263570 431368 263576
rect 431500 263628 431552 263634
rect 431500 263570 431552 263576
rect 431328 263514 431356 263570
rect 431328 263486 431448 263514
rect 431420 253994 431448 263486
rect 431420 253966 431540 253994
rect 431512 244322 431540 253966
rect 431316 244316 431368 244322
rect 431316 244258 431368 244264
rect 431500 244316 431552 244322
rect 431500 244258 431552 244264
rect 431328 244202 431356 244258
rect 431328 244174 431448 244202
rect 431420 234682 431448 244174
rect 431420 234654 431540 234682
rect 431512 225010 431540 234654
rect 431316 225004 431368 225010
rect 431316 224946 431368 224952
rect 431500 225004 431552 225010
rect 431500 224946 431552 224952
rect 431328 224890 431356 224946
rect 431328 224862 431448 224890
rect 431420 215370 431448 224862
rect 431420 215342 431540 215370
rect 431512 205698 431540 215342
rect 431316 205692 431368 205698
rect 431316 205634 431368 205640
rect 431500 205692 431552 205698
rect 431500 205634 431552 205640
rect 431328 205578 431356 205634
rect 431328 205550 431448 205578
rect 431420 196058 431448 205550
rect 431420 196030 431540 196058
rect 431512 186386 431540 196030
rect 431316 186380 431368 186386
rect 431316 186322 431368 186328
rect 431500 186380 431552 186386
rect 431500 186322 431552 186328
rect 431328 176610 431356 186322
rect 431328 176582 431540 176610
rect 431512 167074 431540 176582
rect 431316 167068 431368 167074
rect 431316 167010 431368 167016
rect 431500 167068 431552 167074
rect 431500 167010 431552 167016
rect 431328 99362 431356 167010
rect 431328 99334 431540 99362
rect 431512 89758 431540 99334
rect 431316 89752 431368 89758
rect 431316 89694 431368 89700
rect 431500 89752 431552 89758
rect 431500 89694 431552 89700
rect 431328 86970 431356 89694
rect 431316 86964 431368 86970
rect 431316 86906 431368 86912
rect 431316 77308 431368 77314
rect 431316 77250 431368 77256
rect 431328 77178 431356 77250
rect 431316 77172 431368 77178
rect 431316 77114 431368 77120
rect 431408 67652 431460 67658
rect 431408 67594 431460 67600
rect 431420 60738 431448 67594
rect 431420 60710 431540 60738
rect 431512 51082 431540 60710
rect 431328 51054 431540 51082
rect 431224 3120 431276 3126
rect 431224 3062 431276 3068
rect 431328 2922 431356 51054
rect 431788 6118 431816 336738
rect 431880 6866 431908 340054
rect 432340 336802 432368 340068
rect 432800 337142 432828 340068
rect 432788 337136 432840 337142
rect 432788 337078 432840 337084
rect 432328 336796 432380 336802
rect 432328 336738 432380 336744
rect 433156 336796 433208 336802
rect 433156 336738 433208 336744
rect 431868 6860 431920 6866
rect 431868 6802 431920 6808
rect 433168 6798 433196 336738
rect 433156 6792 433208 6798
rect 433156 6734 433208 6740
rect 433260 6662 433288 340068
rect 433720 336802 433748 340068
rect 434272 337482 434300 340068
rect 434260 337476 434312 337482
rect 434260 337418 434312 337424
rect 434076 337204 434128 337210
rect 434076 337146 434128 337152
rect 433984 336864 434036 336870
rect 433984 336806 434036 336812
rect 433708 336796 433760 336802
rect 433708 336738 433760 336744
rect 433248 6656 433300 6662
rect 433248 6598 433300 6604
rect 431776 6112 431828 6118
rect 431776 6054 431828 6060
rect 433524 5432 433576 5438
rect 433524 5374 433576 5380
rect 432328 2984 432380 2990
rect 432328 2926 432380 2932
rect 431316 2916 431368 2922
rect 431316 2858 431368 2864
rect 432340 480 432368 2926
rect 433536 480 433564 5374
rect 433996 3262 434024 336806
rect 434088 3330 434116 337146
rect 434732 336870 434760 340068
rect 434720 336864 434772 336870
rect 434720 336806 434772 336812
rect 435192 336802 435220 340068
rect 435744 338094 435772 340068
rect 435732 338088 435784 338094
rect 435732 338030 435784 338036
rect 435916 336864 435968 336870
rect 435916 336806 435968 336812
rect 434628 336796 434680 336802
rect 434628 336738 434680 336744
rect 435180 336796 435232 336802
rect 435180 336738 435232 336744
rect 434640 6730 434668 336738
rect 434720 76152 434772 76158
rect 434718 76120 434720 76129
rect 434772 76120 434774 76129
rect 434718 76055 434774 76064
rect 434628 6724 434680 6730
rect 434628 6666 434680 6672
rect 435928 6594 435956 336806
rect 436204 336802 436232 340068
rect 436664 337618 436692 340068
rect 436652 337612 436704 337618
rect 436652 337554 436704 337560
rect 437216 337550 437244 340068
rect 437676 337618 437704 340068
rect 438150 340054 438624 340082
rect 438124 337952 438176 337958
rect 438124 337894 438176 337900
rect 437296 337612 437348 337618
rect 437296 337554 437348 337560
rect 437664 337612 437716 337618
rect 437664 337554 437716 337560
rect 437204 337544 437256 337550
rect 437204 337486 437256 337492
rect 436008 336796 436060 336802
rect 436008 336738 436060 336744
rect 436192 336796 436244 336802
rect 436192 336738 436244 336744
rect 435916 6588 435968 6594
rect 435916 6530 435968 6536
rect 436020 6526 436048 336738
rect 437202 157584 437258 157593
rect 437202 157519 437204 157528
rect 437256 157519 437258 157528
rect 437204 157490 437256 157496
rect 437204 134088 437256 134094
rect 437202 134056 437204 134065
rect 437256 134056 437258 134065
rect 437202 133991 437258 134000
rect 437202 123040 437258 123049
rect 437202 122975 437204 122984
rect 437256 122975 437258 122984
rect 437204 122946 437256 122952
rect 437202 110664 437258 110673
rect 437202 110599 437204 110608
rect 437256 110599 437258 110608
rect 437204 110570 437256 110576
rect 437202 87136 437258 87145
rect 437202 87071 437204 87080
rect 437256 87071 437258 87080
rect 437204 87042 437256 87048
rect 437202 63744 437258 63753
rect 437202 63679 437204 63688
rect 437256 63679 437258 63688
rect 437204 63650 437256 63656
rect 437204 40248 437256 40254
rect 437202 40216 437204 40225
rect 437256 40216 437258 40225
rect 437202 40151 437258 40160
rect 437204 29232 437256 29238
rect 437202 29200 437204 29209
rect 437256 29200 437258 29209
rect 437202 29135 437258 29144
rect 437202 16824 437258 16833
rect 437202 16759 437204 16768
rect 437256 16759 437258 16768
rect 437204 16730 437256 16736
rect 436008 6520 436060 6526
rect 436008 6462 436060 6468
rect 437308 6390 437336 337554
rect 437388 336796 437440 336802
rect 437388 336738 437440 336744
rect 437400 6458 437428 336738
rect 437478 157584 437534 157593
rect 437478 157519 437480 157528
rect 437532 157519 437534 157528
rect 437480 157490 437532 157496
rect 437572 134088 437624 134094
rect 437570 134056 437572 134065
rect 437624 134056 437626 134065
rect 437570 133991 437626 134000
rect 437478 123040 437534 123049
rect 437478 122975 437480 122984
rect 437532 122975 437534 122984
rect 437480 122946 437532 122952
rect 437478 110664 437534 110673
rect 437478 110599 437480 110608
rect 437532 110599 437534 110608
rect 437480 110570 437532 110576
rect 437478 87136 437534 87145
rect 437478 87071 437480 87080
rect 437532 87071 437534 87080
rect 437480 87042 437532 87048
rect 437480 76152 437532 76158
rect 437478 76120 437480 76129
rect 437532 76120 437534 76129
rect 437478 76055 437534 76064
rect 437478 63744 437534 63753
rect 437478 63679 437480 63688
rect 437532 63679 437534 63688
rect 437480 63650 437532 63656
rect 437572 40248 437624 40254
rect 437570 40216 437572 40225
rect 437624 40216 437626 40225
rect 437570 40151 437626 40160
rect 437480 29232 437532 29238
rect 437478 29200 437480 29209
rect 437532 29200 437534 29209
rect 437478 29135 437534 29144
rect 437478 16824 437534 16833
rect 437478 16759 437480 16768
rect 437532 16759 437534 16768
rect 437480 16730 437532 16736
rect 437388 6452 437440 6458
rect 437388 6394 437440 6400
rect 437296 6384 437348 6390
rect 437296 6326 437348 6332
rect 437020 4140 437072 4146
rect 437020 4082 437072 4088
rect 434076 3324 434128 3330
rect 434076 3266 434128 3272
rect 433984 3256 434036 3262
rect 433984 3198 434036 3204
rect 434628 3188 434680 3194
rect 434628 3130 434680 3136
rect 434640 480 434668 3130
rect 435824 3052 435876 3058
rect 435824 2994 435876 3000
rect 435836 480 435864 2994
rect 437032 480 437060 4082
rect 438136 2854 438164 337894
rect 438596 337736 438624 340054
rect 438688 337958 438716 340068
rect 438676 337952 438728 337958
rect 438676 337894 438728 337900
rect 439148 337754 439176 340068
rect 439622 340054 440096 340082
rect 439136 337748 439188 337754
rect 438596 337708 438808 337736
rect 438676 337612 438728 337618
rect 438676 337554 438728 337560
rect 438688 6322 438716 337554
rect 438676 6316 438728 6322
rect 438676 6258 438728 6264
rect 438780 6254 438808 337708
rect 439136 337690 439188 337696
rect 439504 337476 439556 337482
rect 439504 337418 439556 337424
rect 438768 6248 438820 6254
rect 438768 6190 438820 6196
rect 439412 4072 439464 4078
rect 439412 4014 439464 4020
rect 438216 3392 438268 3398
rect 438216 3334 438268 3340
rect 438124 2848 438176 2854
rect 438124 2790 438176 2796
rect 438228 480 438256 3334
rect 439424 480 439452 4014
rect 439516 3262 439544 337418
rect 440068 7342 440096 340054
rect 440160 338026 440188 340068
rect 440148 338020 440200 338026
rect 440148 337962 440200 337968
rect 440148 337748 440200 337754
rect 440148 337690 440200 337696
rect 440056 7336 440108 7342
rect 440056 7278 440108 7284
rect 440160 6186 440188 337690
rect 440620 337618 440648 340068
rect 441094 340054 441476 340082
rect 440608 337612 440660 337618
rect 440608 337554 440660 337560
rect 441448 7410 441476 340054
rect 441632 337618 441660 340068
rect 442092 337686 442120 340068
rect 442566 340054 442856 340082
rect 442264 337816 442316 337822
rect 442264 337758 442316 337764
rect 442080 337680 442132 337686
rect 442080 337622 442132 337628
rect 441528 337612 441580 337618
rect 441528 337554 441580 337560
rect 441620 337612 441672 337618
rect 441620 337554 441672 337560
rect 441436 7404 441488 7410
rect 441436 7346 441488 7352
rect 440148 6180 440200 6186
rect 440148 6122 440200 6128
rect 440608 5364 440660 5370
rect 440608 5306 440660 5312
rect 439504 3256 439556 3262
rect 439504 3198 439556 3204
rect 440620 480 440648 5306
rect 441540 4282 441568 337554
rect 441528 4276 441580 4282
rect 441528 4218 441580 4224
rect 442276 4078 442304 337758
rect 442356 337544 442408 337550
rect 442356 337486 442408 337492
rect 442264 4072 442316 4078
rect 442264 4014 442316 4020
rect 442368 3330 442396 337486
rect 442828 7478 442856 340054
rect 442908 337680 442960 337686
rect 442908 337622 442960 337628
rect 442816 7472 442868 7478
rect 442816 7414 442868 7420
rect 442920 4350 442948 337622
rect 443104 337482 443132 340068
rect 443564 337686 443592 340068
rect 444038 340054 444236 340082
rect 443552 337680 443604 337686
rect 443552 337622 443604 337628
rect 443644 337612 443696 337618
rect 443644 337554 443696 337560
rect 443092 337476 443144 337482
rect 443092 337418 443144 337424
rect 442908 4344 442960 4350
rect 442908 4286 442960 4292
rect 443000 3868 443052 3874
rect 443000 3810 443052 3816
rect 441804 3324 441856 3330
rect 441804 3266 441856 3272
rect 442356 3324 442408 3330
rect 442356 3266 442408 3272
rect 441816 480 441844 3266
rect 443012 480 443040 3810
rect 443656 3398 443684 337554
rect 444208 7546 444236 340054
rect 444576 337822 444604 340068
rect 444564 337816 444616 337822
rect 444564 337758 444616 337764
rect 445036 337686 445064 340068
rect 444288 337680 444340 337686
rect 444288 337622 444340 337628
rect 445024 337680 445076 337686
rect 445024 337622 445076 337628
rect 444196 7540 444248 7546
rect 444196 7482 444248 7488
rect 444196 5296 444248 5302
rect 444196 5238 444248 5244
rect 443644 3392 443696 3398
rect 443644 3334 443696 3340
rect 444208 480 444236 5238
rect 444300 4418 444328 337622
rect 444392 337074 444788 337090
rect 444380 337068 444800 337074
rect 444432 337062 444748 337068
rect 444380 337010 444432 337016
rect 444748 337010 444800 337016
rect 444380 336932 444432 336938
rect 444380 336874 444432 336880
rect 444392 336802 444420 336874
rect 444380 336796 444432 336802
rect 444380 336738 444432 336744
rect 445496 8294 445524 340068
rect 446048 337822 446076 340068
rect 445668 337816 445720 337822
rect 445668 337758 445720 337764
rect 446036 337816 446088 337822
rect 446036 337758 446088 337764
rect 445576 337680 445628 337686
rect 445576 337622 445628 337628
rect 445484 8288 445536 8294
rect 445484 8230 445536 8236
rect 445588 4486 445616 337622
rect 445576 4480 445628 4486
rect 445576 4422 445628 4428
rect 444288 4412 444340 4418
rect 444288 4354 444340 4360
rect 445680 4146 445708 337758
rect 446508 337686 446536 340068
rect 446496 337680 446548 337686
rect 446496 337622 446548 337628
rect 446968 8226 446996 340068
rect 447048 337680 447100 337686
rect 447048 337622 447100 337628
rect 446956 8220 447008 8226
rect 446956 8162 447008 8168
rect 447060 4554 447088 337622
rect 447520 337550 447548 340068
rect 447994 340054 448376 340082
rect 448244 337680 448296 337686
rect 448244 337622 448296 337628
rect 447508 337544 447560 337550
rect 447508 337486 447560 337492
rect 448256 8158 448284 337622
rect 448244 8152 448296 8158
rect 448244 8094 448296 8100
rect 447784 5228 447836 5234
rect 447784 5170 447836 5176
rect 447048 4548 447100 4554
rect 447048 4490 447100 4496
rect 445668 4140 445720 4146
rect 445668 4082 445720 4088
rect 446588 4004 446640 4010
rect 446588 3946 446640 3952
rect 445392 3800 445444 3806
rect 445392 3742 445444 3748
rect 445404 480 445432 3742
rect 446600 480 446628 3946
rect 447796 480 447824 5170
rect 448348 4622 448376 340054
rect 448440 337686 448468 340068
rect 448428 337680 448480 337686
rect 448428 337622 448480 337628
rect 448992 337618 449020 340068
rect 449466 340054 449848 340082
rect 449164 337952 449216 337958
rect 449164 337894 449216 337900
rect 448980 337612 449032 337618
rect 448980 337554 449032 337560
rect 448428 337544 448480 337550
rect 448428 337486 448480 337492
rect 448336 4616 448388 4622
rect 448336 4558 448388 4564
rect 448440 4078 448468 337486
rect 448428 4072 448480 4078
rect 448428 4014 448480 4020
rect 449176 3670 449204 337894
rect 449820 4690 449848 340054
rect 449912 337686 449940 340068
rect 450464 337958 450492 340068
rect 450938 340054 451136 340082
rect 450452 337952 450504 337958
rect 450452 337894 450504 337900
rect 449900 337680 449952 337686
rect 449900 337622 449952 337628
rect 451004 337680 451056 337686
rect 451004 337622 451056 337628
rect 451016 8090 451044 337622
rect 451004 8084 451056 8090
rect 451004 8026 451056 8032
rect 451108 4758 451136 340054
rect 451188 337952 451240 337958
rect 451188 337894 451240 337900
rect 451096 4752 451148 4758
rect 451096 4694 451148 4700
rect 449808 4684 449860 4690
rect 449808 4626 449860 4632
rect 451200 4010 451228 337894
rect 451384 337686 451412 340068
rect 451844 337958 451872 340068
rect 452410 340054 452608 340082
rect 451832 337952 451884 337958
rect 451832 337894 451884 337900
rect 451372 337680 451424 337686
rect 451372 337622 451424 337628
rect 452476 337680 452528 337686
rect 452476 337622 452528 337628
rect 452488 8022 452516 337622
rect 452476 8016 452528 8022
rect 452476 7958 452528 7964
rect 452580 5506 452608 340054
rect 452856 337686 452884 340068
rect 453316 337822 453344 340068
rect 453304 337816 453356 337822
rect 453304 337758 453356 337764
rect 452844 337680 452896 337686
rect 452844 337622 452896 337628
rect 453764 337680 453816 337686
rect 453764 337622 453816 337628
rect 453776 7954 453804 337622
rect 453764 7948 453816 7954
rect 453764 7890 453816 7896
rect 452568 5500 452620 5506
rect 452568 5442 452620 5448
rect 453868 5438 453896 340068
rect 453948 337816 454000 337822
rect 453948 337758 454000 337764
rect 453856 5432 453908 5438
rect 453856 5374 453908 5380
rect 451280 5160 451332 5166
rect 451280 5102 451332 5108
rect 451188 4004 451240 4010
rect 451188 3946 451240 3952
rect 450176 3936 450228 3942
rect 450176 3878 450228 3884
rect 449164 3664 449216 3670
rect 449164 3606 449216 3612
rect 448980 2916 449032 2922
rect 448980 2858 449032 2864
rect 448992 480 449020 2858
rect 450188 480 450216 3878
rect 451292 480 451320 5102
rect 453960 3942 453988 337758
rect 454328 337686 454356 340068
rect 454788 338026 454816 340068
rect 454776 338020 454828 338026
rect 454776 337962 454828 337968
rect 454316 337680 454368 337686
rect 454316 337622 454368 337628
rect 455236 337680 455288 337686
rect 455236 337622 455288 337628
rect 454038 87272 454094 87281
rect 454038 87207 454094 87216
rect 454052 87174 454080 87207
rect 454040 87168 454092 87174
rect 454040 87110 454092 87116
rect 455248 7886 455276 337622
rect 455236 7880 455288 7886
rect 455236 7822 455288 7828
rect 455340 5370 455368 340068
rect 455604 337884 455656 337890
rect 455604 337826 455656 337832
rect 455328 5364 455380 5370
rect 455328 5306 455380 5312
rect 454868 5092 454920 5098
rect 454868 5034 454920 5040
rect 453948 3936 454000 3942
rect 453948 3878 454000 3884
rect 453672 3868 453724 3874
rect 453672 3810 453724 3816
rect 452476 3732 452528 3738
rect 452476 3674 452528 3680
rect 452488 480 452516 3674
rect 453684 480 453712 3810
rect 454880 480 454908 5034
rect 455616 2122 455644 337826
rect 455800 337686 455828 340068
rect 456274 340054 456748 340082
rect 455788 337680 455840 337686
rect 455788 337622 455840 337628
rect 456616 337680 456668 337686
rect 456616 337622 456668 337628
rect 456522 134192 456578 134201
rect 456522 134127 456524 134136
rect 456576 134127 456578 134136
rect 456524 134098 456576 134104
rect 456522 123176 456578 123185
rect 456522 123111 456524 123120
rect 456576 123111 456578 123120
rect 456524 123082 456576 123088
rect 456522 110800 456578 110809
rect 456522 110735 456524 110744
rect 456576 110735 456578 110744
rect 456524 110706 456576 110712
rect 456522 63744 456578 63753
rect 456522 63679 456524 63688
rect 456576 63679 456578 63688
rect 456524 63650 456576 63656
rect 456524 40248 456576 40254
rect 456522 40216 456524 40225
rect 456576 40216 456578 40225
rect 456522 40151 456578 40160
rect 456628 7818 456656 337622
rect 456616 7812 456668 7818
rect 456616 7754 456668 7760
rect 456720 3738 456748 340054
rect 456812 337686 456840 340068
rect 456800 337680 456852 337686
rect 456800 337622 456852 337628
rect 457272 336802 457300 340068
rect 457746 340054 458128 340082
rect 458100 337770 458128 340054
rect 458100 337742 458220 337770
rect 458192 337686 458220 337742
rect 458088 337680 458140 337686
rect 458088 337622 458140 337628
rect 458180 337680 458232 337686
rect 458180 337622 458232 337628
rect 457260 336796 457312 336802
rect 457260 336738 457312 336744
rect 457996 336796 458048 336802
rect 457996 336738 458048 336744
rect 457444 134156 457496 134162
rect 457444 134098 457496 134104
rect 457456 134065 457484 134098
rect 457442 134056 457498 134065
rect 457442 133991 457498 134000
rect 457444 123140 457496 123146
rect 457444 123082 457496 123088
rect 457456 123049 457484 123082
rect 457442 123040 457498 123049
rect 457442 122975 457498 122984
rect 457444 110764 457496 110770
rect 457444 110706 457496 110712
rect 457456 110673 457484 110706
rect 457442 110664 457498 110673
rect 457442 110599 457498 110608
rect 456890 63744 456946 63753
rect 456890 63679 456892 63688
rect 456944 63679 456946 63688
rect 456892 63650 456944 63656
rect 456892 40248 456944 40254
rect 456890 40216 456892 40225
rect 456944 40216 456946 40225
rect 456890 40151 456946 40160
rect 458008 7750 458036 336738
rect 457996 7744 458048 7750
rect 457996 7686 458048 7692
rect 458100 4962 458128 337622
rect 458284 336802 458312 340068
rect 458744 337890 458772 340068
rect 458732 337884 458784 337890
rect 458732 337826 458784 337832
rect 459204 336938 459232 340068
rect 459376 337884 459428 337890
rect 459376 337826 459428 337832
rect 459192 336932 459244 336938
rect 459192 336874 459244 336880
rect 458272 336796 458324 336802
rect 458272 336738 458324 336744
rect 459388 7682 459416 337826
rect 459652 336864 459704 336870
rect 459652 336806 459704 336812
rect 459468 336796 459520 336802
rect 459468 336738 459520 336744
rect 459376 7676 459428 7682
rect 459376 7618 459428 7624
rect 459480 5302 459508 336738
rect 459664 331226 459692 336806
rect 459756 336802 459784 340068
rect 460216 336870 460244 340068
rect 460676 337890 460704 340068
rect 460664 337884 460716 337890
rect 460664 337826 460716 337832
rect 460296 336932 460348 336938
rect 460296 336874 460348 336880
rect 460204 336864 460256 336870
rect 460204 336806 460256 336812
rect 459744 336796 459796 336802
rect 459744 336738 459796 336744
rect 459652 331220 459704 331226
rect 459652 331162 459704 331168
rect 460112 331220 460164 331226
rect 460112 331162 460164 331168
rect 460124 323626 460152 331162
rect 460032 323598 460152 323626
rect 460032 318889 460060 323598
rect 460018 318880 460074 318889
rect 460018 318815 460074 318824
rect 460202 318880 460258 318889
rect 460202 318815 460258 318824
rect 460216 317422 460244 318815
rect 460204 317416 460256 317422
rect 460204 317358 460256 317364
rect 460204 307828 460256 307834
rect 460204 307770 460256 307776
rect 460216 302410 460244 307770
rect 460124 302382 460244 302410
rect 460124 299554 460152 302382
rect 460032 299526 460152 299554
rect 460032 298110 460060 299526
rect 460020 298104 460072 298110
rect 460020 298046 460072 298052
rect 460112 288448 460164 288454
rect 460112 288390 460164 288396
rect 460124 283014 460152 288390
rect 460112 283008 460164 283014
rect 460112 282950 460164 282956
rect 460112 282804 460164 282810
rect 460112 282746 460164 282752
rect 460124 280158 460152 282746
rect 460112 280152 460164 280158
rect 460112 280094 460164 280100
rect 460112 273148 460164 273154
rect 460112 273090 460164 273096
rect 460124 270502 460152 273090
rect 460112 270496 460164 270502
rect 460112 270438 460164 270444
rect 460020 260976 460072 260982
rect 460020 260918 460072 260924
rect 460032 260846 460060 260918
rect 460020 260840 460072 260846
rect 460020 260782 460072 260788
rect 460204 260840 460256 260846
rect 460204 260782 460256 260788
rect 460216 253858 460244 260782
rect 460124 253830 460244 253858
rect 460124 251190 460152 253830
rect 460112 251184 460164 251190
rect 460112 251126 460164 251132
rect 460020 241528 460072 241534
rect 460018 241496 460020 241505
rect 460072 241496 460074 241505
rect 460018 241431 460074 241440
rect 460110 234560 460166 234569
rect 460110 234495 460166 234504
rect 460124 225078 460152 234495
rect 460112 225072 460164 225078
rect 460112 225014 460164 225020
rect 460020 224936 460072 224942
rect 460020 224878 460072 224884
rect 460032 220833 460060 224878
rect 459834 220824 459890 220833
rect 459834 220759 459890 220768
rect 460018 220824 460074 220833
rect 460018 220759 460074 220768
rect 459848 215286 459876 220759
rect 459836 215280 459888 215286
rect 459836 215222 459888 215228
rect 460020 215280 460072 215286
rect 460020 215222 460072 215228
rect 460032 211154 460060 215222
rect 460032 211126 460152 211154
rect 460124 205766 460152 211126
rect 460112 205760 460164 205766
rect 460112 205702 460164 205708
rect 460020 205624 460072 205630
rect 460020 205566 460072 205572
rect 460032 196042 460060 205566
rect 460020 196036 460072 196042
rect 460020 195978 460072 195984
rect 460112 195900 460164 195906
rect 460112 195842 460164 195848
rect 460124 193202 460152 195842
rect 460032 193174 460152 193202
rect 460032 186386 460060 193174
rect 460020 186380 460072 186386
rect 460020 186322 460072 186328
rect 460112 186312 460164 186318
rect 460112 186254 460164 186260
rect 460124 183530 460152 186254
rect 460112 183524 460164 183530
rect 460112 183466 460164 183472
rect 460112 176520 460164 176526
rect 460112 176462 460164 176468
rect 460124 169130 460152 176462
rect 459940 169102 460152 169130
rect 459940 164257 459968 169102
rect 459926 164248 459982 164257
rect 459926 164183 459982 164192
rect 460202 164248 460258 164257
rect 460202 164183 460258 164192
rect 460216 157486 460244 164183
rect 460204 157480 460256 157486
rect 460204 157422 460256 157428
rect 460020 157344 460072 157350
rect 460020 157286 460072 157292
rect 460032 147642 460060 157286
rect 460032 147614 460244 147642
rect 460216 144906 460244 147614
rect 459928 144900 459980 144906
rect 459928 144842 459980 144848
rect 460204 144900 460256 144906
rect 460204 144842 460256 144848
rect 459940 135289 459968 144842
rect 459926 135280 459982 135289
rect 459926 135215 459982 135224
rect 460110 135280 460166 135289
rect 460110 135215 460166 135224
rect 460124 128466 460152 135215
rect 460032 128438 460152 128466
rect 460032 128330 460060 128438
rect 460032 128302 460152 128330
rect 460124 109154 460152 128302
rect 460032 109126 460152 109154
rect 460032 109018 460060 109126
rect 460032 108990 460152 109018
rect 460124 106282 460152 108990
rect 459928 106276 459980 106282
rect 459928 106218 459980 106224
rect 460112 106276 460164 106282
rect 460112 106218 460164 106224
rect 459940 96665 459968 106218
rect 459926 96656 459982 96665
rect 459926 96591 459982 96600
rect 460110 96656 460166 96665
rect 460110 96591 460166 96600
rect 460124 80186 460152 96591
rect 460032 80158 460152 80186
rect 460032 70530 460060 80158
rect 460032 70502 460152 70530
rect 460124 70258 460152 70502
rect 459940 70230 460152 70258
rect 459940 67590 459968 70230
rect 459928 67584 459980 67590
rect 459928 67526 459980 67532
rect 460204 67584 460256 67590
rect 460204 67526 460256 67532
rect 460216 58018 460244 67526
rect 460124 57990 460244 58018
rect 460124 57934 460152 57990
rect 460112 57928 460164 57934
rect 460112 57870 460164 57876
rect 460020 48340 460072 48346
rect 460020 48282 460072 48288
rect 460032 48210 460060 48282
rect 460020 48204 460072 48210
rect 460020 48146 460072 48152
rect 460204 41404 460256 41410
rect 460204 41346 460256 41352
rect 460216 38622 460244 41346
rect 460204 38616 460256 38622
rect 460204 38558 460256 38564
rect 460112 31748 460164 31754
rect 460112 31690 460164 31696
rect 460124 22030 460152 31690
rect 460112 22024 460164 22030
rect 460112 21966 460164 21972
rect 459468 5296 459520 5302
rect 459468 5238 459520 5244
rect 458456 5024 458508 5030
rect 458456 4966 458508 4972
rect 458088 4956 458140 4962
rect 458088 4898 458140 4904
rect 456708 3732 456760 3738
rect 456708 3674 456760 3680
rect 457260 3528 457312 3534
rect 457260 3470 457312 3476
rect 455616 2094 456012 2122
rect 455984 626 456012 2094
rect 455984 598 456104 626
rect 456076 480 456104 598
rect 457272 480 457300 3470
rect 458468 480 458496 4966
rect 460308 3738 460336 336874
rect 460756 336864 460808 336870
rect 460756 336806 460808 336812
rect 460388 22024 460440 22030
rect 460388 21966 460440 21972
rect 460400 3806 460428 21966
rect 460768 7614 460796 336806
rect 461228 336802 461256 340068
rect 461688 336938 461716 340068
rect 462162 340054 462268 340082
rect 461676 336932 461728 336938
rect 461676 336874 461728 336880
rect 460848 336796 460900 336802
rect 460848 336738 460900 336744
rect 461216 336796 461268 336802
rect 461216 336738 461268 336744
rect 462136 336796 462188 336802
rect 462136 336738 462188 336744
rect 460756 7608 460808 7614
rect 460756 7550 460808 7556
rect 460860 5234 460888 336738
rect 460848 5228 460900 5234
rect 460848 5170 460900 5176
rect 462148 4826 462176 336738
rect 462136 4820 462188 4826
rect 462136 4762 462188 4768
rect 460388 3800 460440 3806
rect 460388 3742 460440 3748
rect 460296 3732 460348 3738
rect 460296 3674 460348 3680
rect 462240 3602 462268 340054
rect 462700 336802 462728 340068
rect 463174 340054 463464 340082
rect 463436 336920 463464 340054
rect 463620 337278 463648 340068
rect 463792 337816 463844 337822
rect 463792 337758 463844 337764
rect 463608 337272 463660 337278
rect 463608 337214 463660 337220
rect 463436 336892 463648 336920
rect 462688 336796 462740 336802
rect 462688 336738 462740 336744
rect 463516 336796 463568 336802
rect 463516 336738 463568 336744
rect 463422 87170 463478 87179
rect 463422 87105 463478 87114
rect 463528 5166 463556 336738
rect 463516 5160 463568 5166
rect 463516 5102 463568 5108
rect 463240 3800 463292 3806
rect 463240 3742 463292 3748
rect 460848 3596 460900 3602
rect 460848 3538 460900 3544
rect 462228 3596 462280 3602
rect 462228 3538 462280 3544
rect 459652 2984 459704 2990
rect 459652 2926 459704 2932
rect 459664 480 459692 2926
rect 460860 480 460888 3538
rect 462044 2780 462096 2786
rect 462044 2722 462096 2728
rect 462056 480 462084 2722
rect 463252 480 463280 3742
rect 463620 3670 463648 336892
rect 463804 321586 463832 337758
rect 464172 336802 464200 340068
rect 464646 340054 464936 340082
rect 464160 336796 464212 336802
rect 464160 336738 464212 336744
rect 464908 336734 464936 340054
rect 465092 336938 465120 340068
rect 465644 337822 465672 340068
rect 466118 340054 466316 340082
rect 465632 337816 465684 337822
rect 465632 337758 465684 337764
rect 466184 337816 466236 337822
rect 466184 337758 466236 337764
rect 465080 336932 465132 336938
rect 465080 336874 465132 336880
rect 464988 336796 465040 336802
rect 464988 336738 465040 336744
rect 464896 336728 464948 336734
rect 464896 336670 464948 336676
rect 463712 321558 463832 321586
rect 463712 316010 463740 321558
rect 463712 315982 463924 316010
rect 463896 306406 463924 315982
rect 463700 306400 463752 306406
rect 463700 306342 463752 306348
rect 463884 306400 463936 306406
rect 463884 306342 463936 306348
rect 463712 302138 463740 306342
rect 463712 302110 463832 302138
rect 463804 292618 463832 302110
rect 463804 292590 463924 292618
rect 463896 292482 463924 292590
rect 463804 292454 463924 292482
rect 463804 282962 463832 292454
rect 463712 282934 463832 282962
rect 463712 282826 463740 282934
rect 463712 282798 463832 282826
rect 463804 275330 463832 282798
rect 463792 275324 463844 275330
rect 463792 275266 463844 275272
rect 463884 270564 463936 270570
rect 463884 270506 463936 270512
rect 463896 263514 463924 270506
rect 463804 263486 463924 263514
rect 463804 260846 463832 263486
rect 463792 260840 463844 260846
rect 463792 260782 463844 260788
rect 463700 251252 463752 251258
rect 463700 251194 463752 251200
rect 463712 244202 463740 251194
rect 463712 244174 463832 244202
rect 463804 241466 463832 244174
rect 463792 241460 463844 241466
rect 463792 241402 463844 241408
rect 463976 234660 464028 234666
rect 463976 234602 464028 234608
rect 463988 231849 464016 234602
rect 463790 231840 463846 231849
rect 463790 231775 463846 231784
rect 463974 231840 464030 231849
rect 463974 231775 464030 231784
rect 463804 222222 463832 231775
rect 463792 222216 463844 222222
rect 463792 222158 463844 222164
rect 464068 222216 464120 222222
rect 464068 222158 464120 222164
rect 464080 215422 464108 222158
rect 464068 215416 464120 215422
rect 464068 215358 464120 215364
rect 463976 215280 464028 215286
rect 463976 215222 464028 215228
rect 463988 212537 464016 215222
rect 463790 212528 463846 212537
rect 463790 212463 463846 212472
rect 463974 212528 464030 212537
rect 463974 212463 464030 212472
rect 463804 202910 463832 212463
rect 463792 202904 463844 202910
rect 463792 202846 463844 202852
rect 464068 202904 464120 202910
rect 464068 202846 464120 202852
rect 464080 196110 464108 202846
rect 464068 196104 464120 196110
rect 464068 196046 464120 196052
rect 463976 195968 464028 195974
rect 463976 195910 464028 195916
rect 463988 193225 464016 195910
rect 463790 193216 463846 193225
rect 463790 193151 463846 193160
rect 463974 193216 464030 193225
rect 463974 193151 464030 193160
rect 463804 183598 463832 193151
rect 463792 183592 463844 183598
rect 463792 183534 463844 183540
rect 464068 183592 464120 183598
rect 464068 183534 464120 183540
rect 464080 173942 464108 183534
rect 463884 173936 463936 173942
rect 463884 173878 463936 173884
rect 464068 173936 464120 173942
rect 464068 173878 464120 173884
rect 463896 157434 463924 173878
rect 463712 157406 463924 157434
rect 463712 157298 463740 157406
rect 463712 157270 463832 157298
rect 463804 147762 463832 157270
rect 463792 147756 463844 147762
rect 463792 147698 463844 147704
rect 463700 144968 463752 144974
rect 463700 144910 463752 144916
rect 463712 138038 463740 144910
rect 463700 138032 463752 138038
rect 463700 137974 463752 137980
rect 463884 137964 463936 137970
rect 463884 137906 463936 137912
rect 463896 130422 463924 137906
rect 463884 130416 463936 130422
rect 463884 130358 463936 130364
rect 464068 130416 464120 130422
rect 464068 130358 464120 130364
rect 464080 125633 464108 130358
rect 463882 125624 463938 125633
rect 463882 125559 463938 125568
rect 464066 125624 464122 125633
rect 464066 125559 464122 125568
rect 463896 114594 463924 125559
rect 463896 114566 464016 114594
rect 463988 114510 464016 114566
rect 463976 114504 464028 114510
rect 463976 114446 464028 114452
rect 463884 104916 463936 104922
rect 463884 104858 463936 104864
rect 463896 95266 463924 104858
rect 463700 95260 463752 95266
rect 463700 95202 463752 95208
rect 463884 95260 463936 95266
rect 463884 95202 463936 95208
rect 463712 94178 463740 95202
rect 463700 94172 463752 94178
rect 463700 94114 463752 94120
rect 463700 87168 463752 87174
rect 463698 87136 463700 87145
rect 463752 87136 463754 87145
rect 463698 87071 463754 87080
rect 463884 85604 463936 85610
rect 463884 85546 463936 85552
rect 463700 76152 463752 76158
rect 463698 76120 463700 76129
rect 463752 76120 463754 76129
rect 463698 76055 463754 76064
rect 463896 70530 463924 85546
rect 463804 70502 463924 70530
rect 463804 70394 463832 70502
rect 463712 70366 463832 70394
rect 463608 3664 463660 3670
rect 463608 3606 463660 3612
rect 463712 610 463740 70366
rect 463792 16720 463844 16726
rect 463790 16688 463792 16697
rect 463844 16688 463846 16697
rect 463790 16623 463846 16632
rect 465000 5098 465028 336738
rect 465264 29232 465316 29238
rect 465262 29200 465264 29209
rect 465316 29200 465318 29209
rect 465262 29135 465318 29144
rect 464988 5092 465040 5098
rect 464988 5034 465040 5040
rect 465632 5024 465684 5030
rect 465632 4966 465684 4972
rect 463700 604 463752 610
rect 463700 546 463752 552
rect 464436 604 464488 610
rect 464436 546 464488 552
rect 464448 480 464476 546
rect 465644 480 465672 4966
rect 466196 4962 466224 337758
rect 466184 4956 466236 4962
rect 466184 4898 466236 4904
rect 466288 3534 466316 340054
rect 466564 336938 466592 340068
rect 467116 337822 467144 340068
rect 467104 337816 467156 337822
rect 467104 337758 467156 337764
rect 467576 337385 467604 340068
rect 468036 337822 468064 340068
rect 468602 340054 468984 340082
rect 469062 340054 469168 340082
rect 467748 337816 467800 337822
rect 467748 337758 467800 337764
rect 468024 337816 468076 337822
rect 468024 337758 468076 337764
rect 467562 337376 467618 337385
rect 467562 337311 467618 337320
rect 466368 336932 466420 336938
rect 466368 336874 466420 336880
rect 466552 336932 466604 336938
rect 466552 336874 466604 336880
rect 466380 3602 466408 336874
rect 466550 16960 466606 16969
rect 466550 16895 466606 16904
rect 466564 16726 466592 16895
rect 466552 16720 466604 16726
rect 466552 16662 466604 16668
rect 467760 4865 467788 337758
rect 467930 87272 467986 87281
rect 467930 87207 467986 87216
rect 467944 87174 467972 87207
rect 467932 87168 467984 87174
rect 467932 87110 467984 87116
rect 467930 76256 467986 76265
rect 467930 76191 467986 76200
rect 467944 76158 467972 76191
rect 467932 76152 467984 76158
rect 467932 76094 467984 76100
rect 467930 29336 467986 29345
rect 467930 29271 467986 29280
rect 467944 29238 467972 29271
rect 467932 29232 467984 29238
rect 467932 29174 467984 29180
rect 468852 11756 468904 11762
rect 468852 11698 468904 11704
rect 467746 4856 467802 4865
rect 467746 4791 467802 4800
rect 466368 3596 466420 3602
rect 466368 3538 466420 3544
rect 466276 3528 466328 3534
rect 466276 3470 466328 3476
rect 467932 3460 467984 3466
rect 467932 3402 467984 3408
rect 466828 2848 466880 2854
rect 466828 2790 466880 2796
rect 466840 480 466868 2790
rect 467944 480 467972 3402
rect 468864 3369 468892 11698
rect 468956 4826 468984 340054
rect 469036 337816 469088 337822
rect 469036 337758 469088 337764
rect 468944 4820 468996 4826
rect 468944 4762 468996 4768
rect 469048 3466 469076 337758
rect 469140 11762 469168 340054
rect 469508 337278 469536 340068
rect 469496 337272 469548 337278
rect 469496 337214 469548 337220
rect 469220 336864 469272 336870
rect 469220 336806 469272 336812
rect 469128 11756 469180 11762
rect 469128 11698 469180 11704
rect 469128 4888 469180 4894
rect 469128 4830 469180 4836
rect 469036 3460 469088 3466
rect 469036 3402 469088 3408
rect 468850 3360 468906 3369
rect 468850 3295 468906 3304
rect 469140 480 469168 4830
rect 469232 610 469260 336806
rect 469876 299470 469904 580246
rect 469956 579148 470008 579154
rect 469956 579090 470008 579096
rect 469968 322930 469996 579090
rect 470060 346390 470088 581130
rect 470152 393310 470180 581198
rect 470232 579216 470284 579222
rect 470232 579158 470284 579164
rect 470244 405686 470272 579158
rect 470336 416770 470364 581266
rect 470428 440230 470456 581334
rect 470520 463690 470548 581402
rect 471256 546446 471284 583646
rect 580724 583568 580776 583574
rect 580724 583510 580776 583516
rect 580448 583500 580500 583506
rect 580448 583442 580500 583448
rect 580356 583432 580408 583438
rect 580356 583374 580408 583380
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 580242 580212 580751
rect 580172 580236 580224 580242
rect 580172 580178 580224 580184
rect 579896 579080 579948 579086
rect 579896 579022 579948 579028
rect 579804 567180 579856 567186
rect 579804 567122 579856 567128
rect 579816 557666 579844 567122
rect 579804 557660 579856 557666
rect 579804 557602 579856 557608
rect 579804 557524 579856 557530
rect 579804 557466 579856 557472
rect 579816 557297 579844 557466
rect 579802 557288 579858 557297
rect 579802 557223 579858 557232
rect 579712 547868 579764 547874
rect 579712 547810 579764 547816
rect 471244 546440 471296 546446
rect 471244 546382 471296 546388
rect 579724 538286 579752 547810
rect 579804 546440 579856 546446
rect 579804 546382 579856 546388
rect 579816 545601 579844 546382
rect 579802 545592 579858 545601
rect 579802 545527 579858 545536
rect 579712 538280 579764 538286
rect 579712 538222 579764 538228
rect 579804 528556 579856 528562
rect 579804 528498 579856 528504
rect 579816 518974 579844 528498
rect 579804 518968 579856 518974
rect 579804 518910 579856 518916
rect 579804 510604 579856 510610
rect 579804 510546 579856 510552
rect 579816 510377 579844 510546
rect 579802 510368 579858 510377
rect 579802 510303 579858 510312
rect 579804 509244 579856 509250
rect 579804 509186 579856 509192
rect 579816 499662 579844 509186
rect 579804 499656 579856 499662
rect 579804 499598 579856 499604
rect 579804 499520 579856 499526
rect 579804 499462 579856 499468
rect 579816 498681 579844 499462
rect 579802 498672 579858 498681
rect 579802 498607 579858 498616
rect 579804 489864 579856 489870
rect 579804 489806 579856 489812
rect 579816 480282 579844 489806
rect 579804 480276 579856 480282
rect 579804 480218 579856 480224
rect 579712 470552 579764 470558
rect 579712 470494 579764 470500
rect 470508 463684 470560 463690
rect 470508 463626 470560 463632
rect 579724 460970 579752 470494
rect 579804 463684 579856 463690
rect 579804 463626 579856 463632
rect 579816 463457 579844 463626
rect 579802 463448 579858 463457
rect 579802 463383 579858 463392
rect 579712 460964 579764 460970
rect 579712 460906 579764 460912
rect 579908 451761 579936 579022
rect 580080 579012 580132 579018
rect 580080 578954 580132 578960
rect 579988 578944 580040 578950
rect 579988 578886 580040 578892
rect 579894 451752 579950 451761
rect 579894 451687 579950 451696
rect 470416 440224 470468 440230
rect 470416 440166 470468 440172
rect 579896 440224 579948 440230
rect 579896 440166 579948 440172
rect 579908 439929 579936 440166
rect 579894 439920 579950 439929
rect 579894 439855 579950 439864
rect 470324 416764 470376 416770
rect 470324 416706 470376 416712
rect 579896 416764 579948 416770
rect 579896 416706 579948 416712
rect 579908 416537 579936 416706
rect 579894 416528 579950 416537
rect 579894 416463 579950 416472
rect 579804 412616 579856 412622
rect 579804 412558 579856 412564
rect 470232 405680 470284 405686
rect 470232 405622 470284 405628
rect 579816 403034 579844 412558
rect 579896 405680 579948 405686
rect 579896 405622 579948 405628
rect 579908 404841 579936 405622
rect 579894 404832 579950 404841
rect 579894 404767 579950 404776
rect 579804 403028 579856 403034
rect 579804 402970 579856 402976
rect 470140 393304 470192 393310
rect 470140 393246 470192 393252
rect 579896 393304 579948 393310
rect 579896 393246 579948 393252
rect 579804 393236 579856 393242
rect 579804 393178 579856 393184
rect 579816 384334 579844 393178
rect 579908 393009 579936 393246
rect 579894 393000 579950 393009
rect 579894 392935 579950 392944
rect 579804 384328 579856 384334
rect 579804 384270 579856 384276
rect 580000 369617 580028 578886
rect 579986 369608 580042 369617
rect 579986 369543 580042 369552
rect 579988 361276 580040 361282
rect 579988 361218 580040 361224
rect 580000 360194 580028 361218
rect 579804 360188 579856 360194
rect 579804 360130 579856 360136
rect 579988 360188 580040 360194
rect 579988 360130 580040 360136
rect 579816 357626 579844 360130
rect 580092 357921 580120 578954
rect 580172 578876 580224 578882
rect 580172 578818 580224 578824
rect 580078 357912 580134 357921
rect 580078 357847 580134 357856
rect 579816 357598 580120 357626
rect 470048 346384 470100 346390
rect 470048 346326 470100 346332
rect 579804 346384 579856 346390
rect 579804 346326 579856 346332
rect 579816 346089 579844 346326
rect 579802 346080 579858 346089
rect 579802 346015 579858 346024
rect 580092 345098 580120 357598
rect 580080 345092 580132 345098
rect 580080 345034 580132 345040
rect 580080 344956 580132 344962
rect 580080 344898 580132 344904
rect 499580 338088 499632 338094
rect 499580 338030 499632 338036
rect 470600 337340 470652 337346
rect 470600 337282 470652 337288
rect 470692 337340 470744 337346
rect 470692 337282 470744 337288
rect 470506 337240 470562 337249
rect 470506 337175 470562 337184
rect 470520 336938 470548 337175
rect 470508 336932 470560 336938
rect 470508 336874 470560 336880
rect 469956 322924 470008 322930
rect 469956 322866 470008 322872
rect 469864 299464 469916 299470
rect 469864 299406 469916 299412
rect 470612 3346 470640 337282
rect 470704 337249 470732 337282
rect 470690 337240 470746 337249
rect 470690 337175 470746 337184
rect 492680 337204 492732 337210
rect 492680 337146 492732 337152
rect 485780 337136 485832 337142
rect 485780 337078 485832 337084
rect 477592 337068 477644 337074
rect 477592 337010 477644 337016
rect 475384 337000 475436 337006
rect 475384 336942 475436 336948
rect 471886 123176 471942 123185
rect 471886 123111 471942 123120
rect 471900 122777 471928 123111
rect 471886 122768 471942 122777
rect 471886 122703 471942 122712
rect 471886 110800 471942 110809
rect 471886 110735 471942 110744
rect 471900 110401 471928 110735
rect 471886 110392 471942 110401
rect 471886 110327 471942 110336
rect 472716 4208 472768 4214
rect 472716 4150 472768 4156
rect 470612 3318 471560 3346
rect 469220 604 469272 610
rect 469220 546 469272 552
rect 470324 604 470376 610
rect 470324 546 470376 552
rect 470336 480 470364 546
rect 471532 480 471560 3318
rect 472728 480 472756 4150
rect 475396 3058 475424 336942
rect 475568 134088 475620 134094
rect 475566 134056 475568 134065
rect 475620 134056 475622 134065
rect 475566 133991 475622 134000
rect 476026 123176 476082 123185
rect 476026 123111 476082 123120
rect 476040 123026 476068 123111
rect 476210 123040 476266 123049
rect 476040 122998 476210 123026
rect 476210 122975 476266 122984
rect 476026 110800 476082 110809
rect 476026 110735 476082 110744
rect 476040 110650 476068 110735
rect 476210 110664 476266 110673
rect 476040 110622 476210 110650
rect 476210 110599 476266 110608
rect 476026 87272 476082 87281
rect 476026 87207 476082 87216
rect 476040 87122 476068 87207
rect 476210 87136 476266 87145
rect 476040 87094 476210 87122
rect 476210 87071 476266 87080
rect 476026 29336 476082 29345
rect 476026 29271 476082 29280
rect 476040 29186 476068 29271
rect 476210 29200 476266 29209
rect 476040 29158 476210 29186
rect 476210 29135 476266 29144
rect 476304 5772 476356 5778
rect 476304 5714 476356 5720
rect 475108 3052 475160 3058
rect 475108 2994 475160 3000
rect 475384 3052 475436 3058
rect 475384 2994 475436 3000
rect 473912 2916 473964 2922
rect 473912 2858 473964 2864
rect 473924 480 473952 2858
rect 475120 480 475148 2994
rect 476316 480 476344 5714
rect 477604 3346 477632 337010
rect 482928 134088 482980 134094
rect 482926 134056 482928 134065
rect 482980 134056 482982 134065
rect 482926 133991 482982 134000
rect 482926 76528 482982 76537
rect 482926 76463 482982 76472
rect 482940 76129 482968 76463
rect 482926 76120 482982 76129
rect 482926 76055 482982 76064
rect 482926 17232 482982 17241
rect 482926 17167 482982 17176
rect 482940 16833 482968 17167
rect 482926 16824 482982 16833
rect 482926 16759 482982 16768
rect 484584 5976 484636 5982
rect 484584 5918 484636 5924
rect 483480 5908 483532 5914
rect 483480 5850 483532 5856
rect 479892 5840 479944 5846
rect 479892 5782 479944 5788
rect 477604 3318 478736 3346
rect 477500 3052 477552 3058
rect 477500 2994 477552 3000
rect 477512 480 477540 2994
rect 478708 480 478736 3318
rect 479904 480 479932 5782
rect 482284 3052 482336 3058
rect 482284 2994 482336 3000
rect 481088 2984 481140 2990
rect 481088 2926 481140 2932
rect 481100 480 481128 2926
rect 482296 480 482324 2994
rect 483492 480 483520 5850
rect 484596 480 484624 5918
rect 485792 480 485820 337078
rect 487802 134328 487858 134337
rect 487802 134263 487858 134272
rect 487816 133929 487844 134263
rect 487802 133920 487858 133929
rect 487802 133855 487858 133864
rect 487802 123312 487858 123321
rect 487802 123247 487858 123256
rect 487816 122913 487844 123247
rect 487802 122904 487858 122913
rect 487802 122839 487858 122848
rect 487802 110936 487858 110945
rect 487802 110871 487858 110880
rect 487816 110537 487844 110871
rect 487802 110528 487858 110537
rect 487802 110463 487858 110472
rect 491206 87408 491262 87417
rect 491206 87343 491262 87352
rect 491220 87009 491248 87343
rect 491206 87000 491262 87009
rect 491206 86935 491262 86944
rect 487802 76392 487858 76401
rect 487802 76327 487858 76336
rect 487816 75993 487844 76327
rect 487802 75984 487858 75993
rect 487802 75919 487858 75928
rect 491206 29472 491262 29481
rect 491206 29407 491262 29416
rect 491220 29073 491248 29407
rect 491206 29064 491262 29073
rect 491206 28999 491262 29008
rect 487802 17096 487858 17105
rect 487802 17031 487858 17040
rect 487816 16697 487844 17031
rect 487802 16688 487858 16697
rect 487802 16623 487858 16632
rect 490564 6860 490616 6866
rect 490564 6802 490616 6808
rect 488172 6112 488224 6118
rect 488172 6054 488224 6060
rect 486976 6044 487028 6050
rect 486976 5986 487028 5992
rect 486988 480 487016 5986
rect 488184 480 488212 6054
rect 489368 3188 489420 3194
rect 489368 3130 489420 3136
rect 489380 480 489408 3130
rect 490576 480 490604 6802
rect 491760 6792 491812 6798
rect 491760 6734 491812 6740
rect 491772 480 491800 6734
rect 492692 3482 492720 337146
rect 494612 87168 494664 87174
rect 494612 87110 494664 87116
rect 494624 87009 494652 87110
rect 494610 87000 494666 87009
rect 494610 86935 494666 86944
rect 492772 29096 492824 29102
rect 492770 29064 492772 29073
rect 492824 29064 492826 29073
rect 492770 28999 492826 29008
rect 495348 6724 495400 6730
rect 495348 6666 495400 6672
rect 494152 6656 494204 6662
rect 494152 6598 494204 6604
rect 492692 3454 492996 3482
rect 492968 480 492996 3454
rect 494164 480 494192 6598
rect 495360 480 495388 6666
rect 497740 6588 497792 6594
rect 497740 6530 497792 6536
rect 496544 3256 496596 3262
rect 496544 3198 496596 3204
rect 496556 480 496584 3198
rect 497752 480 497780 6530
rect 498936 6520 498988 6526
rect 498936 6462 498988 6468
rect 498948 480 498976 6462
rect 499592 3482 499620 338030
rect 527824 338020 527876 338026
rect 527824 337962 527876 337968
rect 525064 337952 525116 337958
rect 525064 337894 525116 337900
rect 523684 337884 523736 337890
rect 523684 337826 523736 337832
rect 521016 337816 521068 337822
rect 521016 337758 521068 337764
rect 506480 337748 506532 337754
rect 506480 337690 506532 337696
rect 505744 336796 505796 336802
rect 505744 336738 505796 336744
rect 502246 87272 502302 87281
rect 502246 87207 502302 87216
rect 502260 87174 502288 87207
rect 502248 87168 502300 87174
rect 502248 87110 502300 87116
rect 502246 29336 502302 29345
rect 502246 29271 502302 29280
rect 502260 29102 502288 29271
rect 502248 29096 502300 29102
rect 502248 29038 502300 29044
rect 501236 6452 501288 6458
rect 501236 6394 501288 6400
rect 499592 3454 500172 3482
rect 500144 480 500172 3454
rect 501248 480 501276 6394
rect 502432 6384 502484 6390
rect 502432 6326 502484 6332
rect 502444 480 502472 6326
rect 504824 6316 504876 6322
rect 504824 6258 504876 6264
rect 503628 3324 503680 3330
rect 503628 3266 503680 3272
rect 503640 480 503668 3266
rect 504836 480 504864 6258
rect 505756 3194 505784 336738
rect 506020 6248 506072 6254
rect 506020 6190 506072 6196
rect 505744 3188 505796 3194
rect 505744 3130 505796 3136
rect 506032 480 506060 6190
rect 506492 3482 506520 337690
rect 520924 337680 520976 337686
rect 520924 337622 520976 337628
rect 518164 337612 518216 337618
rect 518164 337554 518216 337560
rect 514024 337544 514076 337550
rect 514024 337486 514076 337492
rect 510620 337408 510672 337414
rect 510620 337350 510672 337356
rect 512642 337376 512698 337385
rect 509884 336864 509936 336870
rect 509884 336806 509936 336812
rect 509608 7336 509660 7342
rect 509608 7278 509660 7284
rect 508412 6180 508464 6186
rect 508412 6122 508464 6128
rect 506492 3454 507256 3482
rect 507228 480 507256 3454
rect 508424 480 508452 6122
rect 509620 480 509648 7278
rect 509896 3058 509924 336806
rect 510632 3482 510660 337350
rect 512642 337311 512698 337320
rect 512000 4276 512052 4282
rect 512000 4218 512052 4224
rect 510632 3454 510844 3482
rect 509884 3052 509936 3058
rect 509884 2994 509936 3000
rect 510816 480 510844 3454
rect 512012 480 512040 4218
rect 512656 3262 512684 337311
rect 513196 7404 513248 7410
rect 513196 7346 513248 7352
rect 512644 3256 512696 3262
rect 512644 3198 512696 3204
rect 513208 480 513236 7346
rect 514036 3398 514064 337486
rect 516784 337476 516836 337482
rect 516784 337418 516836 337424
rect 516796 11778 516824 337418
rect 516704 11750 516824 11778
rect 516704 6934 516732 11750
rect 516784 7472 516836 7478
rect 516784 7414 516836 7420
rect 516692 6928 516744 6934
rect 516692 6870 516744 6876
rect 515588 4344 515640 4350
rect 515588 4286 515640 4292
rect 514024 3392 514076 3398
rect 514024 3334 514076 3340
rect 514392 3324 514444 3330
rect 514392 3266 514444 3272
rect 514404 480 514432 3266
rect 515600 480 515628 4286
rect 516796 480 516824 7414
rect 516876 6928 516928 6934
rect 516876 6870 516928 6876
rect 516888 3330 516916 6870
rect 517888 3392 517940 3398
rect 517888 3334 517940 3340
rect 516876 3324 516928 3330
rect 516876 3266 516928 3272
rect 517900 480 517928 3334
rect 518176 2854 518204 337554
rect 520280 7540 520332 7546
rect 520280 7482 520332 7488
rect 519084 4412 519136 4418
rect 519084 4354 519136 4360
rect 518164 2848 518216 2854
rect 518164 2790 518216 2796
rect 519096 480 519124 4354
rect 520292 480 520320 7482
rect 520936 2922 520964 337622
rect 521028 2990 521056 337758
rect 522672 4480 522724 4486
rect 522672 4422 522724 4428
rect 521476 4140 521528 4146
rect 521476 4082 521528 4088
rect 521016 2984 521068 2990
rect 521016 2926 521068 2932
rect 520924 2916 520976 2922
rect 520924 2858 520976 2864
rect 521488 480 521516 4082
rect 522684 480 522712 4422
rect 523696 3058 523724 337826
rect 523868 8288 523920 8294
rect 523868 8230 523920 8236
rect 523684 3052 523736 3058
rect 523684 2994 523736 3000
rect 523880 480 523908 8230
rect 525076 6882 525104 337894
rect 527456 8220 527508 8226
rect 527456 8162 527508 8168
rect 524984 6854 525104 6882
rect 524984 3126 525012 6854
rect 526260 4548 526312 4554
rect 526260 4490 526312 4496
rect 525064 3392 525116 3398
rect 525064 3334 525116 3340
rect 524972 3120 525024 3126
rect 524972 3062 525024 3068
rect 525076 480 525104 3334
rect 526272 480 526300 4490
rect 527468 480 527496 8162
rect 527836 3398 527864 337962
rect 529204 337340 529256 337346
rect 529204 337282 529256 337288
rect 529216 4146 529244 337282
rect 530584 337272 530636 337278
rect 530584 337214 530636 337220
rect 529848 4616 529900 4622
rect 529848 4558 529900 4564
rect 529204 4140 529256 4146
rect 529204 4082 529256 4088
rect 528652 4072 528704 4078
rect 528652 4014 528704 4020
rect 527824 3392 527876 3398
rect 527824 3334 527876 3340
rect 528664 480 528692 4014
rect 529860 480 529888 4558
rect 530596 4078 530624 337214
rect 580092 335442 580120 344898
rect 580080 335436 580132 335442
rect 580080 335378 580132 335384
rect 580080 335300 580132 335306
rect 580080 335242 580132 335248
rect 580092 325718 580120 335242
rect 580080 325712 580132 325718
rect 579986 325680 580042 325689
rect 580080 325654 580132 325660
rect 579986 325615 580042 325624
rect 580000 316130 580028 325615
rect 580080 322924 580132 322930
rect 580080 322866 580132 322872
rect 580092 322697 580120 322866
rect 580078 322688 580134 322697
rect 580078 322623 580134 322632
rect 579988 316124 580040 316130
rect 579988 316066 580040 316072
rect 580080 315988 580132 315994
rect 580080 315930 580132 315936
rect 580092 306406 580120 315930
rect 580184 310865 580212 578818
rect 580264 578672 580316 578678
rect 580264 578614 580316 578620
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 580080 306400 580132 306406
rect 580078 306368 580080 306377
rect 580132 306368 580134 306377
rect 580078 306303 580134 306312
rect 580092 296818 580120 306303
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 299169 580212 299406
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580080 296812 580132 296818
rect 580080 296754 580132 296760
rect 580172 296676 580224 296682
rect 580172 296618 580224 296624
rect 580184 287094 580212 296618
rect 580172 287088 580224 287094
rect 580172 287030 580224 287036
rect 580172 277364 580224 277370
rect 580172 277306 580224 277312
rect 580184 275777 580212 277306
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580276 170105 580304 578614
rect 580368 181937 580396 583374
rect 580460 205329 580488 583442
rect 580632 581052 580684 581058
rect 580632 580994 580684 581000
rect 580540 578740 580592 578746
rect 580540 578682 580592 578688
rect 580552 217025 580580 578682
rect 580644 228857 580672 580994
rect 580736 252249 580764 583510
rect 580908 581120 580960 581126
rect 580908 581062 580960 581068
rect 580816 578808 580868 578814
rect 580816 578750 580868 578756
rect 580828 263945 580856 578750
rect 580920 567186 580948 581062
rect 580908 567180 580960 567186
rect 580908 567122 580960 567128
rect 580908 557592 580960 557598
rect 580908 557534 580960 557540
rect 580920 547874 580948 557534
rect 580908 547868 580960 547874
rect 580908 547810 580960 547816
rect 580908 538280 580960 538286
rect 580908 538222 580960 538228
rect 580920 528562 580948 538222
rect 580908 528556 580960 528562
rect 580908 528498 580960 528504
rect 580908 518968 580960 518974
rect 580908 518910 580960 518916
rect 580920 509250 580948 518910
rect 580908 509244 580960 509250
rect 580908 509186 580960 509192
rect 580908 499588 580960 499594
rect 580908 499530 580960 499536
rect 580920 489870 580948 499530
rect 580908 489864 580960 489870
rect 580908 489806 580960 489812
rect 580908 480276 580960 480282
rect 580908 480218 580960 480224
rect 580920 470558 580948 480218
rect 580908 470552 580960 470558
rect 580908 470494 580960 470500
rect 580908 460964 580960 460970
rect 580908 460906 580960 460912
rect 580920 412622 580948 460906
rect 580908 412616 580960 412622
rect 580908 412558 580960 412564
rect 580908 403028 580960 403034
rect 580908 402970 580960 402976
rect 580920 393310 580948 402970
rect 580908 393304 580960 393310
rect 580908 393246 580960 393252
rect 580908 384328 580960 384334
rect 580908 384270 580960 384276
rect 580920 361282 580948 384270
rect 580908 361276 580960 361282
rect 580908 361218 580960 361224
rect 580908 345092 580960 345098
rect 580908 345034 580960 345040
rect 580920 344962 580948 345034
rect 580908 344956 580960 344962
rect 580908 344898 580960 344904
rect 581000 335436 581052 335442
rect 581000 335378 581052 335384
rect 581012 335306 581040 335378
rect 581000 335300 581052 335306
rect 581000 335242 581052 335248
rect 580908 325712 580960 325718
rect 580906 325680 580908 325689
rect 580960 325680 580962 325689
rect 580906 325615 580962 325624
rect 581000 316124 581052 316130
rect 581000 316066 581052 316072
rect 581012 315994 581040 316066
rect 581000 315988 581052 315994
rect 581000 315930 581052 315936
rect 580908 306400 580960 306406
rect 580906 306368 580908 306377
rect 580960 306368 580962 306377
rect 580906 306303 580962 306312
rect 581000 296812 581052 296818
rect 581000 296754 581052 296760
rect 581012 296682 581040 296754
rect 581000 296676 581052 296682
rect 581000 296618 581052 296624
rect 580908 287088 580960 287094
rect 580908 287030 580960 287036
rect 580920 277370 580948 287030
rect 580908 277364 580960 277370
rect 580908 277306 580960 277312
rect 580814 263936 580870 263945
rect 580814 263871 580870 263880
rect 580722 252240 580778 252249
rect 580722 252175 580778 252184
rect 580630 228848 580686 228857
rect 580630 228783 580686 228792
rect 580538 217016 580594 217025
rect 580538 216951 580594 216960
rect 580446 205320 580502 205329
rect 580446 205255 580502 205264
rect 580354 181928 580410 181937
rect 580354 181863 580410 181872
rect 580262 170096 580318 170105
rect 580262 170031 580318 170040
rect 531044 8152 531096 8158
rect 531044 8094 531096 8100
rect 530584 4072 530636 4078
rect 530584 4014 530636 4020
rect 531056 480 531084 8094
rect 534540 8084 534592 8090
rect 534540 8026 534592 8032
rect 533436 4684 533488 4690
rect 533436 4626 533488 4632
rect 532240 2848 532292 2854
rect 532240 2790 532292 2796
rect 532252 480 532280 2790
rect 533448 480 533476 4626
rect 534552 480 534580 8026
rect 538128 8016 538180 8022
rect 538128 7958 538180 7964
rect 536932 4752 536984 4758
rect 536932 4694 536984 4700
rect 535736 4004 535788 4010
rect 535736 3946 535788 3952
rect 535748 480 535776 3946
rect 536944 480 536972 4694
rect 538140 480 538168 7958
rect 541716 7948 541768 7954
rect 541716 7890 541768 7896
rect 540520 5500 540572 5506
rect 540520 5442 540572 5448
rect 539324 2916 539376 2922
rect 539324 2858 539376 2864
rect 539336 480 539364 2858
rect 540532 480 540560 5442
rect 541728 480 541756 7890
rect 545304 7880 545356 7886
rect 545304 7822 545356 7828
rect 544108 5432 544160 5438
rect 544108 5374 544160 5380
rect 542912 3936 542964 3942
rect 542912 3878 542964 3884
rect 542924 480 542952 3878
rect 544120 480 544148 5374
rect 545316 480 545344 7822
rect 548892 7812 548944 7818
rect 548892 7754 548944 7760
rect 547696 5364 547748 5370
rect 547696 5306 547748 5312
rect 546500 2984 546552 2990
rect 546500 2926 546552 2932
rect 546512 480 546540 2926
rect 547708 480 547736 5306
rect 548904 480 548932 7754
rect 552388 7744 552440 7750
rect 552388 7686 552440 7692
rect 551192 5296 551244 5302
rect 551192 5238 551244 5244
rect 550088 3868 550140 3874
rect 550088 3810 550140 3816
rect 550100 480 550128 3810
rect 551204 480 551232 5238
rect 552400 480 552428 7686
rect 555976 7676 556028 7682
rect 555976 7618 556028 7624
rect 554780 5228 554832 5234
rect 554780 5170 554832 5176
rect 553584 3052 553636 3058
rect 553584 2994 553636 3000
rect 553596 480 553624 2994
rect 554792 480 554820 5170
rect 555988 480 556016 7618
rect 559564 7608 559616 7614
rect 559564 7550 559616 7556
rect 558368 5160 558420 5166
rect 558368 5102 558420 5108
rect 557172 3800 557224 3806
rect 557172 3742 557224 3748
rect 557184 480 557212 3742
rect 558380 480 558408 5102
rect 559576 480 559604 7550
rect 561956 5092 562008 5098
rect 561956 5034 562008 5040
rect 560760 3120 560812 3126
rect 560760 3062 560812 3068
rect 560772 480 560800 3062
rect 561968 480 561996 5034
rect 565544 5024 565596 5030
rect 565544 4966 565596 4972
rect 564348 3732 564400 3738
rect 564348 3674 564400 3680
rect 563152 3188 563204 3194
rect 563152 3130 563204 3136
rect 563164 480 563192 3130
rect 564360 480 564388 3674
rect 565556 480 565584 4966
rect 569040 4956 569092 4962
rect 569040 4898 569092 4904
rect 566740 3664 566792 3670
rect 566740 3606 566792 3612
rect 566752 480 566780 3606
rect 567844 3392 567896 3398
rect 567844 3334 567896 3340
rect 567856 480 567884 3334
rect 569052 480 569080 4898
rect 572628 4888 572680 4894
rect 572628 4830 572680 4836
rect 576214 4856 576270 4865
rect 571432 3596 571484 3602
rect 571432 3538 571484 3544
rect 570236 3256 570288 3262
rect 570236 3198 570288 3204
rect 570248 480 570276 3198
rect 571444 480 571472 3538
rect 572640 480 572668 4830
rect 576214 4791 576270 4800
rect 579804 4820 579856 4826
rect 575020 4140 575072 4146
rect 575020 4082 575072 4088
rect 573824 3528 573876 3534
rect 573824 3470 573876 3476
rect 573836 480 573864 3470
rect 575032 480 575060 4082
rect 576228 480 576256 4791
rect 579804 4762 579856 4768
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 577412 3324 577464 3330
rect 577412 3266 577464 3272
rect 577424 480 577452 3266
rect 578620 480 578648 3402
rect 579816 480 579844 4762
rect 582196 4072 582248 4078
rect 582196 4014 582248 4020
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582208 480 582236 4014
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 4802 583344 4858 583400
rect 3146 567296 3202 567352
rect 3146 553016 3202 553072
rect 3054 538600 3110 538656
rect 3146 509904 3202 509960
rect 2778 495488 2834 495544
rect 3146 481072 3202 481128
rect 3238 452376 3294 452432
rect 2778 437960 2834 438016
rect 2778 423680 2834 423736
rect 3238 394984 3294 395040
rect 2778 380568 2834 380624
rect 3330 366152 3386 366208
rect 3330 323040 3386 323096
rect 3330 280100 3332 280120
rect 3332 280100 3384 280120
rect 3384 280100 3386 280120
rect 3330 280064 3386 280100
rect 3146 252456 3202 252512
rect 3146 251232 3202 251288
rect 3330 236952 3386 237008
rect 2778 222536 2834 222592
rect 3330 150728 3386 150784
rect 2778 136312 2834 136368
rect 2778 122032 2834 122088
rect 4066 308760 4122 308816
rect 3974 294344 4030 294400
rect 3882 265648 3938 265704
rect 3790 208120 3846 208176
rect 3698 193840 3754 193896
rect 3606 179424 3662 179480
rect 3514 107616 3570 107672
rect 3422 93200 3478 93256
rect 2778 78920 2834 78976
rect 3330 64504 3386 64560
rect 2778 50088 2834 50144
rect 10322 337320 10378 337376
rect 3146 35844 3148 35864
rect 3148 35844 3200 35864
rect 3200 35844 3202 35864
rect 3146 35808 3202 35844
rect 3146 11600 3202 11656
rect 3146 7112 3202 7168
rect 6458 3304 6514 3360
rect 31022 582528 31078 582584
rect 293958 583072 294014 583128
rect 300306 583208 300362 583264
rect 378138 700304 378194 700360
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 460294 583344 460350 583400
rect 420274 582936 420330 582992
rect 432970 582800 433026 582856
rect 445574 582664 445630 582720
rect 462410 582528 462466 582584
rect 231122 579264 231178 579320
rect 232962 579264 233018 579320
rect 235262 579264 235318 579320
rect 237194 579264 237250 579320
rect 239402 579264 239458 579320
rect 241426 579264 241482 579320
rect 243634 579264 243690 579320
rect 245382 579264 245438 579320
rect 247866 579264 247922 579320
rect 249522 579264 249578 579320
rect 466458 579264 466514 579320
rect 468574 579264 468630 579320
rect 51630 6160 51686 6216
rect 132498 337220 132500 337240
rect 132500 337220 132552 337240
rect 132552 337220 132554 337240
rect 132498 337184 132554 337220
rect 142066 337220 142068 337240
rect 142068 337220 142120 337240
rect 142120 337220 142122 337240
rect 142066 337184 142122 337220
rect 151818 337220 151820 337240
rect 151820 337220 151872 337240
rect 151872 337220 151874 337240
rect 151818 337184 151874 337220
rect 161386 337220 161388 337240
rect 161388 337220 161440 337240
rect 161440 337220 161442 337240
rect 161386 337184 161442 337220
rect 171138 337220 171140 337240
rect 171140 337220 171192 337240
rect 171192 337220 171194 337240
rect 171138 337184 171194 337220
rect 180706 337220 180708 337240
rect 180708 337220 180760 337240
rect 180760 337220 180762 337240
rect 180706 337184 180762 337220
rect 190458 337220 190460 337240
rect 190460 337220 190512 337240
rect 190512 337220 190514 337240
rect 190458 337184 190514 337220
rect 200026 337220 200028 337240
rect 200028 337220 200080 337240
rect 200080 337220 200082 337240
rect 200026 337184 200082 337220
rect 209778 337220 209780 337240
rect 209780 337220 209832 337240
rect 209832 337220 209834 337240
rect 209778 337184 209834 337220
rect 219346 337220 219348 337240
rect 219348 337220 219400 337240
rect 219400 337220 219402 337240
rect 219346 337184 219402 337220
rect 132590 8880 132646 8936
rect 129002 7520 129058 7576
rect 208674 4800 208730 4856
rect 229190 337220 229192 337240
rect 229192 337220 229244 337240
rect 229244 337220 229246 337240
rect 229190 337184 229246 337220
rect 231950 337320 232006 337376
rect 230754 202816 230810 202872
rect 231030 202816 231086 202872
rect 230754 183504 230810 183560
rect 231030 183504 231086 183560
rect 230662 153176 230718 153232
rect 230846 153176 230902 153232
rect 232042 3304 232098 3360
rect 234618 337220 234620 337240
rect 234620 337220 234672 337240
rect 234672 337220 234674 337240
rect 234618 337184 234674 337220
rect 234894 241440 234950 241496
rect 235078 241440 235134 241496
rect 234894 222128 234950 222184
rect 235078 222128 235134 222184
rect 236274 241440 236330 241496
rect 236458 241440 236514 241496
rect 236274 222128 236330 222184
rect 236458 222128 236514 222184
rect 236274 202816 236330 202872
rect 236458 202816 236514 202872
rect 236274 183504 236330 183560
rect 236458 183504 236514 183560
rect 236274 154536 236330 154592
rect 236458 154536 236514 154592
rect 236274 135224 236330 135280
rect 236458 135224 236514 135280
rect 236274 115912 236330 115968
rect 236458 115912 236514 115968
rect 236274 96600 236330 96656
rect 236458 96600 236514 96656
rect 238114 5344 238170 5400
rect 244370 249736 244426 249792
rect 244554 249736 244610 249792
rect 245934 278704 245990 278760
rect 246118 278704 246174 278760
rect 245842 259392 245898 259448
rect 246026 259392 246082 259448
rect 245842 249772 245844 249792
rect 245844 249772 245896 249792
rect 245896 249772 245898 249792
rect 245842 249736 245898 249772
rect 246118 249736 246174 249792
rect 247314 220768 247370 220824
rect 247222 211132 247278 211168
rect 247222 211112 247224 211132
rect 247224 211112 247276 211132
rect 247276 211112 247278 211132
rect 246946 201456 247002 201512
rect 247130 201456 247186 201512
rect 244370 144880 244426 144936
rect 244554 144880 244610 144936
rect 244554 66408 244610 66464
rect 244370 66272 244426 66328
rect 245566 48184 245622 48240
rect 245750 159976 245806 160032
rect 246118 159976 246174 160032
rect 245842 143540 245898 143576
rect 245842 143520 245844 143540
rect 245844 143520 245896 143540
rect 245896 143520 245898 143540
rect 246026 143520 246082 143576
rect 245750 140664 245806 140720
rect 245934 140664 245990 140720
rect 247038 133864 247094 133920
rect 247314 133728 247370 133784
rect 245934 48320 245990 48376
rect 245750 5480 245806 5536
rect 248418 110764 248474 110800
rect 248418 110744 248420 110764
rect 248420 110744 248472 110764
rect 248472 110744 248474 110764
rect 249982 201456 250038 201512
rect 250166 201476 250222 201512
rect 250166 201456 250168 201476
rect 250168 201456 250220 201476
rect 250220 201456 250222 201476
rect 250166 116048 250222 116104
rect 250074 115912 250130 115968
rect 249982 6160 250038 6216
rect 251178 280064 251234 280120
rect 251178 260752 251234 260808
rect 251178 249736 251234 249792
rect 251086 240080 251142 240136
rect 251546 307672 251602 307728
rect 251546 298152 251602 298208
rect 251362 280064 251418 280120
rect 251362 260752 251418 260808
rect 251454 249736 251510 249792
rect 251362 240116 251364 240136
rect 251364 240116 251416 240136
rect 251416 240116 251418 240136
rect 251362 240080 251418 240116
rect 251362 230460 251364 230480
rect 251364 230460 251416 230480
rect 251416 230460 251418 230480
rect 251362 230424 251418 230460
rect 251546 230424 251602 230480
rect 251362 193160 251418 193216
rect 251546 193160 251602 193216
rect 251178 76064 251234 76120
rect 251178 75656 251234 75712
rect 251454 77288 251510 77344
rect 251638 77288 251694 77344
rect 251362 19216 251418 19272
rect 251638 19080 251694 19136
rect 251454 9696 251510 9752
rect 251638 9696 251694 9752
rect 253110 29280 253166 29336
rect 254122 110608 254178 110664
rect 257986 29180 257988 29200
rect 257988 29180 258040 29200
rect 258040 29180 258042 29200
rect 257986 29144 258042 29180
rect 259366 110628 259422 110664
rect 259366 110608 259368 110628
rect 259368 110608 259420 110628
rect 259420 110608 259422 110628
rect 259642 222128 259698 222184
rect 259734 221856 259790 221912
rect 259642 202816 259698 202872
rect 259918 202816 259974 202872
rect 259642 183504 259698 183560
rect 259918 183504 259974 183560
rect 259734 122712 259790 122768
rect 259918 122712 259974 122768
rect 262310 248376 262366 248432
rect 262586 269048 262642 269104
rect 262678 268912 262734 268968
rect 262494 248376 262550 248432
rect 262586 202852 262588 202872
rect 262588 202852 262640 202872
rect 262640 202852 262642 202872
rect 262586 202816 262642 202852
rect 262678 202680 262734 202736
rect 262586 183504 262642 183560
rect 262678 183368 262734 183424
rect 262678 135224 262734 135280
rect 262862 135224 262918 135280
rect 262678 66136 262734 66192
rect 262954 66136 263010 66192
rect 264978 193160 265034 193216
rect 265254 275984 265310 276040
rect 265530 275984 265586 276040
rect 265162 266328 265218 266384
rect 265346 266328 265402 266384
rect 265162 222164 265164 222184
rect 265164 222164 265216 222184
rect 265216 222164 265218 222184
rect 265162 222128 265218 222164
rect 265346 222164 265348 222184
rect 265348 222164 265400 222184
rect 265400 222164 265402 222184
rect 265346 222128 265402 222164
rect 265162 202816 265218 202872
rect 265346 202816 265402 202872
rect 265254 193196 265256 193216
rect 265256 193196 265308 193216
rect 265308 193196 265310 193216
rect 265254 193160 265310 193196
rect 265162 183540 265164 183560
rect 265164 183540 265216 183560
rect 265216 183540 265218 183560
rect 265162 183504 265218 183540
rect 265346 183504 265402 183560
rect 265254 125704 265310 125760
rect 265254 125568 265310 125624
rect 265622 16904 265678 16960
rect 265622 16360 265678 16416
rect 267830 306312 267886 306368
rect 268014 306312 268070 306368
rect 267738 269048 267794 269104
rect 267830 268912 267886 268968
rect 267738 222128 267794 222184
rect 267738 221992 267794 222048
rect 266634 220768 266690 220824
rect 266818 220768 266874 220824
rect 267738 202816 267794 202872
rect 267922 202816 267978 202872
rect 267738 180784 267794 180840
rect 267922 180804 267978 180840
rect 267922 180784 267924 180804
rect 267924 180784 267976 180804
rect 267976 180784 267978 180804
rect 267646 134544 267702 134600
rect 267646 134272 267702 134328
rect 266726 125704 266782 125760
rect 267830 125704 267886 125760
rect 266634 125568 266690 125624
rect 267738 125568 267794 125624
rect 267646 110472 267702 110528
rect 267738 48320 267794 48376
rect 267922 48184 267978 48240
rect 264978 8336 265034 8392
rect 265162 8336 265218 8392
rect 270498 212472 270554 212528
rect 270498 202852 270500 202872
rect 270500 202852 270552 202872
rect 270552 202852 270554 202872
rect 270498 202816 270554 202852
rect 270498 193196 270500 193216
rect 270500 193196 270552 193216
rect 270552 193196 270554 193216
rect 270498 193160 270554 193196
rect 270498 183540 270500 183560
rect 270500 183540 270552 183560
rect 270552 183540 270554 183560
rect 270498 183504 270554 183540
rect 270314 134272 270370 134328
rect 270498 134272 270554 134328
rect 270498 75964 270500 75984
rect 270500 75964 270552 75984
rect 270552 75964 270554 75984
rect 270498 75928 270554 75964
rect 270406 40160 270462 40216
rect 270406 40024 270462 40080
rect 270774 212508 270776 212528
rect 270776 212508 270828 212528
rect 270828 212508 270830 212528
rect 270774 212472 270830 212508
rect 270682 202852 270684 202872
rect 270684 202852 270736 202872
rect 270736 202852 270738 202872
rect 270682 202816 270738 202852
rect 270774 193196 270776 193216
rect 270776 193196 270828 193216
rect 270828 193196 270830 193216
rect 270774 193160 270830 193196
rect 270682 183540 270684 183560
rect 270684 183540 270736 183560
rect 270736 183540 270738 183560
rect 270682 183504 270738 183540
rect 272154 278704 272210 278760
rect 272338 278704 272394 278760
rect 272154 240080 272210 240136
rect 272338 240080 272394 240136
rect 272062 220768 272118 220824
rect 272246 220768 272302 220824
rect 272062 211112 272118 211168
rect 272246 211112 272302 211168
rect 272154 202816 272210 202872
rect 272338 202680 272394 202736
rect 272154 183504 272210 183560
rect 272338 183368 272394 183424
rect 272062 172488 272118 172544
rect 272246 172488 272302 172544
rect 272246 125704 272302 125760
rect 272154 125568 272210 125624
rect 273074 87080 273130 87136
rect 273258 87080 273314 87136
rect 273074 29144 273130 29200
rect 273258 29144 273314 29200
rect 273534 241440 273590 241496
rect 273718 241440 273774 241496
rect 273534 222128 273590 222184
rect 273718 222128 273774 222184
rect 273534 202816 273590 202872
rect 273718 202816 273774 202872
rect 273534 183504 273590 183560
rect 273718 183504 273774 183560
rect 273534 125704 273590 125760
rect 273534 125568 273590 125624
rect 273718 123256 273774 123312
rect 273902 123256 273958 123312
rect 275374 76064 275430 76120
rect 281722 278704 281778 278760
rect 281814 278568 281870 278624
rect 281722 193196 281724 193216
rect 281724 193196 281776 193216
rect 281776 193196 281778 193216
rect 281722 193160 281778 193196
rect 281906 193196 281908 193216
rect 281908 193196 281960 193216
rect 281960 193196 281962 193216
rect 281906 193160 281962 193196
rect 281722 173884 281724 173904
rect 281724 173884 281776 173904
rect 281776 173884 281778 173904
rect 281722 173848 281778 173884
rect 281906 173884 281908 173904
rect 281908 173884 281960 173904
rect 281960 173884 281962 173904
rect 281906 173848 281962 173884
rect 281722 125704 281778 125760
rect 281722 125568 281778 125624
rect 283102 7520 283158 7576
rect 284666 278704 284722 278760
rect 284850 278704 284906 278760
rect 284666 193196 284668 193216
rect 284668 193196 284720 193216
rect 284720 193196 284722 193216
rect 284666 193160 284722 193196
rect 284850 193196 284852 193216
rect 284852 193196 284904 193216
rect 284904 193196 284906 193216
rect 284850 193160 284906 193196
rect 284666 173884 284668 173904
rect 284668 173884 284720 173904
rect 284720 173884 284722 173904
rect 284666 173848 284722 173884
rect 284850 173884 284852 173904
rect 284852 173884 284904 173904
rect 284904 173884 284906 173904
rect 284850 173848 284906 173884
rect 284758 125704 284814 125760
rect 284666 125568 284722 125624
rect 284666 76064 284722 76120
rect 284758 75928 284814 75984
rect 284482 8880 284538 8936
rect 285770 325624 285826 325680
rect 285770 124208 285826 124264
rect 285954 325624 286010 325680
rect 286046 316004 286048 316024
rect 286048 316004 286100 316024
rect 286100 316004 286102 316024
rect 286046 315968 286102 316004
rect 286230 315968 286286 316024
rect 286046 238856 286102 238912
rect 285954 238740 286010 238776
rect 285954 238720 285956 238740
rect 285956 238720 286008 238740
rect 286008 238720 286010 238740
rect 285954 182144 286010 182200
rect 286138 182144 286194 182200
rect 285954 173848 286010 173904
rect 286138 173848 286194 173904
rect 286966 134136 287022 134192
rect 286966 133728 287022 133784
rect 285954 124208 286010 124264
rect 286230 87216 286286 87272
rect 286230 86944 286286 87000
rect 286046 56616 286102 56672
rect 286230 56616 286286 56672
rect 288346 16904 288402 16960
rect 288346 16768 288402 16824
rect 288714 335280 288770 335336
rect 288990 335280 289046 335336
rect 288714 306348 288716 306368
rect 288716 306348 288768 306368
rect 288768 306348 288770 306368
rect 288714 306312 288770 306348
rect 288898 306312 288954 306368
rect 288806 220768 288862 220824
rect 288714 220632 288770 220688
rect 288714 193196 288716 193216
rect 288716 193196 288768 193216
rect 288768 193196 288770 193216
rect 288714 193160 288770 193196
rect 288898 193196 288900 193216
rect 288900 193196 288952 193216
rect 288952 193196 288954 193216
rect 288898 193160 288954 193196
rect 290186 220804 290188 220824
rect 290188 220804 290240 220824
rect 290240 220804 290242 220824
rect 290186 220768 290242 220804
rect 290186 220632 290242 220688
rect 290002 60696 290058 60752
rect 290186 60696 290242 60752
rect 291658 306312 291714 306368
rect 291842 306312 291898 306368
rect 291382 258032 291438 258088
rect 291566 258052 291622 258088
rect 291566 258032 291568 258052
rect 291568 258032 291620 258052
rect 291620 258032 291622 258052
rect 291474 164192 291530 164248
rect 291658 164192 291714 164248
rect 291842 134000 291898 134056
rect 291842 133728 291898 133784
rect 294234 45464 294290 45520
rect 294142 35944 294198 36000
rect 295706 258052 295762 258088
rect 295706 258032 295708 258052
rect 295708 258032 295760 258052
rect 295760 258032 295762 258052
rect 295890 258032 295946 258088
rect 296626 140800 296682 140856
rect 296534 123256 296590 123312
rect 296534 122984 296590 123040
rect 296810 277380 296812 277400
rect 296812 277380 296864 277400
rect 296864 277380 296866 277400
rect 296810 277344 296866 277380
rect 297086 277344 297142 277400
rect 296810 258032 296866 258088
rect 296994 258032 297050 258088
rect 296810 140800 296866 140856
rect 299386 16768 299442 16824
rect 302606 220768 302662 220824
rect 302514 220632 302570 220688
rect 303986 45736 304042 45792
rect 303802 45600 303858 45656
rect 306010 123020 306012 123040
rect 306012 123020 306064 123040
rect 306064 123020 306066 123040
rect 306010 122984 306066 123020
rect 306378 157548 306434 157584
rect 306378 157528 306380 157548
rect 306380 157528 306432 157548
rect 306432 157528 306434 157548
rect 306286 110780 306288 110800
rect 306288 110780 306340 110800
rect 306340 110780 306342 110800
rect 306286 110744 306342 110780
rect 306286 28908 306288 28928
rect 306288 28908 306340 28928
rect 306340 28908 306342 28928
rect 306286 28872 306342 28908
rect 306654 24792 306710 24848
rect 307022 24792 307078 24848
rect 309046 134036 309048 134056
rect 309048 134036 309100 134056
rect 309100 134036 309102 134056
rect 309046 134000 309102 134036
rect 307390 3304 307446 3360
rect 310426 75792 310482 75848
rect 310426 66272 310482 66328
rect 310794 193160 310850 193216
rect 311070 193160 311126 193216
rect 310886 153312 310942 153368
rect 310794 153196 310850 153232
rect 310794 153176 310796 153196
rect 310796 153176 310848 153196
rect 310848 153176 310850 153196
rect 310794 75792 310850 75848
rect 310794 66272 310850 66328
rect 311162 17040 311218 17096
rect 314566 123256 314622 123312
rect 314566 28908 314568 28928
rect 314568 28908 314620 28928
rect 314620 28908 314622 28928
rect 314566 28872 314622 28908
rect 315946 157392 316002 157448
rect 315946 134136 316002 134192
rect 315946 110780 315948 110800
rect 315948 110780 316000 110800
rect 316000 110780 316002 110800
rect 315946 110744 316002 110780
rect 314658 4800 314714 4856
rect 317418 337728 317474 337784
rect 317326 157664 317382 157720
rect 317326 157392 317382 157448
rect 317326 17040 317382 17096
rect 317326 16632 317382 16688
rect 322202 16768 322258 16824
rect 322202 16360 322258 16416
rect 323306 296656 323362 296712
rect 323490 296656 323546 296712
rect 323398 229064 323454 229120
rect 323582 229064 323638 229120
rect 323398 200062 323454 200118
rect 323398 199824 323454 199880
rect 323306 135224 323362 135280
rect 323490 135224 323546 135280
rect 324502 277344 324558 277400
rect 324778 277344 324834 277400
rect 324594 238720 324650 238776
rect 324778 238720 324834 238776
rect 324686 231820 324688 231840
rect 324688 231820 324740 231840
rect 324740 231820 324742 231840
rect 324686 231784 324742 231820
rect 324778 231648 324834 231704
rect 324594 125568 324650 125624
rect 324778 125568 324834 125624
rect 325606 123528 325662 123584
rect 325606 122984 325662 123040
rect 325606 111016 325662 111072
rect 325606 110744 325662 110800
rect 325606 29144 325662 29200
rect 325606 28872 325662 28928
rect 326986 337728 327042 337784
rect 325882 202852 325884 202872
rect 325884 202852 325936 202872
rect 325936 202852 325938 202872
rect 325882 202816 325938 202852
rect 325974 202680 326030 202736
rect 325882 144900 325938 144936
rect 325882 144880 325884 144900
rect 325884 144880 325936 144900
rect 325936 144880 325938 144900
rect 326066 144900 326122 144936
rect 326066 144880 326068 144900
rect 326068 144880 326120 144900
rect 326120 144880 326122 144900
rect 325882 125568 325938 125624
rect 326066 125568 326122 125624
rect 326986 29280 327042 29336
rect 326986 28872 327042 28928
rect 327170 337748 327226 337784
rect 327170 337728 327172 337748
rect 327172 337728 327224 337748
rect 327224 337728 327226 337748
rect 327170 259392 327226 259448
rect 327354 259256 327410 259312
rect 327262 162832 327318 162888
rect 327446 162832 327502 162888
rect 327170 113328 327226 113384
rect 327170 113192 327226 113248
rect 328458 134136 328514 134192
rect 328458 133864 328514 133920
rect 328458 123120 328514 123176
rect 328458 122984 328514 123040
rect 329930 248376 329986 248432
rect 329930 172508 329986 172544
rect 329930 172488 329932 172508
rect 329932 172488 329984 172508
rect 329984 172488 329986 172508
rect 329930 162832 329986 162888
rect 329930 125568 329986 125624
rect 330298 248376 330354 248432
rect 330206 240080 330262 240136
rect 330390 240080 330446 240136
rect 330298 190440 330354 190496
rect 330482 190440 330538 190496
rect 330114 182144 330170 182200
rect 330298 182144 330354 182200
rect 330206 172508 330262 172544
rect 330206 172488 330208 172508
rect 330208 172488 330260 172508
rect 330260 172488 330262 172508
rect 330114 162832 330170 162888
rect 330114 125588 330170 125624
rect 330114 125568 330116 125588
rect 330116 125568 330168 125588
rect 330168 125568 330170 125588
rect 329930 48184 329986 48240
rect 330298 48320 330354 48376
rect 331126 48184 331182 48240
rect 331402 180784 331458 180840
rect 331586 180784 331642 180840
rect 331494 151816 331550 151872
rect 331678 151816 331734 151872
rect 331862 87352 331918 87408
rect 331862 87080 331918 87136
rect 331402 66136 331458 66192
rect 331586 66000 331642 66056
rect 331586 48320 331642 48376
rect 331494 27784 331550 27840
rect 331402 27648 331458 27704
rect 335174 110744 335230 110800
rect 335174 110608 335230 110664
rect 336186 337748 336242 337784
rect 336186 337728 336188 337748
rect 336188 337728 336240 337748
rect 336240 337728 336242 337748
rect 336738 157548 336794 157584
rect 336738 157528 336740 157548
rect 336740 157528 336792 157548
rect 336792 157528 336794 157548
rect 336738 87100 336794 87136
rect 336738 87080 336740 87100
rect 336740 87080 336792 87100
rect 336792 87080 336794 87100
rect 336646 29280 336702 29336
rect 336646 29008 336702 29064
rect 336646 17040 336702 17096
rect 336646 16632 336702 16688
rect 337198 318960 337254 319016
rect 337106 318824 337162 318880
rect 337106 269048 337162 269104
rect 337290 269048 337346 269104
rect 337106 240080 337162 240136
rect 337290 240080 337346 240136
rect 337106 220768 337162 220824
rect 337290 220768 337346 220824
rect 337198 135360 337254 135416
rect 337198 135244 337254 135280
rect 337198 135224 337200 135244
rect 337200 135224 337252 135244
rect 337252 135224 337254 135244
rect 339774 182144 339830 182200
rect 339958 182144 340014 182200
rect 340878 154536 340934 154592
rect 341246 299376 341302 299432
rect 341246 289856 341302 289912
rect 341246 280064 341302 280120
rect 341246 270544 341302 270600
rect 341246 260752 341302 260808
rect 341246 251232 341302 251288
rect 341154 240080 341210 240136
rect 341430 240080 341486 240136
rect 341154 202852 341156 202872
rect 341156 202852 341208 202872
rect 341208 202852 341210 202872
rect 341154 202816 341210 202852
rect 341430 202816 341486 202872
rect 341338 154536 341394 154592
rect 341154 28872 341210 28928
rect 341338 28872 341394 28928
rect 340878 3032 340934 3088
rect 346306 157392 346362 157448
rect 346306 86944 346362 87000
rect 345754 3032 345810 3088
rect 356242 3304 356298 3360
rect 357438 183504 357494 183560
rect 357622 183504 357678 183560
rect 357622 124072 357678 124128
rect 357806 124072 357862 124128
rect 360106 157528 360162 157584
rect 360290 157528 360346 157584
rect 360106 134000 360162 134056
rect 360290 134000 360346 134056
rect 360106 76064 360162 76120
rect 360290 76064 360346 76120
rect 360106 63688 360162 63744
rect 360290 63688 360346 63744
rect 360106 40160 360162 40216
rect 360290 40160 360346 40216
rect 365626 122984 365682 123040
rect 365626 122848 365682 122904
rect 366822 183504 366878 183560
rect 366730 144880 366786 144936
rect 366730 106256 366786 106312
rect 367006 183540 367008 183560
rect 367008 183540 367060 183560
rect 367060 183540 367062 183560
rect 367006 183504 367062 183540
rect 367006 173848 367062 173904
rect 367006 164212 367062 164248
rect 367006 164192 367008 164212
rect 367008 164192 367060 164212
rect 367060 164192 367062 164212
rect 367006 144900 367062 144936
rect 367006 144880 367008 144900
rect 367008 144880 367060 144900
rect 367060 144880 367062 144900
rect 367006 106276 367062 106312
rect 367006 106256 367008 106276
rect 367008 106256 367060 106276
rect 367060 106256 367062 106276
rect 367006 87216 367062 87272
rect 367006 87080 367062 87136
rect 366914 48456 366970 48512
rect 366914 48320 366970 48376
rect 367098 29144 367154 29200
rect 367098 29008 367154 29064
rect 369674 122848 369730 122904
rect 372526 241440 372582 241496
rect 372710 241440 372766 241496
rect 372526 222128 372582 222184
rect 372710 222128 372766 222184
rect 372526 202816 372582 202872
rect 372710 202816 372766 202872
rect 372526 154536 372582 154592
rect 372710 154536 372766 154592
rect 375838 125588 375894 125624
rect 375838 125568 375840 125588
rect 375840 125568 375892 125588
rect 375892 125568 375894 125588
rect 376942 241440 376998 241496
rect 377126 241440 377182 241496
rect 376942 222128 376998 222184
rect 377126 222128 377182 222184
rect 376942 202816 376998 202872
rect 377126 202816 377182 202872
rect 376942 183504 376998 183560
rect 377126 183504 377182 183560
rect 376114 125568 376170 125624
rect 376666 123120 376722 123176
rect 378230 157700 378232 157720
rect 378232 157700 378284 157720
rect 378284 157700 378286 157720
rect 378230 157664 378286 157700
rect 378230 134172 378232 134192
rect 378232 134172 378284 134192
rect 378284 134172 378286 134192
rect 378230 134136 378286 134172
rect 379058 87100 379114 87136
rect 379058 87080 379060 87100
rect 379060 87080 379112 87100
rect 379112 87080 379114 87100
rect 378230 76236 378232 76256
rect 378232 76236 378284 76256
rect 378284 76236 378286 76256
rect 378230 76200 378286 76236
rect 378230 63860 378232 63880
rect 378232 63860 378284 63880
rect 378284 63860 378286 63880
rect 378230 63824 378286 63860
rect 386326 157700 386328 157720
rect 386328 157700 386380 157720
rect 386380 157700 386382 157720
rect 386326 157664 386382 157700
rect 386326 134172 386328 134192
rect 386328 134172 386380 134192
rect 386380 134172 386382 134192
rect 386326 134136 386382 134172
rect 386326 86944 386382 87000
rect 386326 76236 386328 76256
rect 386328 76236 386380 76256
rect 386380 76236 386382 76256
rect 386326 76200 386382 76236
rect 386326 63860 386328 63880
rect 386328 63860 386380 63880
rect 386380 63860 386382 63880
rect 386326 63824 386382 63860
rect 389270 231784 389326 231840
rect 389454 231784 389510 231840
rect 389270 212472 389326 212528
rect 389454 212472 389510 212528
rect 389270 193160 389326 193216
rect 389454 193160 389510 193216
rect 389362 16496 389418 16552
rect 389546 16496 389602 16552
rect 393594 259392 393650 259448
rect 393778 259392 393834 259448
rect 393318 229064 393374 229120
rect 393502 229064 393558 229120
rect 393318 219408 393374 219464
rect 393502 219408 393558 219464
rect 393318 172488 393374 172544
rect 393594 172488 393650 172544
rect 393594 162968 393650 163024
rect 393686 162852 393742 162888
rect 393686 162832 393688 162852
rect 393688 162832 393740 162852
rect 393740 162832 393742 162852
rect 393594 121624 393650 121680
rect 393594 121488 393650 121544
rect 393502 55120 393558 55176
rect 393686 55120 393742 55176
rect 393410 37304 393466 37360
rect 393594 37304 393650 37360
rect 396078 87100 396134 87136
rect 396078 87080 396080 87100
rect 396080 87080 396132 87100
rect 396132 87080 396134 87100
rect 405554 86944 405610 87000
rect 417882 157548 417938 157584
rect 417882 157528 417884 157548
rect 417884 157528 417936 157548
rect 417936 157528 417938 157548
rect 417882 134020 417938 134056
rect 417882 134000 417884 134020
rect 417884 134000 417936 134020
rect 417936 134000 417938 134020
rect 417882 123004 417938 123040
rect 417882 122984 417884 123004
rect 417884 122984 417936 123004
rect 417936 122984 417938 123004
rect 417882 110628 417938 110664
rect 417882 110608 417884 110628
rect 417884 110608 417936 110628
rect 417936 110608 417938 110628
rect 417882 87116 417884 87136
rect 417884 87116 417936 87136
rect 417936 87116 417938 87136
rect 417882 87080 417938 87116
rect 417882 76084 417938 76120
rect 417882 76064 417884 76084
rect 417884 76064 417936 76084
rect 417936 76064 417938 76084
rect 417882 63708 417938 63744
rect 417882 63688 417884 63708
rect 417884 63688 417936 63708
rect 417936 63688 417938 63708
rect 417882 40180 417938 40216
rect 417882 40160 417884 40180
rect 417884 40160 417936 40180
rect 417936 40160 417938 40180
rect 417882 29164 417938 29200
rect 417882 29144 417884 29164
rect 417884 29144 417936 29164
rect 417936 29144 417938 29164
rect 417882 16788 417938 16824
rect 417882 16768 417884 16788
rect 417884 16768 417936 16788
rect 417936 16768 417938 16788
rect 418158 157548 418214 157584
rect 418158 157528 418160 157548
rect 418160 157528 418212 157548
rect 418212 157528 418214 157548
rect 418158 134020 418214 134056
rect 418158 134000 418160 134020
rect 418160 134000 418212 134020
rect 418212 134000 418214 134020
rect 419354 123004 419410 123040
rect 419354 122984 419356 123004
rect 419356 122984 419408 123004
rect 419408 122984 419410 123004
rect 418158 110628 418214 110664
rect 418158 110608 418160 110628
rect 418160 110608 418212 110628
rect 418212 110608 418214 110628
rect 418618 87116 418620 87136
rect 418620 87116 418672 87136
rect 418672 87116 418674 87136
rect 418618 87080 418674 87116
rect 419354 76084 419410 76120
rect 419354 76064 419356 76084
rect 419356 76064 419408 76084
rect 419408 76064 419410 76084
rect 418158 63708 418214 63744
rect 418158 63688 418160 63708
rect 418160 63688 418212 63708
rect 418212 63688 418214 63708
rect 418158 40180 418214 40216
rect 418158 40160 418160 40180
rect 418160 40160 418212 40180
rect 418212 40160 418214 40180
rect 418158 29164 418214 29200
rect 418158 29144 418160 29164
rect 418160 29144 418212 29164
rect 418212 29144 418214 29164
rect 418158 16788 418214 16824
rect 418158 16768 418160 16788
rect 418160 16768 418212 16788
rect 418212 16768 418214 16788
rect 434718 76100 434720 76120
rect 434720 76100 434772 76120
rect 434772 76100 434774 76120
rect 434718 76064 434774 76100
rect 437202 157548 437258 157584
rect 437202 157528 437204 157548
rect 437204 157528 437256 157548
rect 437256 157528 437258 157548
rect 437202 134036 437204 134056
rect 437204 134036 437256 134056
rect 437256 134036 437258 134056
rect 437202 134000 437258 134036
rect 437202 123004 437258 123040
rect 437202 122984 437204 123004
rect 437204 122984 437256 123004
rect 437256 122984 437258 123004
rect 437202 110628 437258 110664
rect 437202 110608 437204 110628
rect 437204 110608 437256 110628
rect 437256 110608 437258 110628
rect 437202 87100 437258 87136
rect 437202 87080 437204 87100
rect 437204 87080 437256 87100
rect 437256 87080 437258 87100
rect 437202 63708 437258 63744
rect 437202 63688 437204 63708
rect 437204 63688 437256 63708
rect 437256 63688 437258 63708
rect 437202 40196 437204 40216
rect 437204 40196 437256 40216
rect 437256 40196 437258 40216
rect 437202 40160 437258 40196
rect 437202 29180 437204 29200
rect 437204 29180 437256 29200
rect 437256 29180 437258 29200
rect 437202 29144 437258 29180
rect 437202 16788 437258 16824
rect 437202 16768 437204 16788
rect 437204 16768 437256 16788
rect 437256 16768 437258 16788
rect 437478 157548 437534 157584
rect 437478 157528 437480 157548
rect 437480 157528 437532 157548
rect 437532 157528 437534 157548
rect 437570 134036 437572 134056
rect 437572 134036 437624 134056
rect 437624 134036 437626 134056
rect 437570 134000 437626 134036
rect 437478 123004 437534 123040
rect 437478 122984 437480 123004
rect 437480 122984 437532 123004
rect 437532 122984 437534 123004
rect 437478 110628 437534 110664
rect 437478 110608 437480 110628
rect 437480 110608 437532 110628
rect 437532 110608 437534 110628
rect 437478 87100 437534 87136
rect 437478 87080 437480 87100
rect 437480 87080 437532 87100
rect 437532 87080 437534 87100
rect 437478 76100 437480 76120
rect 437480 76100 437532 76120
rect 437532 76100 437534 76120
rect 437478 76064 437534 76100
rect 437478 63708 437534 63744
rect 437478 63688 437480 63708
rect 437480 63688 437532 63708
rect 437532 63688 437534 63708
rect 437570 40196 437572 40216
rect 437572 40196 437624 40216
rect 437624 40196 437626 40216
rect 437570 40160 437626 40196
rect 437478 29180 437480 29200
rect 437480 29180 437532 29200
rect 437532 29180 437534 29200
rect 437478 29144 437534 29180
rect 437478 16788 437534 16824
rect 437478 16768 437480 16788
rect 437480 16768 437532 16788
rect 437532 16768 437534 16788
rect 454038 87216 454094 87272
rect 456522 134156 456578 134192
rect 456522 134136 456524 134156
rect 456524 134136 456576 134156
rect 456576 134136 456578 134156
rect 456522 123140 456578 123176
rect 456522 123120 456524 123140
rect 456524 123120 456576 123140
rect 456576 123120 456578 123140
rect 456522 110764 456578 110800
rect 456522 110744 456524 110764
rect 456524 110744 456576 110764
rect 456576 110744 456578 110764
rect 456522 63708 456578 63744
rect 456522 63688 456524 63708
rect 456524 63688 456576 63708
rect 456576 63688 456578 63708
rect 456522 40196 456524 40216
rect 456524 40196 456576 40216
rect 456576 40196 456578 40216
rect 456522 40160 456578 40196
rect 457442 134000 457498 134056
rect 457442 122984 457498 123040
rect 457442 110608 457498 110664
rect 456890 63708 456946 63744
rect 456890 63688 456892 63708
rect 456892 63688 456944 63708
rect 456944 63688 456946 63708
rect 456890 40196 456892 40216
rect 456892 40196 456944 40216
rect 456944 40196 456946 40216
rect 456890 40160 456946 40196
rect 460018 318824 460074 318880
rect 460202 318824 460258 318880
rect 460018 241476 460020 241496
rect 460020 241476 460072 241496
rect 460072 241476 460074 241496
rect 460018 241440 460074 241476
rect 460110 234504 460166 234560
rect 459834 220768 459890 220824
rect 460018 220768 460074 220824
rect 459926 164192 459982 164248
rect 460202 164192 460258 164248
rect 459926 135224 459982 135280
rect 460110 135224 460166 135280
rect 459926 96600 459982 96656
rect 460110 96600 460166 96656
rect 463422 87168 463478 87170
rect 463422 87116 463424 87168
rect 463424 87116 463476 87168
rect 463476 87116 463478 87168
rect 463422 87114 463478 87116
rect 463790 231784 463846 231840
rect 463974 231784 464030 231840
rect 463790 212472 463846 212528
rect 463974 212472 464030 212528
rect 463790 193160 463846 193216
rect 463974 193160 464030 193216
rect 463882 125568 463938 125624
rect 464066 125568 464122 125624
rect 463698 87116 463700 87136
rect 463700 87116 463752 87136
rect 463752 87116 463754 87136
rect 463698 87080 463754 87116
rect 463698 76100 463700 76120
rect 463700 76100 463752 76120
rect 463752 76100 463754 76120
rect 463698 76064 463754 76100
rect 463790 16668 463792 16688
rect 463792 16668 463844 16688
rect 463844 16668 463846 16688
rect 463790 16632 463846 16668
rect 465262 29180 465264 29200
rect 465264 29180 465316 29200
rect 465316 29180 465318 29200
rect 465262 29144 465318 29180
rect 467562 337320 467618 337376
rect 466550 16904 466606 16960
rect 467930 87216 467986 87272
rect 467930 76200 467986 76256
rect 467930 29280 467986 29336
rect 467746 4800 467802 4856
rect 468850 3304 468906 3360
rect 580170 580760 580226 580816
rect 579802 557232 579858 557288
rect 579802 545536 579858 545592
rect 579802 510312 579858 510368
rect 579802 498616 579858 498672
rect 579802 463392 579858 463448
rect 579894 451696 579950 451752
rect 579894 439864 579950 439920
rect 579894 416472 579950 416528
rect 579894 404776 579950 404832
rect 579894 392944 579950 393000
rect 579986 369552 580042 369608
rect 580078 357856 580134 357912
rect 579802 346024 579858 346080
rect 470506 337184 470562 337240
rect 470690 337184 470746 337240
rect 471886 123120 471942 123176
rect 471886 122712 471942 122768
rect 471886 110744 471942 110800
rect 471886 110336 471942 110392
rect 475566 134036 475568 134056
rect 475568 134036 475620 134056
rect 475620 134036 475622 134056
rect 475566 134000 475622 134036
rect 476026 123120 476082 123176
rect 476210 122984 476266 123040
rect 476026 110744 476082 110800
rect 476210 110608 476266 110664
rect 476026 87216 476082 87272
rect 476210 87080 476266 87136
rect 476026 29280 476082 29336
rect 476210 29144 476266 29200
rect 482926 134036 482928 134056
rect 482928 134036 482980 134056
rect 482980 134036 482982 134056
rect 482926 134000 482982 134036
rect 482926 76472 482982 76528
rect 482926 76064 482982 76120
rect 482926 17176 482982 17232
rect 482926 16768 482982 16824
rect 487802 134272 487858 134328
rect 487802 133864 487858 133920
rect 487802 123256 487858 123312
rect 487802 122848 487858 122904
rect 487802 110880 487858 110936
rect 487802 110472 487858 110528
rect 491206 87352 491262 87408
rect 491206 86944 491262 87000
rect 487802 76336 487858 76392
rect 487802 75928 487858 75984
rect 491206 29416 491262 29472
rect 491206 29008 491262 29064
rect 487802 17040 487858 17096
rect 487802 16632 487858 16688
rect 494610 86944 494666 87000
rect 492770 29044 492772 29064
rect 492772 29044 492824 29064
rect 492824 29044 492826 29064
rect 492770 29008 492826 29044
rect 502246 87216 502302 87272
rect 502246 29280 502302 29336
rect 512642 337320 512698 337376
rect 579986 325624 580042 325680
rect 580078 322632 580134 322688
rect 580170 310800 580226 310856
rect 580078 306348 580080 306368
rect 580080 306348 580132 306368
rect 580132 306348 580134 306368
rect 580078 306312 580134 306348
rect 580170 299104 580226 299160
rect 580170 275712 580226 275768
rect 580906 325660 580908 325680
rect 580908 325660 580960 325680
rect 580960 325660 580962 325680
rect 580906 325624 580962 325660
rect 580906 306348 580908 306368
rect 580908 306348 580960 306368
rect 580960 306348 580962 306368
rect 580906 306312 580962 306348
rect 580814 263880 580870 263936
rect 580722 252184 580778 252240
rect 580630 228792 580686 228848
rect 580538 216960 580594 217016
rect 580446 205264 580502 205320
rect 580354 181872 580410 181928
rect 580262 170040 580318 170096
rect 576214 4800 576270 4856
rect 580998 3304 581054 3360
<< metal3 >>
rect 8109 700362 8175 700365
rect 378133 700362 378199 700365
rect 8109 700360 378199 700362
rect 8109 700304 8114 700360
rect 8170 700304 378138 700360
rect 378194 700304 378199 700360
rect 8109 700302 378199 700304
rect 8109 700299 8175 700302
rect 378133 700299 378199 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect 4797 583402 4863 583405
rect 460289 583402 460355 583405
rect 4797 583400 460355 583402
rect 4797 583344 4802 583400
rect 4858 583344 460294 583400
rect 460350 583344 460355 583400
rect 4797 583342 460355 583344
rect 4797 583339 4863 583342
rect 460289 583339 460355 583342
rect 300301 583266 300367 583269
rect 465758 583266 465764 583268
rect 300301 583264 465764 583266
rect 300301 583208 300306 583264
rect 300362 583208 465764 583264
rect 300301 583206 465764 583208
rect 300301 583203 300367 583206
rect 465758 583204 465764 583206
rect 465828 583204 465834 583268
rect 293953 583130 294019 583133
rect 465574 583130 465580 583132
rect 293953 583128 465580 583130
rect 293953 583072 293958 583128
rect 294014 583072 465580 583128
rect 293953 583070 465580 583072
rect 293953 583067 294019 583070
rect 465574 583068 465580 583070
rect 465644 583068 465650 583132
rect 247902 582932 247908 582996
rect 247972 582994 247978 582996
rect 420269 582994 420335 582997
rect 247972 582992 420335 582994
rect 247972 582936 420274 582992
rect 420330 582936 420335 582992
rect 247972 582934 420335 582936
rect 247972 582932 247978 582934
rect 420269 582931 420335 582934
rect 247718 582796 247724 582860
rect 247788 582858 247794 582860
rect 432965 582858 433031 582861
rect 247788 582856 433031 582858
rect 247788 582800 432970 582856
rect 433026 582800 433031 582856
rect 247788 582798 433031 582800
rect 247788 582796 247794 582798
rect 432965 582795 433031 582798
rect 247534 582660 247540 582724
rect 247604 582722 247610 582724
rect 445569 582722 445635 582725
rect 247604 582720 445635 582722
rect 247604 582664 445574 582720
rect 445630 582664 445635 582720
rect 247604 582662 445635 582664
rect 247604 582660 247610 582662
rect 445569 582659 445635 582662
rect 31017 582586 31083 582589
rect 462405 582586 462471 582589
rect 31017 582584 462471 582586
rect 31017 582528 31022 582584
rect 31078 582528 462410 582584
rect 462466 582528 462471 582584
rect 31017 582526 462471 582528
rect 31017 582523 31083 582526
rect 462405 582523 462471 582526
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 231117 579322 231183 579325
rect 232957 579324 233023 579325
rect 231710 579322 231716 579324
rect 231117 579320 231716 579322
rect 231117 579264 231122 579320
rect 231178 579264 231716 579320
rect 231117 579262 231716 579264
rect 231117 579259 231183 579262
rect 231710 579260 231716 579262
rect 231780 579260 231786 579324
rect 232957 579320 233004 579324
rect 233068 579322 233074 579324
rect 235257 579322 235323 579325
rect 237189 579324 237255 579325
rect 235758 579322 235764 579324
rect 232957 579264 232962 579320
rect 232957 579260 233004 579264
rect 233068 579262 233114 579322
rect 235257 579320 235764 579322
rect 235257 579264 235262 579320
rect 235318 579264 235764 579320
rect 235257 579262 235764 579264
rect 233068 579260 233074 579262
rect 232957 579259 233023 579260
rect 235257 579259 235323 579262
rect 235758 579260 235764 579262
rect 235828 579260 235834 579324
rect 237189 579320 237236 579324
rect 237300 579322 237306 579324
rect 239397 579322 239463 579325
rect 239990 579322 239996 579324
rect 237189 579264 237194 579320
rect 237189 579260 237236 579264
rect 237300 579262 237346 579322
rect 239397 579320 239996 579322
rect 239397 579264 239402 579320
rect 239458 579264 239996 579320
rect 239397 579262 239996 579264
rect 237300 579260 237306 579262
rect 237189 579259 237255 579260
rect 239397 579259 239463 579262
rect 239990 579260 239996 579262
rect 240060 579260 240066 579324
rect 241278 579260 241284 579324
rect 241348 579322 241354 579324
rect 241421 579322 241487 579325
rect 241348 579320 241487 579322
rect 241348 579264 241426 579320
rect 241482 579264 241487 579320
rect 241348 579262 241487 579264
rect 241348 579260 241354 579262
rect 241421 579259 241487 579262
rect 243629 579322 243695 579325
rect 245377 579324 245443 579325
rect 244038 579322 244044 579324
rect 243629 579320 244044 579322
rect 243629 579264 243634 579320
rect 243690 579264 244044 579320
rect 243629 579262 244044 579264
rect 243629 579259 243695 579262
rect 244038 579260 244044 579262
rect 244108 579260 244114 579324
rect 245326 579322 245332 579324
rect 245286 579262 245332 579322
rect 245396 579320 245443 579324
rect 245438 579264 245443 579320
rect 245326 579260 245332 579262
rect 245396 579260 245443 579264
rect 245377 579259 245443 579260
rect 247861 579322 247927 579325
rect 248270 579322 248276 579324
rect 247861 579320 248276 579322
rect 247861 579264 247866 579320
rect 247922 579264 248276 579320
rect 247861 579262 248276 579264
rect 247861 579259 247927 579262
rect 248270 579260 248276 579262
rect 248340 579260 248346 579324
rect 249006 579260 249012 579324
rect 249076 579322 249082 579324
rect 249517 579322 249583 579325
rect 249076 579320 249583 579322
rect 249076 579264 249522 579320
rect 249578 579264 249583 579320
rect 249076 579262 249583 579264
rect 249076 579260 249082 579262
rect 249517 579259 249583 579262
rect 466453 579324 466519 579325
rect 466453 579320 466500 579324
rect 466564 579322 466570 579324
rect 466453 579264 466458 579320
rect 466453 579260 466500 579264
rect 466564 579262 466610 579322
rect 466564 579260 466570 579262
rect 467782 579260 467788 579324
rect 467852 579322 467858 579324
rect 468569 579322 468635 579325
rect 467852 579320 468635 579322
rect 467852 579264 468574 579320
rect 468630 579264 468635 579320
rect 467852 579262 468635 579264
rect 467852 579260 467858 579262
rect 466453 579259 466519 579260
rect 468569 579259 468635 579262
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3141 567354 3207 567357
rect -960 567352 3207 567354
rect -960 567296 3146 567352
rect 3202 567296 3207 567352
rect -960 567294 3207 567296
rect -960 567204 480 567294
rect 3141 567291 3207 567294
rect 579797 557290 579863 557293
rect 583520 557290 584960 557380
rect 579797 557288 584960 557290
rect 579797 557232 579802 557288
rect 579858 557232 584960 557288
rect 579797 557230 584960 557232
rect 579797 557227 579863 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 579797 545594 579863 545597
rect 583520 545594 584960 545684
rect 579797 545592 584960 545594
rect 579797 545536 579802 545592
rect 579858 545536 584960 545592
rect 579797 545534 584960 545536
rect 579797 545531 579863 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3049 538658 3115 538661
rect -960 538656 3115 538658
rect -960 538600 3054 538656
rect 3110 538600 3115 538656
rect -960 538598 3115 538600
rect -960 538508 480 538598
rect 3049 538595 3115 538598
rect 583520 533898 584960 533988
rect 583342 533838 584960 533898
rect 465758 533020 465764 533084
rect 465828 533082 465834 533084
rect 465828 533022 470610 533082
rect 465828 533020 465834 533022
rect 470550 532946 470610 533022
rect 480302 533022 489930 533082
rect 470550 532886 480178 532946
rect 480118 532810 480178 532886
rect 480302 532810 480362 533022
rect 489870 532946 489930 533022
rect 499622 533022 509250 533082
rect 489870 532886 499498 532946
rect 480118 532750 480362 532810
rect 499438 532810 499498 532886
rect 499622 532810 499682 533022
rect 509190 532946 509250 533022
rect 518942 533022 528570 533082
rect 509190 532886 518818 532946
rect 499438 532750 499682 532810
rect 518758 532810 518818 532886
rect 518942 532810 519002 533022
rect 528510 532946 528570 533022
rect 538262 533022 547890 533082
rect 528510 532886 538138 532946
rect 518758 532750 519002 532810
rect 538078 532810 538138 532886
rect 538262 532810 538322 533022
rect 547830 532946 547890 533022
rect 557582 533022 567210 533082
rect 547830 532886 557458 532946
rect 538078 532750 538322 532810
rect 557398 532810 557458 532886
rect 557582 532810 557642 533022
rect 567150 532946 567210 533022
rect 583342 532946 583402 533838
rect 583520 533748 584960 533838
rect 567150 532886 576778 532946
rect 557398 532750 557642 532810
rect 576718 532810 576778 532886
rect 576902 532886 583402 532946
rect 576902 532810 576962 532886
rect 576718 532750 576962 532810
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 579797 510370 579863 510373
rect 583520 510370 584960 510460
rect 579797 510368 584960 510370
rect 579797 510312 579802 510368
rect 579858 510312 584960 510368
rect 579797 510310 584960 510312
rect 579797 510307 579863 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3141 509962 3207 509965
rect -960 509960 3207 509962
rect -960 509904 3146 509960
rect 3202 509904 3207 509960
rect -960 509902 3207 509904
rect -960 509812 480 509902
rect 3141 509899 3207 509902
rect 579797 498674 579863 498677
rect 583520 498674 584960 498764
rect 579797 498672 584960 498674
rect 579797 498616 579802 498672
rect 579858 498616 584960 498672
rect 579797 498614 584960 498616
rect 579797 498611 579863 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 2773 495546 2839 495549
rect -960 495544 2839 495546
rect -960 495488 2778 495544
rect 2834 495488 2839 495544
rect -960 495486 2839 495488
rect -960 495396 480 495486
rect 2773 495483 2839 495486
rect 583520 486842 584960 486932
rect 583342 486782 584960 486842
rect 465942 486100 465948 486164
rect 466012 486162 466018 486164
rect 466012 486102 470610 486162
rect 466012 486100 466018 486102
rect 470550 486026 470610 486102
rect 480302 486102 489930 486162
rect 470550 485966 480178 486026
rect 480118 485890 480178 485966
rect 480302 485890 480362 486102
rect 489870 486026 489930 486102
rect 499622 486102 509250 486162
rect 489870 485966 499498 486026
rect 480118 485830 480362 485890
rect 499438 485890 499498 485966
rect 499622 485890 499682 486102
rect 509190 486026 509250 486102
rect 518942 486102 528570 486162
rect 509190 485966 518818 486026
rect 499438 485830 499682 485890
rect 518758 485890 518818 485966
rect 518942 485890 519002 486102
rect 528510 486026 528570 486102
rect 538262 486102 547890 486162
rect 528510 485966 538138 486026
rect 518758 485830 519002 485890
rect 538078 485890 538138 485966
rect 538262 485890 538322 486102
rect 547830 486026 547890 486102
rect 557582 486102 567210 486162
rect 547830 485966 557458 486026
rect 538078 485830 538322 485890
rect 557398 485890 557458 485966
rect 557582 485890 557642 486102
rect 567150 486026 567210 486102
rect 583342 486026 583402 486782
rect 583520 486692 584960 486782
rect 567150 485966 576778 486026
rect 557398 485830 557642 485890
rect 576718 485890 576778 485966
rect 576902 485966 583402 486026
rect 576902 485890 576962 485966
rect 576718 485830 576962 485890
rect -960 481130 480 481220
rect 3141 481130 3207 481133
rect -960 481128 3207 481130
rect -960 481072 3146 481128
rect 3202 481072 3207 481128
rect -960 481070 3207 481072
rect -960 480980 480 481070
rect 3141 481067 3207 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 579797 463450 579863 463453
rect 583520 463450 584960 463540
rect 579797 463448 584960 463450
rect 579797 463392 579802 463448
rect 579858 463392 584960 463448
rect 579797 463390 584960 463392
rect 579797 463387 579863 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 3233 452434 3299 452437
rect -960 452432 3299 452434
rect -960 452376 3238 452432
rect 3294 452376 3299 452432
rect -960 452374 3299 452376
rect -960 452284 480 452374
rect 3233 452371 3299 452374
rect 579889 451754 579955 451757
rect 583520 451754 584960 451844
rect 579889 451752 584960 451754
rect 579889 451696 579894 451752
rect 579950 451696 584960 451752
rect 579889 451694 584960 451696
rect 579889 451691 579955 451694
rect 583520 451604 584960 451694
rect 579889 439922 579955 439925
rect 583520 439922 584960 440012
rect 579889 439920 584960 439922
rect 579889 439864 579894 439920
rect 579950 439864 584960 439920
rect 579889 439862 584960 439864
rect 579889 439859 579955 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 2773 438018 2839 438021
rect -960 438016 2839 438018
rect -960 437960 2778 438016
rect 2834 437960 2839 438016
rect -960 437958 2839 437960
rect -960 437868 480 437958
rect 2773 437955 2839 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 2773 423738 2839 423741
rect -960 423736 2839 423738
rect -960 423680 2778 423736
rect 2834 423680 2839 423736
rect -960 423678 2839 423680
rect -960 423588 480 423678
rect 2773 423675 2839 423678
rect 579889 416530 579955 416533
rect 583520 416530 584960 416620
rect 579889 416528 584960 416530
rect 579889 416472 579894 416528
rect 579950 416472 584960 416528
rect 579889 416470 584960 416472
rect 579889 416467 579955 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 579889 404834 579955 404837
rect 583520 404834 584960 404924
rect 579889 404832 584960 404834
rect 579889 404776 579894 404832
rect 579950 404776 584960 404832
rect 579889 404774 584960 404776
rect 579889 404771 579955 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3233 395042 3299 395045
rect -960 395040 3299 395042
rect -960 394984 3238 395040
rect 3294 394984 3299 395040
rect -960 394982 3299 394984
rect -960 394892 480 394982
rect 3233 394979 3299 394982
rect 579889 393002 579955 393005
rect 583520 393002 584960 393092
rect 579889 393000 584960 393002
rect 579889 392944 579894 393000
rect 579950 392944 584960 393000
rect 579889 392942 584960 392944
rect 579889 392939 579955 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 2773 380626 2839 380629
rect -960 380624 2839 380626
rect -960 380568 2778 380624
rect 2834 380568 2839 380624
rect -960 380566 2839 380568
rect -960 380476 480 380566
rect 2773 380563 2839 380566
rect 579981 369610 580047 369613
rect 583520 369610 584960 369700
rect 579981 369608 584960 369610
rect 579981 369552 579986 369608
rect 580042 369552 584960 369608
rect 579981 369550 584960 369552
rect 579981 369547 580047 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3325 366210 3391 366213
rect -960 366208 3391 366210
rect -960 366152 3330 366208
rect 3386 366152 3391 366208
rect -960 366150 3391 366152
rect -960 366060 480 366150
rect 3325 366147 3391 366150
rect 580073 357914 580139 357917
rect 583520 357914 584960 358004
rect 580073 357912 584960 357914
rect 580073 357856 580078 357912
rect 580134 357856 584960 357912
rect 580073 357854 584960 357856
rect 580073 357851 580139 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579797 346082 579863 346085
rect 583520 346082 584960 346172
rect 579797 346080 584960 346082
rect 579797 346024 579802 346080
rect 579858 346024 584960 346080
rect 579797 346022 584960 346024
rect 579797 346019 579863 346022
rect 583520 345932 584960 346022
rect 247902 338058 247908 338060
rect 614 337998 247908 338058
rect -960 337514 480 337604
rect 614 337514 674 337998
rect 247902 337996 247908 337998
rect 247972 337996 247978 338060
rect 317413 337786 317479 337789
rect 326981 337786 327047 337789
rect 317413 337784 327047 337786
rect 317413 337728 317418 337784
rect 317474 337728 326986 337784
rect 327042 337728 327047 337784
rect 317413 337726 327047 337728
rect 317413 337723 317479 337726
rect 326981 337723 327047 337726
rect 327165 337786 327231 337789
rect 336181 337786 336247 337789
rect 327165 337784 336247 337786
rect 327165 337728 327170 337784
rect 327226 337728 336186 337784
rect 336242 337728 336247 337784
rect 327165 337726 336247 337728
rect 327165 337723 327231 337726
rect 336181 337723 336247 337726
rect -960 337454 674 337514
rect -960 337364 480 337454
rect 10317 337378 10383 337381
rect 231945 337378 232011 337381
rect 10317 337376 232011 337378
rect 10317 337320 10322 337376
rect 10378 337320 231950 337376
rect 232006 337320 232011 337376
rect 10317 337318 232011 337320
rect 10317 337315 10383 337318
rect 231945 337315 232011 337318
rect 467557 337378 467623 337381
rect 512637 337378 512703 337381
rect 467557 337376 512703 337378
rect 467557 337320 467562 337376
rect 467618 337320 512642 337376
rect 512698 337320 512703 337376
rect 467557 337318 512703 337320
rect 467557 337315 467623 337318
rect 512637 337315 512703 337318
rect 132493 337242 132559 337245
rect 142061 337242 142127 337245
rect 132493 337240 142127 337242
rect 132493 337184 132498 337240
rect 132554 337184 142066 337240
rect 142122 337184 142127 337240
rect 132493 337182 142127 337184
rect 132493 337179 132559 337182
rect 142061 337179 142127 337182
rect 151813 337242 151879 337245
rect 161381 337242 161447 337245
rect 151813 337240 161447 337242
rect 151813 337184 151818 337240
rect 151874 337184 161386 337240
rect 161442 337184 161447 337240
rect 151813 337182 161447 337184
rect 151813 337179 151879 337182
rect 161381 337179 161447 337182
rect 171133 337242 171199 337245
rect 180701 337242 180767 337245
rect 171133 337240 180767 337242
rect 171133 337184 171138 337240
rect 171194 337184 180706 337240
rect 180762 337184 180767 337240
rect 171133 337182 180767 337184
rect 171133 337179 171199 337182
rect 180701 337179 180767 337182
rect 190453 337242 190519 337245
rect 200021 337242 200087 337245
rect 190453 337240 200087 337242
rect 190453 337184 190458 337240
rect 190514 337184 200026 337240
rect 200082 337184 200087 337240
rect 190453 337182 200087 337184
rect 190453 337179 190519 337182
rect 200021 337179 200087 337182
rect 209773 337242 209839 337245
rect 219341 337242 219407 337245
rect 209773 337240 219407 337242
rect 209773 337184 209778 337240
rect 209834 337184 219346 337240
rect 219402 337184 219407 337240
rect 209773 337182 219407 337184
rect 209773 337179 209839 337182
rect 219341 337179 219407 337182
rect 229185 337242 229251 337245
rect 234613 337242 234679 337245
rect 229185 337240 234679 337242
rect 229185 337184 229190 337240
rect 229246 337184 234618 337240
rect 234674 337184 234679 337240
rect 229185 337182 234679 337184
rect 229185 337179 229251 337182
rect 234613 337179 234679 337182
rect 470501 337242 470567 337245
rect 470685 337242 470751 337245
rect 470501 337240 470751 337242
rect 470501 337184 470506 337240
rect 470562 337184 470690 337240
rect 470746 337184 470751 337240
rect 470501 337182 470751 337184
rect 470501 337179 470567 337182
rect 470685 337179 470751 337182
rect 288709 335338 288775 335341
rect 288985 335338 289051 335341
rect 288709 335336 289051 335338
rect 288709 335280 288714 335336
rect 288770 335280 288990 335336
rect 289046 335280 289051 335336
rect 288709 335278 289051 335280
rect 288709 335275 288775 335278
rect 288985 335275 289051 335278
rect 583520 334236 584960 334476
rect 285765 325682 285831 325685
rect 285949 325682 286015 325685
rect 285765 325680 286015 325682
rect 285765 325624 285770 325680
rect 285826 325624 285954 325680
rect 286010 325624 286015 325680
rect 285765 325622 286015 325624
rect 285765 325619 285831 325622
rect 285949 325619 286015 325622
rect 579981 325682 580047 325685
rect 580901 325682 580967 325685
rect 579981 325680 580967 325682
rect 579981 325624 579986 325680
rect 580042 325624 580906 325680
rect 580962 325624 580967 325680
rect 579981 325622 580967 325624
rect 579981 325619 580047 325622
rect 580901 325619 580967 325622
rect -960 323098 480 323188
rect 3325 323098 3391 323101
rect -960 323096 3391 323098
rect -960 323040 3330 323096
rect 3386 323040 3391 323096
rect -960 323038 3391 323040
rect -960 322948 480 323038
rect 3325 323035 3391 323038
rect 580073 322690 580139 322693
rect 583520 322690 584960 322780
rect 580073 322688 584960 322690
rect 580073 322632 580078 322688
rect 580134 322632 584960 322688
rect 580073 322630 584960 322632
rect 580073 322627 580139 322630
rect 583520 322540 584960 322630
rect 337193 319018 337259 319021
rect 336966 319016 337259 319018
rect 336966 318960 337198 319016
rect 337254 318960 337259 319016
rect 336966 318958 337259 318960
rect 336966 318882 337026 318958
rect 337193 318955 337259 318958
rect 337101 318882 337167 318885
rect 336966 318880 337167 318882
rect 336966 318824 337106 318880
rect 337162 318824 337167 318880
rect 336966 318822 337167 318824
rect 337101 318819 337167 318822
rect 460013 318882 460079 318885
rect 460197 318882 460263 318885
rect 460013 318880 460263 318882
rect 460013 318824 460018 318880
rect 460074 318824 460202 318880
rect 460258 318824 460263 318880
rect 460013 318822 460263 318824
rect 460013 318819 460079 318822
rect 460197 318819 460263 318822
rect 286041 316026 286107 316029
rect 286225 316026 286291 316029
rect 286041 316024 286291 316026
rect 286041 315968 286046 316024
rect 286102 315968 286230 316024
rect 286286 315968 286291 316024
rect 286041 315966 286291 315968
rect 286041 315963 286107 315966
rect 286225 315963 286291 315966
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 4061 308818 4127 308821
rect -960 308816 4127 308818
rect -960 308760 4066 308816
rect 4122 308760 4127 308816
rect -960 308758 4127 308760
rect -960 308668 480 308758
rect 4061 308755 4127 308758
rect 251398 307668 251404 307732
rect 251468 307730 251474 307732
rect 251541 307730 251607 307733
rect 251468 307728 251607 307730
rect 251468 307672 251546 307728
rect 251602 307672 251607 307728
rect 251468 307670 251607 307672
rect 251468 307668 251474 307670
rect 251541 307667 251607 307670
rect 267825 306370 267891 306373
rect 268009 306370 268075 306373
rect 267825 306368 268075 306370
rect 267825 306312 267830 306368
rect 267886 306312 268014 306368
rect 268070 306312 268075 306368
rect 267825 306310 268075 306312
rect 267825 306307 267891 306310
rect 268009 306307 268075 306310
rect 288709 306370 288775 306373
rect 288893 306370 288959 306373
rect 288709 306368 288959 306370
rect 288709 306312 288714 306368
rect 288770 306312 288898 306368
rect 288954 306312 288959 306368
rect 288709 306310 288959 306312
rect 288709 306307 288775 306310
rect 288893 306307 288959 306310
rect 291653 306370 291719 306373
rect 291837 306370 291903 306373
rect 291653 306368 291903 306370
rect 291653 306312 291658 306368
rect 291714 306312 291842 306368
rect 291898 306312 291903 306368
rect 291653 306310 291903 306312
rect 291653 306307 291719 306310
rect 291837 306307 291903 306310
rect 580073 306370 580139 306373
rect 580901 306370 580967 306373
rect 580073 306368 580967 306370
rect 580073 306312 580078 306368
rect 580134 306312 580906 306368
rect 580962 306312 580967 306368
rect 580073 306310 580967 306312
rect 580073 306307 580139 306310
rect 580901 306307 580967 306310
rect 341241 299434 341307 299437
rect 341374 299434 341380 299436
rect 341241 299432 341380 299434
rect 341241 299376 341246 299432
rect 341302 299376 341380 299432
rect 341241 299374 341380 299376
rect 341241 299371 341307 299374
rect 341374 299372 341380 299374
rect 341444 299372 341450 299436
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect 251398 298148 251404 298212
rect 251468 298210 251474 298212
rect 251541 298210 251607 298213
rect 251468 298208 251607 298210
rect 251468 298152 251546 298208
rect 251602 298152 251607 298208
rect 251468 298150 251607 298152
rect 251468 298148 251474 298150
rect 251541 298147 251607 298150
rect 323301 296714 323367 296717
rect 323485 296714 323551 296717
rect 323301 296712 323551 296714
rect 323301 296656 323306 296712
rect 323362 296656 323490 296712
rect 323546 296656 323551 296712
rect 323301 296654 323551 296656
rect 323301 296651 323367 296654
rect 323485 296651 323551 296654
rect -960 294402 480 294492
rect 3969 294402 4035 294405
rect -960 294400 4035 294402
rect -960 294344 3974 294400
rect 4030 294344 4035 294400
rect -960 294342 4035 294344
rect -960 294252 480 294342
rect 3969 294339 4035 294342
rect 341241 289914 341307 289917
rect 341374 289914 341380 289916
rect 341241 289912 341380 289914
rect 341241 289856 341246 289912
rect 341302 289856 341380 289912
rect 341241 289854 341380 289856
rect 341241 289851 341307 289854
rect 341374 289852 341380 289854
rect 341444 289852 341450 289916
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3325 280122 3391 280125
rect -960 280120 3391 280122
rect -960 280064 3330 280120
rect 3386 280064 3391 280120
rect -960 280062 3391 280064
rect -960 279972 480 280062
rect 3325 280059 3391 280062
rect 251173 280122 251239 280125
rect 251357 280122 251423 280125
rect 251173 280120 251423 280122
rect 251173 280064 251178 280120
rect 251234 280064 251362 280120
rect 251418 280064 251423 280120
rect 251173 280062 251423 280064
rect 251173 280059 251239 280062
rect 251357 280059 251423 280062
rect 341241 280122 341307 280125
rect 341374 280122 341380 280124
rect 341241 280120 341380 280122
rect 341241 280064 341246 280120
rect 341302 280064 341380 280120
rect 341241 280062 341380 280064
rect 341241 280059 341307 280062
rect 341374 280060 341380 280062
rect 341444 280060 341450 280124
rect 245929 278762 245995 278765
rect 246113 278762 246179 278765
rect 245929 278760 246179 278762
rect 245929 278704 245934 278760
rect 245990 278704 246118 278760
rect 246174 278704 246179 278760
rect 245929 278702 246179 278704
rect 245929 278699 245995 278702
rect 246113 278699 246179 278702
rect 272149 278762 272215 278765
rect 272333 278762 272399 278765
rect 281717 278762 281783 278765
rect 272149 278760 272399 278762
rect 272149 278704 272154 278760
rect 272210 278704 272338 278760
rect 272394 278704 272399 278760
rect 272149 278702 272399 278704
rect 272149 278699 272215 278702
rect 272333 278699 272399 278702
rect 281582 278760 281783 278762
rect 281582 278704 281722 278760
rect 281778 278704 281783 278760
rect 281582 278702 281783 278704
rect 281582 278626 281642 278702
rect 281717 278699 281783 278702
rect 284661 278762 284727 278765
rect 284845 278762 284911 278765
rect 284661 278760 284911 278762
rect 284661 278704 284666 278760
rect 284722 278704 284850 278760
rect 284906 278704 284911 278760
rect 284661 278702 284911 278704
rect 284661 278699 284727 278702
rect 284845 278699 284911 278702
rect 281809 278626 281875 278629
rect 281582 278624 281875 278626
rect 281582 278568 281814 278624
rect 281870 278568 281875 278624
rect 281582 278566 281875 278568
rect 281809 278563 281875 278566
rect 296805 277402 296871 277405
rect 297081 277402 297147 277405
rect 296805 277400 297147 277402
rect 296805 277344 296810 277400
rect 296866 277344 297086 277400
rect 297142 277344 297147 277400
rect 296805 277342 297147 277344
rect 296805 277339 296871 277342
rect 297081 277339 297147 277342
rect 324497 277402 324563 277405
rect 324773 277402 324839 277405
rect 324497 277400 324839 277402
rect 324497 277344 324502 277400
rect 324558 277344 324778 277400
rect 324834 277344 324839 277400
rect 324497 277342 324839 277344
rect 324497 277339 324563 277342
rect 324773 277339 324839 277342
rect 265249 276042 265315 276045
rect 265525 276042 265591 276045
rect 265249 276040 265591 276042
rect 265249 275984 265254 276040
rect 265310 275984 265530 276040
rect 265586 275984 265591 276040
rect 265249 275982 265591 275984
rect 265249 275979 265315 275982
rect 265525 275979 265591 275982
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 341241 270602 341307 270605
rect 341374 270602 341380 270604
rect 341241 270600 341380 270602
rect 341241 270544 341246 270600
rect 341302 270544 341380 270600
rect 341241 270542 341380 270544
rect 341241 270539 341307 270542
rect 341374 270540 341380 270542
rect 341444 270540 341450 270604
rect 262581 269106 262647 269109
rect 267733 269106 267799 269109
rect 337101 269106 337167 269109
rect 337285 269106 337351 269109
rect 262581 269104 262690 269106
rect 262581 269048 262586 269104
rect 262642 269048 262690 269104
rect 262581 269043 262690 269048
rect 267733 269104 267842 269106
rect 267733 269048 267738 269104
rect 267794 269048 267842 269104
rect 267733 269043 267842 269048
rect 337101 269104 337351 269106
rect 337101 269048 337106 269104
rect 337162 269048 337290 269104
rect 337346 269048 337351 269104
rect 337101 269046 337351 269048
rect 337101 269043 337167 269046
rect 337285 269043 337351 269046
rect 262630 268973 262690 269043
rect 267782 268973 267842 269043
rect 262630 268968 262739 268973
rect 262630 268912 262678 268968
rect 262734 268912 262739 268968
rect 262630 268910 262739 268912
rect 267782 268968 267891 268973
rect 267782 268912 267830 268968
rect 267886 268912 267891 268968
rect 267782 268910 267891 268912
rect 262673 268907 262739 268910
rect 267825 268907 267891 268910
rect 265157 266386 265223 266389
rect 265341 266386 265407 266389
rect 265157 266384 265407 266386
rect 265157 266328 265162 266384
rect 265218 266328 265346 266384
rect 265402 266328 265407 266384
rect 265157 266326 265407 266328
rect 265157 266323 265223 266326
rect 265341 266323 265407 266326
rect -960 265706 480 265796
rect 3877 265706 3943 265709
rect -960 265704 3943 265706
rect -960 265648 3882 265704
rect 3938 265648 3943 265704
rect -960 265646 3943 265648
rect -960 265556 480 265646
rect 3877 265643 3943 265646
rect 580809 263938 580875 263941
rect 583520 263938 584960 264028
rect 580809 263936 584960 263938
rect 580809 263880 580814 263936
rect 580870 263880 584960 263936
rect 580809 263878 584960 263880
rect 580809 263875 580875 263878
rect 583520 263788 584960 263878
rect 251173 260810 251239 260813
rect 251357 260810 251423 260813
rect 251173 260808 251423 260810
rect 251173 260752 251178 260808
rect 251234 260752 251362 260808
rect 251418 260752 251423 260808
rect 251173 260750 251423 260752
rect 251173 260747 251239 260750
rect 251357 260747 251423 260750
rect 341241 260810 341307 260813
rect 341374 260810 341380 260812
rect 341241 260808 341380 260810
rect 341241 260752 341246 260808
rect 341302 260752 341380 260808
rect 341241 260750 341380 260752
rect 341241 260747 341307 260750
rect 341374 260748 341380 260750
rect 341444 260748 341450 260812
rect 245837 259450 245903 259453
rect 246021 259450 246087 259453
rect 327165 259450 327231 259453
rect 245837 259448 246087 259450
rect 245837 259392 245842 259448
rect 245898 259392 246026 259448
rect 246082 259392 246087 259448
rect 245837 259390 246087 259392
rect 245837 259387 245903 259390
rect 246021 259387 246087 259390
rect 327030 259448 327231 259450
rect 327030 259392 327170 259448
rect 327226 259392 327231 259448
rect 327030 259390 327231 259392
rect 327030 259314 327090 259390
rect 327165 259387 327231 259390
rect 393589 259450 393655 259453
rect 393773 259450 393839 259453
rect 393589 259448 393839 259450
rect 393589 259392 393594 259448
rect 393650 259392 393778 259448
rect 393834 259392 393839 259448
rect 393589 259390 393839 259392
rect 393589 259387 393655 259390
rect 393773 259387 393839 259390
rect 327349 259314 327415 259317
rect 327030 259312 327415 259314
rect 327030 259256 327354 259312
rect 327410 259256 327415 259312
rect 327030 259254 327415 259256
rect 327349 259251 327415 259254
rect 291377 258090 291443 258093
rect 291561 258090 291627 258093
rect 291377 258088 291627 258090
rect 291377 258032 291382 258088
rect 291438 258032 291566 258088
rect 291622 258032 291627 258088
rect 291377 258030 291627 258032
rect 291377 258027 291443 258030
rect 291561 258027 291627 258030
rect 295701 258090 295767 258093
rect 295885 258090 295951 258093
rect 295701 258088 295951 258090
rect 295701 258032 295706 258088
rect 295762 258032 295890 258088
rect 295946 258032 295951 258088
rect 295701 258030 295951 258032
rect 295701 258027 295767 258030
rect 295885 258027 295951 258030
rect 296805 258090 296871 258093
rect 296989 258090 297055 258093
rect 296805 258088 297055 258090
rect 296805 258032 296810 258088
rect 296866 258032 296994 258088
rect 297050 258032 297055 258088
rect 296805 258030 297055 258032
rect 296805 258027 296871 258030
rect 296989 258027 297055 258030
rect 3141 252514 3207 252517
rect 247718 252514 247724 252516
rect 3141 252512 247724 252514
rect 3141 252456 3146 252512
rect 3202 252456 247724 252512
rect 3141 252454 247724 252456
rect 3141 252451 3207 252454
rect 247718 252452 247724 252454
rect 247788 252452 247794 252516
rect 580717 252242 580783 252245
rect 583520 252242 584960 252332
rect 580717 252240 584960 252242
rect 580717 252184 580722 252240
rect 580778 252184 584960 252240
rect 580717 252182 584960 252184
rect 580717 252179 580783 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3141 251290 3207 251293
rect -960 251288 3207 251290
rect -960 251232 3146 251288
rect 3202 251232 3207 251288
rect -960 251230 3207 251232
rect -960 251140 480 251230
rect 3141 251227 3207 251230
rect 341241 251290 341307 251293
rect 341374 251290 341380 251292
rect 341241 251288 341380 251290
rect 341241 251232 341246 251288
rect 341302 251232 341380 251288
rect 341241 251230 341380 251232
rect 341241 251227 341307 251230
rect 341374 251228 341380 251230
rect 341444 251228 341450 251292
rect 244365 249794 244431 249797
rect 244549 249794 244615 249797
rect 244365 249792 244615 249794
rect 244365 249736 244370 249792
rect 244426 249736 244554 249792
rect 244610 249736 244615 249792
rect 244365 249734 244615 249736
rect 244365 249731 244431 249734
rect 244549 249731 244615 249734
rect 245837 249794 245903 249797
rect 246113 249794 246179 249797
rect 245837 249792 246179 249794
rect 245837 249736 245842 249792
rect 245898 249736 246118 249792
rect 246174 249736 246179 249792
rect 245837 249734 246179 249736
rect 245837 249731 245903 249734
rect 246113 249731 246179 249734
rect 251173 249794 251239 249797
rect 251449 249794 251515 249797
rect 251173 249792 251515 249794
rect 251173 249736 251178 249792
rect 251234 249736 251454 249792
rect 251510 249736 251515 249792
rect 251173 249734 251515 249736
rect 251173 249731 251239 249734
rect 251449 249731 251515 249734
rect 262305 248434 262371 248437
rect 262489 248434 262555 248437
rect 262305 248432 262555 248434
rect 262305 248376 262310 248432
rect 262366 248376 262494 248432
rect 262550 248376 262555 248432
rect 262305 248374 262555 248376
rect 262305 248371 262371 248374
rect 262489 248371 262555 248374
rect 329925 248434 329991 248437
rect 330293 248434 330359 248437
rect 329925 248432 330359 248434
rect 329925 248376 329930 248432
rect 329986 248376 330298 248432
rect 330354 248376 330359 248432
rect 329925 248374 330359 248376
rect 329925 248371 329991 248374
rect 330293 248371 330359 248374
rect 234889 241498 234955 241501
rect 235073 241498 235139 241501
rect 234889 241496 235139 241498
rect 234889 241440 234894 241496
rect 234950 241440 235078 241496
rect 235134 241440 235139 241496
rect 234889 241438 235139 241440
rect 234889 241435 234955 241438
rect 235073 241435 235139 241438
rect 236269 241498 236335 241501
rect 236453 241498 236519 241501
rect 236269 241496 236519 241498
rect 236269 241440 236274 241496
rect 236330 241440 236458 241496
rect 236514 241440 236519 241496
rect 236269 241438 236519 241440
rect 236269 241435 236335 241438
rect 236453 241435 236519 241438
rect 273529 241498 273595 241501
rect 273713 241498 273779 241501
rect 273529 241496 273779 241498
rect 273529 241440 273534 241496
rect 273590 241440 273718 241496
rect 273774 241440 273779 241496
rect 273529 241438 273779 241440
rect 273529 241435 273595 241438
rect 273713 241435 273779 241438
rect 372521 241498 372587 241501
rect 372705 241498 372771 241501
rect 372521 241496 372771 241498
rect 372521 241440 372526 241496
rect 372582 241440 372710 241496
rect 372766 241440 372771 241496
rect 372521 241438 372771 241440
rect 372521 241435 372587 241438
rect 372705 241435 372771 241438
rect 376937 241498 377003 241501
rect 377121 241498 377187 241501
rect 376937 241496 377187 241498
rect 376937 241440 376942 241496
rect 376998 241440 377126 241496
rect 377182 241440 377187 241496
rect 376937 241438 377187 241440
rect 376937 241435 377003 241438
rect 377121 241435 377187 241438
rect 460013 241500 460079 241501
rect 460013 241496 460060 241500
rect 460124 241498 460130 241500
rect 460013 241440 460018 241496
rect 460013 241436 460060 241440
rect 460124 241438 460170 241498
rect 460124 241436 460130 241438
rect 460013 241435 460079 241436
rect 583520 240396 584960 240636
rect 251081 240138 251147 240141
rect 251357 240138 251423 240141
rect 251081 240136 251423 240138
rect 251081 240080 251086 240136
rect 251142 240080 251362 240136
rect 251418 240080 251423 240136
rect 251081 240078 251423 240080
rect 251081 240075 251147 240078
rect 251357 240075 251423 240078
rect 272149 240138 272215 240141
rect 272333 240138 272399 240141
rect 272149 240136 272399 240138
rect 272149 240080 272154 240136
rect 272210 240080 272338 240136
rect 272394 240080 272399 240136
rect 272149 240078 272399 240080
rect 272149 240075 272215 240078
rect 272333 240075 272399 240078
rect 330201 240138 330267 240141
rect 330385 240138 330451 240141
rect 330201 240136 330451 240138
rect 330201 240080 330206 240136
rect 330262 240080 330390 240136
rect 330446 240080 330451 240136
rect 330201 240078 330451 240080
rect 330201 240075 330267 240078
rect 330385 240075 330451 240078
rect 337101 240138 337167 240141
rect 337285 240138 337351 240141
rect 337101 240136 337351 240138
rect 337101 240080 337106 240136
rect 337162 240080 337290 240136
rect 337346 240080 337351 240136
rect 337101 240078 337351 240080
rect 337101 240075 337167 240078
rect 337285 240075 337351 240078
rect 341149 240138 341215 240141
rect 341425 240138 341491 240141
rect 341149 240136 341491 240138
rect 341149 240080 341154 240136
rect 341210 240080 341430 240136
rect 341486 240080 341491 240136
rect 341149 240078 341491 240080
rect 341149 240075 341215 240078
rect 341425 240075 341491 240078
rect 286041 238914 286107 238917
rect 285998 238912 286107 238914
rect 285998 238856 286046 238912
rect 286102 238856 286107 238912
rect 285998 238851 286107 238856
rect 285998 238781 286058 238851
rect 285949 238776 286058 238781
rect 285949 238720 285954 238776
rect 286010 238720 286058 238776
rect 285949 238718 286058 238720
rect 324589 238778 324655 238781
rect 324773 238778 324839 238781
rect 324589 238776 324839 238778
rect 324589 238720 324594 238776
rect 324650 238720 324778 238776
rect 324834 238720 324839 238776
rect 324589 238718 324839 238720
rect 285949 238715 286015 238718
rect 324589 238715 324655 238718
rect 324773 238715 324839 238718
rect -960 237010 480 237100
rect 3325 237010 3391 237013
rect -960 237008 3391 237010
rect -960 236952 3330 237008
rect 3386 236952 3391 237008
rect -960 236950 3391 236952
rect -960 236860 480 236950
rect 3325 236947 3391 236950
rect 460105 234564 460171 234565
rect 460054 234562 460060 234564
rect 460014 234502 460060 234562
rect 460124 234560 460171 234564
rect 460166 234504 460171 234560
rect 460054 234500 460060 234502
rect 460124 234500 460171 234504
rect 460105 234499 460171 234500
rect 324681 231842 324747 231845
rect 324638 231840 324747 231842
rect 324638 231784 324686 231840
rect 324742 231784 324747 231840
rect 324638 231779 324747 231784
rect 389265 231842 389331 231845
rect 389449 231842 389515 231845
rect 389265 231840 389515 231842
rect 389265 231784 389270 231840
rect 389326 231784 389454 231840
rect 389510 231784 389515 231840
rect 389265 231782 389515 231784
rect 389265 231779 389331 231782
rect 389449 231779 389515 231782
rect 463785 231842 463851 231845
rect 463969 231842 464035 231845
rect 463785 231840 464035 231842
rect 463785 231784 463790 231840
rect 463846 231784 463974 231840
rect 464030 231784 464035 231840
rect 463785 231782 464035 231784
rect 463785 231779 463851 231782
rect 463969 231779 464035 231782
rect 324638 231706 324698 231779
rect 324773 231706 324839 231709
rect 324638 231704 324839 231706
rect 324638 231648 324778 231704
rect 324834 231648 324839 231704
rect 324638 231646 324839 231648
rect 324773 231643 324839 231646
rect 251357 230482 251423 230485
rect 251541 230482 251607 230485
rect 251357 230480 251607 230482
rect 251357 230424 251362 230480
rect 251418 230424 251546 230480
rect 251602 230424 251607 230480
rect 251357 230422 251607 230424
rect 251357 230419 251423 230422
rect 251541 230419 251607 230422
rect 323393 229122 323459 229125
rect 323577 229122 323643 229125
rect 323393 229120 323643 229122
rect 323393 229064 323398 229120
rect 323454 229064 323582 229120
rect 323638 229064 323643 229120
rect 323393 229062 323643 229064
rect 323393 229059 323459 229062
rect 323577 229059 323643 229062
rect 393313 229122 393379 229125
rect 393497 229122 393563 229125
rect 393313 229120 393563 229122
rect 393313 229064 393318 229120
rect 393374 229064 393502 229120
rect 393558 229064 393563 229120
rect 393313 229062 393563 229064
rect 393313 229059 393379 229062
rect 393497 229059 393563 229062
rect 580625 228850 580691 228853
rect 583520 228850 584960 228940
rect 580625 228848 584960 228850
rect 580625 228792 580630 228848
rect 580686 228792 584960 228848
rect 580625 228790 584960 228792
rect 580625 228787 580691 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 2773 222594 2839 222597
rect -960 222592 2839 222594
rect -960 222536 2778 222592
rect 2834 222536 2839 222592
rect -960 222534 2839 222536
rect -960 222444 480 222534
rect 2773 222531 2839 222534
rect 234889 222186 234955 222189
rect 235073 222186 235139 222189
rect 234889 222184 235139 222186
rect 234889 222128 234894 222184
rect 234950 222128 235078 222184
rect 235134 222128 235139 222184
rect 234889 222126 235139 222128
rect 234889 222123 234955 222126
rect 235073 222123 235139 222126
rect 236269 222186 236335 222189
rect 236453 222186 236519 222189
rect 259637 222186 259703 222189
rect 236269 222184 236519 222186
rect 236269 222128 236274 222184
rect 236330 222128 236458 222184
rect 236514 222128 236519 222184
rect 236269 222126 236519 222128
rect 236269 222123 236335 222126
rect 236453 222123 236519 222126
rect 259502 222184 259703 222186
rect 259502 222128 259642 222184
rect 259698 222128 259703 222184
rect 259502 222126 259703 222128
rect 259502 221914 259562 222126
rect 259637 222123 259703 222126
rect 265157 222186 265223 222189
rect 265341 222186 265407 222189
rect 265157 222184 265407 222186
rect 265157 222128 265162 222184
rect 265218 222128 265346 222184
rect 265402 222128 265407 222184
rect 265157 222126 265407 222128
rect 265157 222123 265223 222126
rect 265341 222123 265407 222126
rect 267733 222186 267799 222189
rect 273529 222186 273595 222189
rect 273713 222186 273779 222189
rect 267733 222184 267842 222186
rect 267733 222128 267738 222184
rect 267794 222128 267842 222184
rect 267733 222123 267842 222128
rect 273529 222184 273779 222186
rect 273529 222128 273534 222184
rect 273590 222128 273718 222184
rect 273774 222128 273779 222184
rect 273529 222126 273779 222128
rect 273529 222123 273595 222126
rect 273713 222123 273779 222126
rect 372521 222186 372587 222189
rect 372705 222186 372771 222189
rect 372521 222184 372771 222186
rect 372521 222128 372526 222184
rect 372582 222128 372710 222184
rect 372766 222128 372771 222184
rect 372521 222126 372771 222128
rect 372521 222123 372587 222126
rect 372705 222123 372771 222126
rect 376937 222186 377003 222189
rect 377121 222186 377187 222189
rect 376937 222184 377187 222186
rect 376937 222128 376942 222184
rect 376998 222128 377126 222184
rect 377182 222128 377187 222184
rect 376937 222126 377187 222128
rect 376937 222123 377003 222126
rect 377121 222123 377187 222126
rect 267782 222053 267842 222123
rect 267733 222048 267842 222053
rect 267733 221992 267738 222048
rect 267794 221992 267842 222048
rect 267733 221990 267842 221992
rect 267733 221987 267799 221990
rect 259729 221914 259795 221917
rect 259502 221912 259795 221914
rect 259502 221856 259734 221912
rect 259790 221856 259795 221912
rect 259502 221854 259795 221856
rect 259729 221851 259795 221854
rect 247166 220764 247172 220828
rect 247236 220826 247242 220828
rect 247309 220826 247375 220829
rect 247236 220824 247375 220826
rect 247236 220768 247314 220824
rect 247370 220768 247375 220824
rect 247236 220766 247375 220768
rect 247236 220764 247242 220766
rect 247309 220763 247375 220766
rect 266629 220826 266695 220829
rect 266813 220826 266879 220829
rect 266629 220824 266879 220826
rect 266629 220768 266634 220824
rect 266690 220768 266818 220824
rect 266874 220768 266879 220824
rect 266629 220766 266879 220768
rect 266629 220763 266695 220766
rect 266813 220763 266879 220766
rect 272057 220826 272123 220829
rect 272241 220826 272307 220829
rect 288801 220826 288867 220829
rect 272057 220824 272307 220826
rect 272057 220768 272062 220824
rect 272118 220768 272246 220824
rect 272302 220768 272307 220824
rect 272057 220766 272307 220768
rect 272057 220763 272123 220766
rect 272241 220763 272307 220766
rect 288758 220824 288867 220826
rect 288758 220768 288806 220824
rect 288862 220768 288867 220824
rect 288758 220763 288867 220768
rect 290181 220826 290247 220829
rect 302601 220826 302667 220829
rect 290181 220824 290290 220826
rect 290181 220768 290186 220824
rect 290242 220768 290290 220824
rect 290181 220763 290290 220768
rect 288758 220693 288818 220763
rect 290230 220693 290290 220763
rect 302558 220824 302667 220826
rect 302558 220768 302606 220824
rect 302662 220768 302667 220824
rect 302558 220763 302667 220768
rect 337101 220826 337167 220829
rect 337285 220826 337351 220829
rect 337101 220824 337351 220826
rect 337101 220768 337106 220824
rect 337162 220768 337290 220824
rect 337346 220768 337351 220824
rect 337101 220766 337351 220768
rect 337101 220763 337167 220766
rect 337285 220763 337351 220766
rect 459829 220826 459895 220829
rect 460013 220826 460079 220829
rect 459829 220824 460079 220826
rect 459829 220768 459834 220824
rect 459890 220768 460018 220824
rect 460074 220768 460079 220824
rect 459829 220766 460079 220768
rect 459829 220763 459895 220766
rect 460013 220763 460079 220766
rect 302558 220693 302618 220763
rect 288709 220688 288818 220693
rect 288709 220632 288714 220688
rect 288770 220632 288818 220688
rect 288709 220630 288818 220632
rect 290181 220688 290290 220693
rect 290181 220632 290186 220688
rect 290242 220632 290290 220688
rect 290181 220630 290290 220632
rect 302509 220688 302618 220693
rect 302509 220632 302514 220688
rect 302570 220632 302618 220688
rect 302509 220630 302618 220632
rect 288709 220627 288775 220630
rect 290181 220627 290247 220630
rect 302509 220627 302575 220630
rect 393313 219466 393379 219469
rect 393497 219466 393563 219469
rect 393313 219464 393563 219466
rect 393313 219408 393318 219464
rect 393374 219408 393502 219464
rect 393558 219408 393563 219464
rect 393313 219406 393563 219408
rect 393313 219403 393379 219406
rect 393497 219403 393563 219406
rect 580533 217018 580599 217021
rect 583520 217018 584960 217108
rect 580533 217016 584960 217018
rect 580533 216960 580538 217016
rect 580594 216960 584960 217016
rect 580533 216958 584960 216960
rect 580533 216955 580599 216958
rect 583520 216868 584960 216958
rect 270493 212530 270559 212533
rect 270769 212530 270835 212533
rect 270493 212528 270835 212530
rect 270493 212472 270498 212528
rect 270554 212472 270774 212528
rect 270830 212472 270835 212528
rect 270493 212470 270835 212472
rect 270493 212467 270559 212470
rect 270769 212467 270835 212470
rect 389265 212530 389331 212533
rect 389449 212530 389515 212533
rect 389265 212528 389515 212530
rect 389265 212472 389270 212528
rect 389326 212472 389454 212528
rect 389510 212472 389515 212528
rect 389265 212470 389515 212472
rect 389265 212467 389331 212470
rect 389449 212467 389515 212470
rect 463785 212530 463851 212533
rect 463969 212530 464035 212533
rect 463785 212528 464035 212530
rect 463785 212472 463790 212528
rect 463846 212472 463974 212528
rect 464030 212472 464035 212528
rect 463785 212470 464035 212472
rect 463785 212467 463851 212470
rect 463969 212467 464035 212470
rect 247217 211172 247283 211173
rect 247166 211108 247172 211172
rect 247236 211170 247283 211172
rect 272057 211170 272123 211173
rect 272241 211170 272307 211173
rect 247236 211168 247328 211170
rect 247278 211112 247328 211168
rect 247236 211110 247328 211112
rect 272057 211168 272307 211170
rect 272057 211112 272062 211168
rect 272118 211112 272246 211168
rect 272302 211112 272307 211168
rect 272057 211110 272307 211112
rect 247236 211108 247283 211110
rect 247217 211107 247283 211108
rect 272057 211107 272123 211110
rect 272241 211107 272307 211110
rect -960 208178 480 208268
rect 3785 208178 3851 208181
rect -960 208176 3851 208178
rect -960 208120 3790 208176
rect 3846 208120 3851 208176
rect -960 208118 3851 208120
rect -960 208028 480 208118
rect 3785 208115 3851 208118
rect 580441 205322 580507 205325
rect 583520 205322 584960 205412
rect 580441 205320 584960 205322
rect 580441 205264 580446 205320
rect 580502 205264 584960 205320
rect 580441 205262 584960 205264
rect 580441 205259 580507 205262
rect 583520 205172 584960 205262
rect 230749 202874 230815 202877
rect 231025 202874 231091 202877
rect 230749 202872 231091 202874
rect 230749 202816 230754 202872
rect 230810 202816 231030 202872
rect 231086 202816 231091 202872
rect 230749 202814 231091 202816
rect 230749 202811 230815 202814
rect 231025 202811 231091 202814
rect 236269 202874 236335 202877
rect 236453 202874 236519 202877
rect 236269 202872 236519 202874
rect 236269 202816 236274 202872
rect 236330 202816 236458 202872
rect 236514 202816 236519 202872
rect 236269 202814 236519 202816
rect 236269 202811 236335 202814
rect 236453 202811 236519 202814
rect 259637 202874 259703 202877
rect 259913 202874 259979 202877
rect 259637 202872 259979 202874
rect 259637 202816 259642 202872
rect 259698 202816 259918 202872
rect 259974 202816 259979 202872
rect 259637 202814 259979 202816
rect 259637 202811 259703 202814
rect 259913 202811 259979 202814
rect 262581 202874 262647 202877
rect 265157 202874 265223 202877
rect 265341 202874 265407 202877
rect 262581 202872 262690 202874
rect 262581 202816 262586 202872
rect 262642 202816 262690 202872
rect 262581 202811 262690 202816
rect 265157 202872 265407 202874
rect 265157 202816 265162 202872
rect 265218 202816 265346 202872
rect 265402 202816 265407 202872
rect 265157 202814 265407 202816
rect 265157 202811 265223 202814
rect 265341 202811 265407 202814
rect 267733 202874 267799 202877
rect 267917 202874 267983 202877
rect 267733 202872 267983 202874
rect 267733 202816 267738 202872
rect 267794 202816 267922 202872
rect 267978 202816 267983 202872
rect 267733 202814 267983 202816
rect 267733 202811 267799 202814
rect 267917 202811 267983 202814
rect 270493 202874 270559 202877
rect 270677 202874 270743 202877
rect 272149 202874 272215 202877
rect 270493 202872 270743 202874
rect 270493 202816 270498 202872
rect 270554 202816 270682 202872
rect 270738 202816 270743 202872
rect 270493 202814 270743 202816
rect 270493 202811 270559 202814
rect 270677 202811 270743 202814
rect 272014 202872 272215 202874
rect 272014 202816 272154 202872
rect 272210 202816 272215 202872
rect 272014 202814 272215 202816
rect 262630 202741 262690 202811
rect 262630 202736 262739 202741
rect 262630 202680 262678 202736
rect 262734 202680 262739 202736
rect 262630 202678 262739 202680
rect 272014 202738 272074 202814
rect 272149 202811 272215 202814
rect 273529 202874 273595 202877
rect 273713 202874 273779 202877
rect 273529 202872 273779 202874
rect 273529 202816 273534 202872
rect 273590 202816 273718 202872
rect 273774 202816 273779 202872
rect 273529 202814 273779 202816
rect 273529 202811 273595 202814
rect 273713 202811 273779 202814
rect 325877 202874 325943 202877
rect 341149 202874 341215 202877
rect 341425 202874 341491 202877
rect 325877 202872 325986 202874
rect 325877 202816 325882 202872
rect 325938 202816 325986 202872
rect 325877 202811 325986 202816
rect 341149 202872 341491 202874
rect 341149 202816 341154 202872
rect 341210 202816 341430 202872
rect 341486 202816 341491 202872
rect 341149 202814 341491 202816
rect 341149 202811 341215 202814
rect 341425 202811 341491 202814
rect 372521 202874 372587 202877
rect 372705 202874 372771 202877
rect 372521 202872 372771 202874
rect 372521 202816 372526 202872
rect 372582 202816 372710 202872
rect 372766 202816 372771 202872
rect 372521 202814 372771 202816
rect 372521 202811 372587 202814
rect 372705 202811 372771 202814
rect 376937 202874 377003 202877
rect 377121 202874 377187 202877
rect 376937 202872 377187 202874
rect 376937 202816 376942 202872
rect 376998 202816 377126 202872
rect 377182 202816 377187 202872
rect 376937 202814 377187 202816
rect 376937 202811 377003 202814
rect 377121 202811 377187 202814
rect 325926 202741 325986 202811
rect 272333 202738 272399 202741
rect 272014 202736 272399 202738
rect 272014 202680 272338 202736
rect 272394 202680 272399 202736
rect 272014 202678 272399 202680
rect 325926 202736 326035 202741
rect 325926 202680 325974 202736
rect 326030 202680 326035 202736
rect 325926 202678 326035 202680
rect 262673 202675 262739 202678
rect 272333 202675 272399 202678
rect 325969 202675 326035 202678
rect 246941 201514 247007 201517
rect 247125 201514 247191 201517
rect 246941 201512 247191 201514
rect 246941 201456 246946 201512
rect 247002 201456 247130 201512
rect 247186 201456 247191 201512
rect 246941 201454 247191 201456
rect 246941 201451 247007 201454
rect 247125 201451 247191 201454
rect 249977 201514 250043 201517
rect 250161 201514 250227 201517
rect 249977 201512 250227 201514
rect 249977 201456 249982 201512
rect 250038 201456 250166 201512
rect 250222 201456 250227 201512
rect 249977 201454 250227 201456
rect 249977 201451 250043 201454
rect 250161 201451 250227 201454
rect 323393 200120 323459 200123
rect 323393 200118 323594 200120
rect 323393 200062 323398 200118
rect 323454 200062 323594 200118
rect 323393 200060 323594 200062
rect 323393 200057 323459 200060
rect 323393 199882 323459 199885
rect 323534 199882 323594 200060
rect 323393 199880 323594 199882
rect 323393 199824 323398 199880
rect 323454 199824 323594 199880
rect 323393 199822 323594 199824
rect 323393 199819 323459 199822
rect -960 193898 480 193988
rect 3693 193898 3759 193901
rect -960 193896 3759 193898
rect -960 193840 3698 193896
rect 3754 193840 3759 193896
rect -960 193838 3759 193840
rect -960 193748 480 193838
rect 3693 193835 3759 193838
rect 583520 193476 584960 193716
rect 251357 193218 251423 193221
rect 251541 193218 251607 193221
rect 251357 193216 251607 193218
rect 251357 193160 251362 193216
rect 251418 193160 251546 193216
rect 251602 193160 251607 193216
rect 251357 193158 251607 193160
rect 251357 193155 251423 193158
rect 251541 193155 251607 193158
rect 264973 193218 265039 193221
rect 265249 193218 265315 193221
rect 264973 193216 265315 193218
rect 264973 193160 264978 193216
rect 265034 193160 265254 193216
rect 265310 193160 265315 193216
rect 264973 193158 265315 193160
rect 264973 193155 265039 193158
rect 265249 193155 265315 193158
rect 270493 193218 270559 193221
rect 270769 193218 270835 193221
rect 270493 193216 270835 193218
rect 270493 193160 270498 193216
rect 270554 193160 270774 193216
rect 270830 193160 270835 193216
rect 270493 193158 270835 193160
rect 270493 193155 270559 193158
rect 270769 193155 270835 193158
rect 281717 193218 281783 193221
rect 281901 193218 281967 193221
rect 281717 193216 281967 193218
rect 281717 193160 281722 193216
rect 281778 193160 281906 193216
rect 281962 193160 281967 193216
rect 281717 193158 281967 193160
rect 281717 193155 281783 193158
rect 281901 193155 281967 193158
rect 284661 193218 284727 193221
rect 284845 193218 284911 193221
rect 284661 193216 284911 193218
rect 284661 193160 284666 193216
rect 284722 193160 284850 193216
rect 284906 193160 284911 193216
rect 284661 193158 284911 193160
rect 284661 193155 284727 193158
rect 284845 193155 284911 193158
rect 288709 193218 288775 193221
rect 288893 193218 288959 193221
rect 288709 193216 288959 193218
rect 288709 193160 288714 193216
rect 288770 193160 288898 193216
rect 288954 193160 288959 193216
rect 288709 193158 288959 193160
rect 288709 193155 288775 193158
rect 288893 193155 288959 193158
rect 310789 193218 310855 193221
rect 311065 193218 311131 193221
rect 310789 193216 311131 193218
rect 310789 193160 310794 193216
rect 310850 193160 311070 193216
rect 311126 193160 311131 193216
rect 310789 193158 311131 193160
rect 310789 193155 310855 193158
rect 311065 193155 311131 193158
rect 389265 193218 389331 193221
rect 389449 193218 389515 193221
rect 389265 193216 389515 193218
rect 389265 193160 389270 193216
rect 389326 193160 389454 193216
rect 389510 193160 389515 193216
rect 389265 193158 389515 193160
rect 389265 193155 389331 193158
rect 389449 193155 389515 193158
rect 463785 193218 463851 193221
rect 463969 193218 464035 193221
rect 463785 193216 464035 193218
rect 463785 193160 463790 193216
rect 463846 193160 463974 193216
rect 464030 193160 464035 193216
rect 463785 193158 464035 193160
rect 463785 193155 463851 193158
rect 463969 193155 464035 193158
rect 330293 190498 330359 190501
rect 330477 190498 330543 190501
rect 330293 190496 330543 190498
rect 330293 190440 330298 190496
rect 330354 190440 330482 190496
rect 330538 190440 330543 190496
rect 330293 190438 330543 190440
rect 330293 190435 330359 190438
rect 330477 190435 330543 190438
rect 230749 183562 230815 183565
rect 231025 183562 231091 183565
rect 230749 183560 231091 183562
rect 230749 183504 230754 183560
rect 230810 183504 231030 183560
rect 231086 183504 231091 183560
rect 230749 183502 231091 183504
rect 230749 183499 230815 183502
rect 231025 183499 231091 183502
rect 236269 183562 236335 183565
rect 236453 183562 236519 183565
rect 236269 183560 236519 183562
rect 236269 183504 236274 183560
rect 236330 183504 236458 183560
rect 236514 183504 236519 183560
rect 236269 183502 236519 183504
rect 236269 183499 236335 183502
rect 236453 183499 236519 183502
rect 259637 183562 259703 183565
rect 259913 183562 259979 183565
rect 259637 183560 259979 183562
rect 259637 183504 259642 183560
rect 259698 183504 259918 183560
rect 259974 183504 259979 183560
rect 259637 183502 259979 183504
rect 259637 183499 259703 183502
rect 259913 183499 259979 183502
rect 262581 183562 262647 183565
rect 265157 183562 265223 183565
rect 265341 183562 265407 183565
rect 262581 183560 262690 183562
rect 262581 183504 262586 183560
rect 262642 183504 262690 183560
rect 262581 183499 262690 183504
rect 265157 183560 265407 183562
rect 265157 183504 265162 183560
rect 265218 183504 265346 183560
rect 265402 183504 265407 183560
rect 265157 183502 265407 183504
rect 265157 183499 265223 183502
rect 265341 183499 265407 183502
rect 270493 183562 270559 183565
rect 270677 183562 270743 183565
rect 272149 183562 272215 183565
rect 270493 183560 270743 183562
rect 270493 183504 270498 183560
rect 270554 183504 270682 183560
rect 270738 183504 270743 183560
rect 270493 183502 270743 183504
rect 270493 183499 270559 183502
rect 270677 183499 270743 183502
rect 272014 183560 272215 183562
rect 272014 183504 272154 183560
rect 272210 183504 272215 183560
rect 272014 183502 272215 183504
rect 262630 183429 262690 183499
rect 262630 183424 262739 183429
rect 262630 183368 262678 183424
rect 262734 183368 262739 183424
rect 262630 183366 262739 183368
rect 272014 183426 272074 183502
rect 272149 183499 272215 183502
rect 273529 183562 273595 183565
rect 273713 183562 273779 183565
rect 273529 183560 273779 183562
rect 273529 183504 273534 183560
rect 273590 183504 273718 183560
rect 273774 183504 273779 183560
rect 273529 183502 273779 183504
rect 273529 183499 273595 183502
rect 273713 183499 273779 183502
rect 357433 183562 357499 183565
rect 357617 183562 357683 183565
rect 357433 183560 357683 183562
rect 357433 183504 357438 183560
rect 357494 183504 357622 183560
rect 357678 183504 357683 183560
rect 357433 183502 357683 183504
rect 357433 183499 357499 183502
rect 357617 183499 357683 183502
rect 366817 183562 366883 183565
rect 367001 183562 367067 183565
rect 366817 183560 367067 183562
rect 366817 183504 366822 183560
rect 366878 183504 367006 183560
rect 367062 183504 367067 183560
rect 366817 183502 367067 183504
rect 366817 183499 366883 183502
rect 367001 183499 367067 183502
rect 376937 183562 377003 183565
rect 377121 183562 377187 183565
rect 376937 183560 377187 183562
rect 376937 183504 376942 183560
rect 376998 183504 377126 183560
rect 377182 183504 377187 183560
rect 376937 183502 377187 183504
rect 376937 183499 377003 183502
rect 377121 183499 377187 183502
rect 272333 183426 272399 183429
rect 272014 183424 272399 183426
rect 272014 183368 272338 183424
rect 272394 183368 272399 183424
rect 272014 183366 272399 183368
rect 262673 183363 262739 183366
rect 272333 183363 272399 183366
rect 285949 182202 286015 182205
rect 286133 182202 286199 182205
rect 285949 182200 286199 182202
rect 285949 182144 285954 182200
rect 286010 182144 286138 182200
rect 286194 182144 286199 182200
rect 285949 182142 286199 182144
rect 285949 182139 286015 182142
rect 286133 182139 286199 182142
rect 330109 182202 330175 182205
rect 330293 182202 330359 182205
rect 330109 182200 330359 182202
rect 330109 182144 330114 182200
rect 330170 182144 330298 182200
rect 330354 182144 330359 182200
rect 330109 182142 330359 182144
rect 330109 182139 330175 182142
rect 330293 182139 330359 182142
rect 339769 182202 339835 182205
rect 339953 182202 340019 182205
rect 339769 182200 340019 182202
rect 339769 182144 339774 182200
rect 339830 182144 339958 182200
rect 340014 182144 340019 182200
rect 339769 182142 340019 182144
rect 339769 182139 339835 182142
rect 339953 182139 340019 182142
rect 580349 181930 580415 181933
rect 583520 181930 584960 182020
rect 580349 181928 584960 181930
rect 580349 181872 580354 181928
rect 580410 181872 584960 181928
rect 580349 181870 584960 181872
rect 580349 181867 580415 181870
rect 583520 181780 584960 181870
rect 267733 180842 267799 180845
rect 267917 180842 267983 180845
rect 267733 180840 267983 180842
rect 267733 180784 267738 180840
rect 267794 180784 267922 180840
rect 267978 180784 267983 180840
rect 267733 180782 267983 180784
rect 267733 180779 267799 180782
rect 267917 180779 267983 180782
rect 331397 180842 331463 180845
rect 331581 180842 331647 180845
rect 331397 180840 331647 180842
rect 331397 180784 331402 180840
rect 331458 180784 331586 180840
rect 331642 180784 331647 180840
rect 331397 180782 331647 180784
rect 331397 180779 331463 180782
rect 331581 180779 331647 180782
rect -960 179482 480 179572
rect 3601 179482 3667 179485
rect -960 179480 3667 179482
rect -960 179424 3606 179480
rect 3662 179424 3667 179480
rect -960 179422 3667 179424
rect -960 179332 480 179422
rect 3601 179419 3667 179422
rect 281717 173906 281783 173909
rect 281901 173906 281967 173909
rect 281717 173904 281967 173906
rect 281717 173848 281722 173904
rect 281778 173848 281906 173904
rect 281962 173848 281967 173904
rect 281717 173846 281967 173848
rect 281717 173843 281783 173846
rect 281901 173843 281967 173846
rect 284661 173906 284727 173909
rect 284845 173906 284911 173909
rect 284661 173904 284911 173906
rect 284661 173848 284666 173904
rect 284722 173848 284850 173904
rect 284906 173848 284911 173904
rect 284661 173846 284911 173848
rect 284661 173843 284727 173846
rect 284845 173843 284911 173846
rect 285949 173906 286015 173909
rect 286133 173906 286199 173909
rect 367001 173908 367067 173909
rect 366950 173906 366956 173908
rect 285949 173904 286199 173906
rect 285949 173848 285954 173904
rect 286010 173848 286138 173904
rect 286194 173848 286199 173904
rect 285949 173846 286199 173848
rect 366910 173846 366956 173906
rect 367020 173904 367067 173908
rect 367062 173848 367067 173904
rect 285949 173843 286015 173846
rect 286133 173843 286199 173846
rect 366950 173844 366956 173846
rect 367020 173844 367067 173848
rect 367001 173843 367067 173844
rect 272057 172546 272123 172549
rect 272241 172546 272307 172549
rect 272057 172544 272307 172546
rect 272057 172488 272062 172544
rect 272118 172488 272246 172544
rect 272302 172488 272307 172544
rect 272057 172486 272307 172488
rect 272057 172483 272123 172486
rect 272241 172483 272307 172486
rect 329925 172546 329991 172549
rect 330201 172546 330267 172549
rect 329925 172544 330267 172546
rect 329925 172488 329930 172544
rect 329986 172488 330206 172544
rect 330262 172488 330267 172544
rect 329925 172486 330267 172488
rect 329925 172483 329991 172486
rect 330201 172483 330267 172486
rect 393313 172546 393379 172549
rect 393589 172546 393655 172549
rect 393313 172544 393655 172546
rect 393313 172488 393318 172544
rect 393374 172488 393594 172544
rect 393650 172488 393655 172544
rect 393313 172486 393655 172488
rect 393313 172483 393379 172486
rect 393589 172483 393655 172486
rect 580257 170098 580323 170101
rect 583520 170098 584960 170188
rect 580257 170096 584960 170098
rect 580257 170040 580262 170096
rect 580318 170040 584960 170096
rect 580257 170038 584960 170040
rect 580257 170035 580323 170038
rect 583520 169948 584960 170038
rect 247534 165610 247540 165612
rect 614 165550 247540 165610
rect -960 165066 480 165156
rect 614 165066 674 165550
rect 247534 165548 247540 165550
rect 247604 165548 247610 165612
rect -960 165006 674 165066
rect -960 164916 480 165006
rect 291469 164250 291535 164253
rect 291653 164250 291719 164253
rect 367001 164252 367067 164253
rect 366950 164250 366956 164252
rect 291469 164248 291719 164250
rect 291469 164192 291474 164248
rect 291530 164192 291658 164248
rect 291714 164192 291719 164248
rect 291469 164190 291719 164192
rect 366910 164190 366956 164250
rect 367020 164248 367067 164252
rect 367062 164192 367067 164248
rect 291469 164187 291535 164190
rect 291653 164187 291719 164190
rect 366950 164188 366956 164190
rect 367020 164188 367067 164192
rect 367001 164187 367067 164188
rect 459921 164250 459987 164253
rect 460197 164250 460263 164253
rect 459921 164248 460263 164250
rect 459921 164192 459926 164248
rect 459982 164192 460202 164248
rect 460258 164192 460263 164248
rect 459921 164190 460263 164192
rect 459921 164187 459987 164190
rect 460197 164187 460263 164190
rect 393589 163026 393655 163029
rect 393589 163024 393698 163026
rect 393589 162968 393594 163024
rect 393650 162968 393698 163024
rect 393589 162963 393698 162968
rect 393638 162893 393698 162963
rect 327257 162890 327323 162893
rect 327441 162890 327507 162893
rect 327257 162888 327507 162890
rect 327257 162832 327262 162888
rect 327318 162832 327446 162888
rect 327502 162832 327507 162888
rect 327257 162830 327507 162832
rect 327257 162827 327323 162830
rect 327441 162827 327507 162830
rect 329925 162890 329991 162893
rect 330109 162890 330175 162893
rect 329925 162888 330175 162890
rect 329925 162832 329930 162888
rect 329986 162832 330114 162888
rect 330170 162832 330175 162888
rect 329925 162830 330175 162832
rect 393638 162888 393747 162893
rect 393638 162832 393686 162888
rect 393742 162832 393747 162888
rect 393638 162830 393747 162832
rect 329925 162827 329991 162830
rect 330109 162827 330175 162830
rect 393681 162827 393747 162830
rect 245745 160034 245811 160037
rect 246113 160034 246179 160037
rect 245745 160032 246179 160034
rect 245745 159976 245750 160032
rect 245806 159976 246118 160032
rect 246174 159976 246179 160032
rect 245745 159974 246179 159976
rect 245745 159971 245811 159974
rect 246113 159971 246179 159974
rect 583520 158402 584960 158492
rect 583342 158342 584960 158402
rect 405406 157858 405412 157860
rect 398606 157798 405412 157858
rect 317321 157722 317387 157725
rect 378225 157722 378291 157725
rect 317321 157720 330586 157722
rect 317321 157664 317326 157720
rect 317382 157664 330586 157720
rect 317321 157662 330586 157664
rect 317321 157659 317387 157662
rect 249006 157524 249012 157588
rect 249076 157586 249082 157588
rect 306373 157586 306439 157589
rect 249076 157526 254042 157586
rect 249076 157524 249082 157526
rect 253982 157450 254042 157526
rect 275326 157584 306439 157586
rect 275326 157528 306378 157584
rect 306434 157528 306439 157584
rect 275326 157526 306439 157528
rect 330526 157586 330586 157662
rect 369902 157720 378291 157722
rect 369902 157664 378230 157720
rect 378286 157664 378291 157720
rect 369902 157662 378291 157664
rect 336733 157586 336799 157589
rect 360101 157586 360167 157589
rect 330526 157584 336799 157586
rect 330526 157528 336738 157584
rect 336794 157528 336799 157584
rect 330526 157526 336799 157528
rect 275326 157450 275386 157526
rect 306373 157523 306439 157526
rect 336733 157523 336799 157526
rect 350582 157584 360167 157586
rect 350582 157528 360106 157584
rect 360162 157528 360167 157584
rect 350582 157526 360167 157528
rect 253982 157390 275386 157450
rect 315941 157450 316007 157453
rect 317321 157450 317387 157453
rect 315941 157448 317387 157450
rect 315941 157392 315946 157448
rect 316002 157392 317326 157448
rect 317382 157392 317387 157448
rect 315941 157390 317387 157392
rect 315941 157387 316007 157390
rect 317321 157387 317387 157390
rect 346301 157450 346367 157453
rect 350582 157450 350642 157526
rect 360101 157523 360167 157526
rect 360285 157586 360351 157589
rect 360285 157584 369778 157586
rect 360285 157528 360290 157584
rect 360346 157528 369778 157584
rect 360285 157526 369778 157528
rect 360285 157523 360351 157526
rect 346301 157448 350642 157450
rect 346301 157392 346306 157448
rect 346362 157392 350642 157448
rect 346301 157390 350642 157392
rect 369718 157450 369778 157526
rect 369902 157450 369962 157662
rect 378225 157659 378291 157662
rect 386321 157722 386387 157725
rect 386321 157720 389098 157722
rect 386321 157664 386326 157720
rect 386382 157664 389098 157720
rect 386321 157662 389098 157664
rect 386321 157659 386387 157662
rect 369718 157390 369962 157450
rect 389038 157450 389098 157662
rect 398606 157586 398666 157798
rect 405406 157796 405412 157798
rect 405476 157796 405482 157860
rect 470550 157662 480178 157722
rect 417877 157586 417943 157589
rect 389222 157526 398666 157586
rect 408542 157584 417943 157586
rect 408542 157528 417882 157584
rect 417938 157528 417943 157584
rect 408542 157526 417943 157528
rect 389222 157450 389282 157526
rect 389038 157390 389282 157450
rect 346301 157387 346367 157390
rect 405590 157388 405596 157452
rect 405660 157450 405666 157452
rect 408542 157450 408602 157526
rect 417877 157523 417943 157526
rect 418153 157586 418219 157589
rect 437197 157586 437263 157589
rect 418153 157584 424978 157586
rect 418153 157528 418158 157584
rect 418214 157528 424978 157584
rect 418153 157526 424978 157528
rect 418153 157523 418219 157526
rect 405660 157390 408602 157450
rect 424918 157450 424978 157526
rect 427862 157584 437263 157586
rect 427862 157528 437202 157584
rect 437258 157528 437263 157584
rect 427862 157526 437263 157528
rect 427862 157450 427922 157526
rect 437197 157523 437263 157526
rect 437473 157586 437539 157589
rect 437473 157584 444298 157586
rect 437473 157528 437478 157584
rect 437534 157528 444298 157584
rect 437473 157526 444298 157528
rect 437473 157523 437539 157526
rect 424918 157390 427922 157450
rect 444238 157450 444298 157526
rect 447182 157526 463618 157586
rect 447182 157450 447242 157526
rect 444238 157390 447242 157450
rect 463558 157450 463618 157526
rect 470550 157450 470610 157662
rect 463558 157390 470610 157450
rect 480118 157450 480178 157662
rect 480302 157662 489930 157722
rect 480302 157450 480362 157662
rect 489870 157586 489930 157662
rect 499622 157662 509250 157722
rect 489870 157526 499498 157586
rect 480118 157390 480362 157450
rect 499438 157450 499498 157526
rect 499622 157450 499682 157662
rect 509190 157586 509250 157662
rect 518942 157662 528570 157722
rect 509190 157526 518818 157586
rect 499438 157390 499682 157450
rect 518758 157450 518818 157526
rect 518942 157450 519002 157662
rect 528510 157586 528570 157662
rect 538262 157662 547890 157722
rect 528510 157526 538138 157586
rect 518758 157390 519002 157450
rect 538078 157450 538138 157526
rect 538262 157450 538322 157662
rect 547830 157586 547890 157662
rect 557582 157662 567210 157722
rect 547830 157526 557458 157586
rect 538078 157390 538322 157450
rect 557398 157450 557458 157526
rect 557582 157450 557642 157662
rect 567150 157586 567210 157662
rect 583342 157586 583402 158342
rect 583520 158252 584960 158342
rect 567150 157526 576778 157586
rect 557398 157390 557642 157450
rect 576718 157450 576778 157526
rect 576902 157526 583402 157586
rect 576902 157450 576962 157526
rect 576718 157390 576962 157450
rect 405660 157388 405666 157390
rect 236269 154594 236335 154597
rect 236453 154594 236519 154597
rect 236269 154592 236519 154594
rect 236269 154536 236274 154592
rect 236330 154536 236458 154592
rect 236514 154536 236519 154592
rect 236269 154534 236519 154536
rect 236269 154531 236335 154534
rect 236453 154531 236519 154534
rect 340873 154594 340939 154597
rect 341333 154594 341399 154597
rect 340873 154592 341399 154594
rect 340873 154536 340878 154592
rect 340934 154536 341338 154592
rect 341394 154536 341399 154592
rect 340873 154534 341399 154536
rect 340873 154531 340939 154534
rect 341333 154531 341399 154534
rect 372521 154594 372587 154597
rect 372705 154594 372771 154597
rect 372521 154592 372771 154594
rect 372521 154536 372526 154592
rect 372582 154536 372710 154592
rect 372766 154536 372771 154592
rect 372521 154534 372771 154536
rect 372521 154531 372587 154534
rect 372705 154531 372771 154534
rect 310881 153370 310947 153373
rect 310838 153368 310947 153370
rect 310838 153312 310886 153368
rect 310942 153312 310947 153368
rect 310838 153307 310947 153312
rect 310838 153237 310898 153307
rect 230657 153234 230723 153237
rect 230841 153234 230907 153237
rect 230657 153232 230907 153234
rect 230657 153176 230662 153232
rect 230718 153176 230846 153232
rect 230902 153176 230907 153232
rect 230657 153174 230907 153176
rect 230657 153171 230723 153174
rect 230841 153171 230907 153174
rect 310789 153232 310898 153237
rect 310789 153176 310794 153232
rect 310850 153176 310898 153232
rect 310789 153174 310898 153176
rect 310789 153171 310855 153174
rect 331489 151874 331555 151877
rect 331673 151874 331739 151877
rect 331489 151872 331739 151874
rect 331489 151816 331494 151872
rect 331550 151816 331678 151872
rect 331734 151816 331739 151872
rect 331489 151814 331739 151816
rect 331489 151811 331555 151814
rect 331673 151811 331739 151814
rect -960 150786 480 150876
rect 3325 150786 3391 150789
rect -960 150784 3391 150786
rect -960 150728 3330 150784
rect 3386 150728 3391 150784
rect -960 150726 3391 150728
rect -960 150636 480 150726
rect 3325 150723 3391 150726
rect 583520 146556 584960 146796
rect 244365 144938 244431 144941
rect 244549 144938 244615 144941
rect 244365 144936 244615 144938
rect 244365 144880 244370 144936
rect 244426 144880 244554 144936
rect 244610 144880 244615 144936
rect 244365 144878 244615 144880
rect 244365 144875 244431 144878
rect 244549 144875 244615 144878
rect 325877 144938 325943 144941
rect 326061 144938 326127 144941
rect 325877 144936 326127 144938
rect 325877 144880 325882 144936
rect 325938 144880 326066 144936
rect 326122 144880 326127 144936
rect 325877 144878 326127 144880
rect 325877 144875 325943 144878
rect 326061 144875 326127 144878
rect 366725 144938 366791 144941
rect 367001 144938 367067 144941
rect 366725 144936 367067 144938
rect 366725 144880 366730 144936
rect 366786 144880 367006 144936
rect 367062 144880 367067 144936
rect 366725 144878 367067 144880
rect 366725 144875 366791 144878
rect 367001 144875 367067 144878
rect 245837 143578 245903 143581
rect 246021 143578 246087 143581
rect 245837 143576 246087 143578
rect 245837 143520 245842 143576
rect 245898 143520 246026 143576
rect 246082 143520 246087 143576
rect 245837 143518 246087 143520
rect 245837 143515 245903 143518
rect 246021 143515 246087 143518
rect 296621 140858 296687 140861
rect 296805 140858 296871 140861
rect 296621 140856 296871 140858
rect 296621 140800 296626 140856
rect 296682 140800 296810 140856
rect 296866 140800 296871 140856
rect 296621 140798 296871 140800
rect 296621 140795 296687 140798
rect 296805 140795 296871 140798
rect 245745 140722 245811 140725
rect 245929 140722 245995 140725
rect 245745 140720 245995 140722
rect 245745 140664 245750 140720
rect 245806 140664 245934 140720
rect 245990 140664 245995 140720
rect 245745 140662 245995 140664
rect 245745 140659 245811 140662
rect 245929 140659 245995 140662
rect -960 136370 480 136460
rect 2773 136370 2839 136373
rect -960 136368 2839 136370
rect -960 136312 2778 136368
rect 2834 136312 2839 136368
rect -960 136310 2839 136312
rect -960 136220 480 136310
rect 2773 136307 2839 136310
rect 337193 135418 337259 135421
rect 337193 135416 337394 135418
rect 337193 135360 337198 135416
rect 337254 135360 337394 135416
rect 337193 135358 337394 135360
rect 337193 135355 337259 135358
rect 236269 135282 236335 135285
rect 236453 135282 236519 135285
rect 236269 135280 236519 135282
rect 236269 135224 236274 135280
rect 236330 135224 236458 135280
rect 236514 135224 236519 135280
rect 236269 135222 236519 135224
rect 236269 135219 236335 135222
rect 236453 135219 236519 135222
rect 262673 135282 262739 135285
rect 262857 135282 262923 135285
rect 262673 135280 262923 135282
rect 262673 135224 262678 135280
rect 262734 135224 262862 135280
rect 262918 135224 262923 135280
rect 262673 135222 262923 135224
rect 262673 135219 262739 135222
rect 262857 135219 262923 135222
rect 323301 135282 323367 135285
rect 323485 135282 323551 135285
rect 323301 135280 323551 135282
rect 323301 135224 323306 135280
rect 323362 135224 323490 135280
rect 323546 135224 323551 135280
rect 323301 135222 323551 135224
rect 323301 135219 323367 135222
rect 323485 135219 323551 135222
rect 337193 135282 337259 135285
rect 337334 135282 337394 135358
rect 337193 135280 337394 135282
rect 337193 135224 337198 135280
rect 337254 135224 337394 135280
rect 337193 135222 337394 135224
rect 459921 135282 459987 135285
rect 460105 135282 460171 135285
rect 459921 135280 460171 135282
rect 459921 135224 459926 135280
rect 459982 135224 460110 135280
rect 460166 135224 460171 135280
rect 459921 135222 460171 135224
rect 337193 135219 337259 135222
rect 459921 135219 459987 135222
rect 460105 135219 460171 135222
rect 583520 134874 584960 134964
rect 583342 134814 584960 134874
rect 258022 134540 258028 134604
rect 258092 134602 258098 134604
rect 267641 134602 267707 134605
rect 258092 134600 267707 134602
rect 258092 134544 267646 134600
rect 267702 134544 267707 134600
rect 258092 134542 267707 134544
rect 258092 134540 258098 134542
rect 267641 134539 267707 134542
rect 267641 134330 267707 134333
rect 270309 134330 270375 134333
rect 267641 134328 270375 134330
rect 267641 134272 267646 134328
rect 267702 134272 270314 134328
rect 270370 134272 270375 134328
rect 267641 134270 270375 134272
rect 267641 134267 267707 134270
rect 270309 134267 270375 134270
rect 270493 134330 270559 134333
rect 487797 134330 487863 134333
rect 270493 134328 272626 134330
rect 270493 134272 270498 134328
rect 270554 134272 272626 134328
rect 270493 134270 272626 134272
rect 270493 134267 270559 134270
rect 245326 134132 245332 134196
rect 245396 134194 245402 134196
rect 258022 134194 258028 134196
rect 245396 134134 258028 134194
rect 245396 134132 245402 134134
rect 258022 134132 258028 134134
rect 258092 134132 258098 134196
rect 272566 134194 272626 134270
rect 396030 134270 405658 134330
rect 286961 134194 287027 134197
rect 272566 134192 287027 134194
rect 272566 134136 286966 134192
rect 287022 134136 287027 134192
rect 272566 134134 287027 134136
rect 286961 134131 287027 134134
rect 315941 134194 316007 134197
rect 328453 134194 328519 134197
rect 378225 134194 378291 134197
rect 315941 134192 323594 134194
rect 315941 134136 315946 134192
rect 316002 134136 323594 134192
rect 315941 134134 323594 134136
rect 315941 134131 316007 134134
rect 291837 134058 291903 134061
rect 309041 134058 309107 134061
rect 291837 134056 309107 134058
rect 291837 134000 291842 134056
rect 291898 134000 309046 134056
rect 309102 134000 309107 134056
rect 291837 133998 309107 134000
rect 291837 133995 291903 133998
rect 309041 133995 309107 133998
rect 247033 133922 247099 133925
rect 323534 133922 323594 134134
rect 328453 134192 340890 134194
rect 328453 134136 328458 134192
rect 328514 134136 340890 134192
rect 328453 134134 340890 134136
rect 328453 134131 328519 134134
rect 328453 133922 328519 133925
rect 247033 133920 247234 133922
rect 247033 133864 247038 133920
rect 247094 133864 247234 133920
rect 247033 133862 247234 133864
rect 323534 133920 328519 133922
rect 323534 133864 328458 133920
rect 328514 133864 328519 133920
rect 323534 133862 328519 133864
rect 340830 133922 340890 134134
rect 369902 134192 378291 134194
rect 369902 134136 378230 134192
rect 378286 134136 378291 134192
rect 369902 134134 378291 134136
rect 360101 134058 360167 134061
rect 350582 134056 360167 134058
rect 350582 134000 360106 134056
rect 360162 134000 360167 134056
rect 350582 133998 360167 134000
rect 350582 133922 350642 133998
rect 360101 133995 360167 133998
rect 360285 134058 360351 134061
rect 360285 134056 369778 134058
rect 360285 134000 360290 134056
rect 360346 134000 369778 134056
rect 360285 133998 369778 134000
rect 360285 133995 360351 133998
rect 340830 133862 350642 133922
rect 369718 133922 369778 133998
rect 369902 133922 369962 134134
rect 378225 134131 378291 134134
rect 386321 134194 386387 134197
rect 386321 134192 389098 134194
rect 386321 134136 386326 134192
rect 386382 134136 389098 134192
rect 386321 134134 389098 134136
rect 386321 134131 386387 134134
rect 369718 133862 369962 133922
rect 389038 133922 389098 134134
rect 396030 134058 396090 134270
rect 405598 134196 405658 134270
rect 483062 134328 487863 134330
rect 483062 134272 487802 134328
rect 487858 134272 487863 134328
rect 483062 134270 487863 134272
rect 405590 134132 405596 134196
rect 405660 134132 405666 134196
rect 456517 134194 456583 134197
rect 447182 134192 456583 134194
rect 447182 134136 456522 134192
rect 456578 134136 456583 134192
rect 447182 134134 456583 134136
rect 417877 134058 417943 134061
rect 389222 133998 396090 134058
rect 408542 134056 417943 134058
rect 408542 134000 417882 134056
rect 417938 134000 417943 134056
rect 408542 133998 417943 134000
rect 389222 133922 389282 133998
rect 389038 133862 389282 133922
rect 247033 133859 247099 133862
rect 247174 133786 247234 133862
rect 328453 133859 328519 133862
rect 405590 133860 405596 133924
rect 405660 133922 405666 133924
rect 408542 133922 408602 133998
rect 417877 133995 417943 133998
rect 418153 134058 418219 134061
rect 437197 134058 437263 134061
rect 418153 134056 424978 134058
rect 418153 134000 418158 134056
rect 418214 134000 424978 134056
rect 418153 133998 424978 134000
rect 418153 133995 418219 133998
rect 405660 133862 408602 133922
rect 424918 133922 424978 133998
rect 427862 134056 437263 134058
rect 427862 134000 437202 134056
rect 437258 134000 437263 134056
rect 427862 133998 437263 134000
rect 427862 133922 427922 133998
rect 437197 133995 437263 133998
rect 437565 134058 437631 134061
rect 437565 134056 444298 134058
rect 437565 134000 437570 134056
rect 437626 134000 444298 134056
rect 437565 133998 444298 134000
rect 437565 133995 437631 133998
rect 424918 133862 427922 133922
rect 444238 133922 444298 133998
rect 447182 133922 447242 134134
rect 456517 134131 456583 134134
rect 457437 134058 457503 134061
rect 475561 134058 475627 134061
rect 457437 134056 475627 134058
rect 457437 134000 457442 134056
rect 457498 134000 475566 134056
rect 475622 134000 475627 134056
rect 457437 133998 475627 134000
rect 457437 133995 457503 133998
rect 475561 133995 475627 133998
rect 482921 134058 482987 134061
rect 483062 134058 483122 134270
rect 487797 134267 487863 134270
rect 492622 134132 492628 134196
rect 492692 134194 492698 134196
rect 492692 134134 509250 134194
rect 492692 134132 492698 134134
rect 482921 134056 483122 134058
rect 482921 134000 482926 134056
rect 482982 134000 483122 134056
rect 482921 133998 483122 134000
rect 509190 134058 509250 134134
rect 518942 134134 528570 134194
rect 509190 133998 518818 134058
rect 482921 133995 482987 133998
rect 444238 133862 447242 133922
rect 487797 133922 487863 133925
rect 492622 133922 492628 133924
rect 487797 133920 492628 133922
rect 487797 133864 487802 133920
rect 487858 133864 492628 133920
rect 487797 133862 492628 133864
rect 405660 133860 405666 133862
rect 487797 133859 487863 133862
rect 492622 133860 492628 133862
rect 492692 133860 492698 133924
rect 518758 133922 518818 133998
rect 518942 133922 519002 134134
rect 528510 134058 528570 134134
rect 538262 134134 547890 134194
rect 528510 133998 538138 134058
rect 518758 133862 519002 133922
rect 538078 133922 538138 133998
rect 538262 133922 538322 134134
rect 547830 134058 547890 134134
rect 557582 134134 567210 134194
rect 547830 133998 557458 134058
rect 538078 133862 538322 133922
rect 557398 133922 557458 133998
rect 557582 133922 557642 134134
rect 567150 134058 567210 134134
rect 583342 134058 583402 134814
rect 583520 134724 584960 134814
rect 567150 133998 576778 134058
rect 557398 133862 557642 133922
rect 576718 133922 576778 133998
rect 576902 133998 583402 134058
rect 576902 133922 576962 133998
rect 576718 133862 576962 133922
rect 247309 133786 247375 133789
rect 247174 133784 247375 133786
rect 247174 133728 247314 133784
rect 247370 133728 247375 133784
rect 247174 133726 247375 133728
rect 247309 133723 247375 133726
rect 286961 133786 287027 133789
rect 291837 133786 291903 133789
rect 286961 133784 291903 133786
rect 286961 133728 286966 133784
rect 287022 133728 291842 133784
rect 291898 133728 291903 133784
rect 286961 133726 291903 133728
rect 286961 133723 287027 133726
rect 291837 133723 291903 133726
rect 265249 125762 265315 125765
rect 266721 125762 266787 125765
rect 267825 125762 267891 125765
rect 272241 125762 272307 125765
rect 273529 125762 273595 125765
rect 265206 125760 265315 125762
rect 265206 125704 265254 125760
rect 265310 125704 265315 125760
rect 265206 125699 265315 125704
rect 266678 125760 266787 125762
rect 266678 125704 266726 125760
rect 266782 125704 266787 125760
rect 266678 125699 266787 125704
rect 267782 125760 267891 125762
rect 267782 125704 267830 125760
rect 267886 125704 267891 125760
rect 267782 125699 267891 125704
rect 272198 125760 272307 125762
rect 272198 125704 272246 125760
rect 272302 125704 272307 125760
rect 272198 125699 272307 125704
rect 273486 125760 273595 125762
rect 273486 125704 273534 125760
rect 273590 125704 273595 125760
rect 273486 125699 273595 125704
rect 281717 125762 281783 125765
rect 284753 125762 284819 125765
rect 281717 125760 281826 125762
rect 281717 125704 281722 125760
rect 281778 125704 281826 125760
rect 281717 125699 281826 125704
rect 265206 125629 265266 125699
rect 266678 125629 266738 125699
rect 267782 125629 267842 125699
rect 272198 125629 272258 125699
rect 265206 125624 265315 125629
rect 265206 125568 265254 125624
rect 265310 125568 265315 125624
rect 265206 125566 265315 125568
rect 265249 125563 265315 125566
rect 266629 125624 266738 125629
rect 266629 125568 266634 125624
rect 266690 125568 266738 125624
rect 266629 125566 266738 125568
rect 267733 125624 267842 125629
rect 267733 125568 267738 125624
rect 267794 125568 267842 125624
rect 267733 125566 267842 125568
rect 272149 125624 272258 125629
rect 272149 125568 272154 125624
rect 272210 125568 272258 125624
rect 272149 125566 272258 125568
rect 273486 125629 273546 125699
rect 281766 125629 281826 125699
rect 284710 125760 284819 125762
rect 284710 125704 284758 125760
rect 284814 125704 284819 125760
rect 284710 125699 284819 125704
rect 284710 125629 284770 125699
rect 273486 125624 273595 125629
rect 273486 125568 273534 125624
rect 273590 125568 273595 125624
rect 273486 125566 273595 125568
rect 266629 125563 266695 125566
rect 267733 125563 267799 125566
rect 272149 125563 272215 125566
rect 273529 125563 273595 125566
rect 281717 125624 281826 125629
rect 281717 125568 281722 125624
rect 281778 125568 281826 125624
rect 281717 125566 281826 125568
rect 284661 125624 284770 125629
rect 284661 125568 284666 125624
rect 284722 125568 284770 125624
rect 284661 125566 284770 125568
rect 324589 125626 324655 125629
rect 324773 125626 324839 125629
rect 324589 125624 324839 125626
rect 324589 125568 324594 125624
rect 324650 125568 324778 125624
rect 324834 125568 324839 125624
rect 324589 125566 324839 125568
rect 281717 125563 281783 125566
rect 284661 125563 284727 125566
rect 324589 125563 324655 125566
rect 324773 125563 324839 125566
rect 325877 125626 325943 125629
rect 326061 125626 326127 125629
rect 325877 125624 326127 125626
rect 325877 125568 325882 125624
rect 325938 125568 326066 125624
rect 326122 125568 326127 125624
rect 325877 125566 326127 125568
rect 325877 125563 325943 125566
rect 326061 125563 326127 125566
rect 329925 125626 329991 125629
rect 330109 125626 330175 125629
rect 329925 125624 330175 125626
rect 329925 125568 329930 125624
rect 329986 125568 330114 125624
rect 330170 125568 330175 125624
rect 329925 125566 330175 125568
rect 329925 125563 329991 125566
rect 330109 125563 330175 125566
rect 375833 125626 375899 125629
rect 376109 125626 376175 125629
rect 375833 125624 376175 125626
rect 375833 125568 375838 125624
rect 375894 125568 376114 125624
rect 376170 125568 376175 125624
rect 375833 125566 376175 125568
rect 375833 125563 375899 125566
rect 376109 125563 376175 125566
rect 463877 125626 463943 125629
rect 464061 125626 464127 125629
rect 463877 125624 464127 125626
rect 463877 125568 463882 125624
rect 463938 125568 464066 125624
rect 464122 125568 464127 125624
rect 463877 125566 464127 125568
rect 463877 125563 463943 125566
rect 464061 125563 464127 125566
rect 285765 124266 285831 124269
rect 285949 124266 286015 124269
rect 285765 124264 286015 124266
rect 285765 124208 285770 124264
rect 285826 124208 285954 124264
rect 286010 124208 286015 124264
rect 285765 124206 286015 124208
rect 285765 124203 285831 124206
rect 285949 124203 286015 124206
rect 357617 124130 357683 124133
rect 357801 124130 357867 124133
rect 357617 124128 357867 124130
rect 357617 124072 357622 124128
rect 357678 124072 357806 124128
rect 357862 124072 357867 124128
rect 357617 124070 357867 124072
rect 357617 124067 357683 124070
rect 357801 124067 357867 124070
rect 315982 123524 315988 123588
rect 316052 123586 316058 123588
rect 325601 123586 325667 123589
rect 316052 123584 325667 123586
rect 316052 123528 325606 123584
rect 325662 123528 325667 123584
rect 316052 123526 325667 123528
rect 316052 123524 316058 123526
rect 325601 123523 325667 123526
rect 267774 123252 267780 123316
rect 267844 123314 267850 123316
rect 273713 123314 273779 123317
rect 267844 123312 273779 123314
rect 267844 123256 273718 123312
rect 273774 123256 273779 123312
rect 267844 123254 273779 123256
rect 267844 123252 267850 123254
rect 273713 123251 273779 123254
rect 273897 123314 273963 123317
rect 296529 123314 296595 123317
rect 273897 123312 296595 123314
rect 273897 123256 273902 123312
rect 273958 123256 296534 123312
rect 296590 123256 296595 123312
rect 273897 123254 296595 123256
rect 273897 123251 273963 123254
rect 296529 123251 296595 123254
rect 314561 123314 314627 123317
rect 315982 123314 315988 123316
rect 314561 123312 315988 123314
rect 314561 123256 314566 123312
rect 314622 123256 315988 123312
rect 314561 123254 315988 123256
rect 314561 123251 314627 123254
rect 315982 123252 315988 123254
rect 316052 123252 316058 123316
rect 487797 123314 487863 123317
rect 398606 123254 405658 123314
rect 248270 123116 248276 123180
rect 248340 123178 248346 123180
rect 328453 123178 328519 123181
rect 376661 123178 376727 123181
rect 248340 123118 254042 123178
rect 248340 123116 248346 123118
rect 253982 123042 254042 123118
rect 328453 123176 340890 123178
rect 328453 123120 328458 123176
rect 328514 123120 340890 123176
rect 328453 123118 340890 123120
rect 328453 123115 328519 123118
rect 267774 123042 267780 123044
rect 253982 122982 267780 123042
rect 267774 122980 267780 122982
rect 267844 122980 267850 123044
rect 296529 123042 296595 123045
rect 306005 123042 306071 123045
rect 296529 123040 306071 123042
rect 296529 122984 296534 123040
rect 296590 122984 306010 123040
rect 306066 122984 306071 123040
rect 296529 122982 306071 122984
rect 296529 122979 296595 122982
rect 306005 122979 306071 122982
rect 325601 123042 325667 123045
rect 328453 123042 328519 123045
rect 325601 123040 328519 123042
rect 325601 122984 325606 123040
rect 325662 122984 328458 123040
rect 328514 122984 328519 123040
rect 325601 122982 328519 122984
rect 325601 122979 325667 122982
rect 328453 122979 328519 122982
rect 340830 122906 340890 123118
rect 376661 123176 379530 123178
rect 376661 123120 376666 123176
rect 376722 123120 379530 123176
rect 376661 123118 379530 123120
rect 376661 123115 376727 123118
rect 365621 123042 365687 123045
rect 350582 123040 365687 123042
rect 350582 122984 365626 123040
rect 365682 122984 365687 123040
rect 350582 122982 365687 122984
rect 350582 122906 350642 122982
rect 365621 122979 365687 122982
rect 340830 122846 350642 122906
rect 365621 122906 365687 122909
rect 369669 122906 369735 122909
rect 365621 122904 369735 122906
rect 365621 122848 365626 122904
rect 365682 122848 369674 122904
rect 369730 122848 369735 122904
rect 365621 122846 369735 122848
rect 379470 122906 379530 123118
rect 398606 123042 398666 123254
rect 388486 122982 398666 123042
rect 388486 122906 388546 122982
rect 379470 122846 388546 122906
rect 405598 122906 405658 123254
rect 483062 123312 487863 123314
rect 483062 123256 487802 123312
rect 487858 123256 487863 123312
rect 483062 123254 487863 123256
rect 456517 123178 456583 123181
rect 447182 123176 456583 123178
rect 447182 123120 456522 123176
rect 456578 123120 456583 123176
rect 447182 123118 456583 123120
rect 417877 123042 417943 123045
rect 408542 123040 417943 123042
rect 408542 122984 417882 123040
rect 417938 122984 417943 123040
rect 408542 122982 417943 122984
rect 408542 122906 408602 122982
rect 417877 122979 417943 122982
rect 419349 123042 419415 123045
rect 437197 123042 437263 123045
rect 419349 123040 424978 123042
rect 419349 122984 419354 123040
rect 419410 122984 424978 123040
rect 419349 122982 424978 122984
rect 419349 122979 419415 122982
rect 405598 122846 408602 122906
rect 424918 122906 424978 122982
rect 427862 123040 437263 123042
rect 427862 122984 437202 123040
rect 437258 122984 437263 123040
rect 427862 122982 437263 122984
rect 427862 122906 427922 122982
rect 437197 122979 437263 122982
rect 437473 123042 437539 123045
rect 437473 123040 444298 123042
rect 437473 122984 437478 123040
rect 437534 122984 444298 123040
rect 437473 122982 444298 122984
rect 437473 122979 437539 122982
rect 424918 122846 427922 122906
rect 444238 122906 444298 122982
rect 447182 122906 447242 123118
rect 456517 123115 456583 123118
rect 471881 123178 471947 123181
rect 476021 123178 476087 123181
rect 471881 123176 476087 123178
rect 471881 123120 471886 123176
rect 471942 123120 476026 123176
rect 476082 123120 476087 123176
rect 471881 123118 476087 123120
rect 471881 123115 471947 123118
rect 476021 123115 476087 123118
rect 457437 123042 457503 123045
rect 462262 123042 462268 123044
rect 457437 123040 462268 123042
rect 457437 122984 457442 123040
rect 457498 122984 462268 123040
rect 457437 122982 462268 122984
rect 457437 122979 457503 122982
rect 462262 122980 462268 122982
rect 462332 122980 462338 123044
rect 476205 123042 476271 123045
rect 483062 123042 483122 123254
rect 487797 123251 487863 123254
rect 492622 123116 492628 123180
rect 492692 123178 492698 123180
rect 583520 123178 584960 123268
rect 492692 123118 509250 123178
rect 492692 123116 492698 123118
rect 476205 123040 483122 123042
rect 476205 122984 476210 123040
rect 476266 122984 483122 123040
rect 476205 122982 483122 122984
rect 509190 123042 509250 123118
rect 518942 123118 528570 123178
rect 509190 122982 518818 123042
rect 476205 122979 476271 122982
rect 444238 122846 447242 122906
rect 487797 122906 487863 122909
rect 492622 122906 492628 122908
rect 487797 122904 492628 122906
rect 487797 122848 487802 122904
rect 487858 122848 492628 122904
rect 487797 122846 492628 122848
rect 365621 122843 365687 122846
rect 369669 122843 369735 122846
rect 487797 122843 487863 122846
rect 492622 122844 492628 122846
rect 492692 122844 492698 122908
rect 518758 122906 518818 122982
rect 518942 122906 519002 123118
rect 528510 123042 528570 123118
rect 538262 123118 547890 123178
rect 528510 122982 538138 123042
rect 518758 122846 519002 122906
rect 538078 122906 538138 122982
rect 538262 122906 538322 123118
rect 547830 123042 547890 123118
rect 557582 123118 567210 123178
rect 547830 122982 557458 123042
rect 538078 122846 538322 122906
rect 557398 122906 557458 122982
rect 557582 122906 557642 123118
rect 567150 123042 567210 123118
rect 583342 123118 584960 123178
rect 583342 123042 583402 123118
rect 567150 122982 576778 123042
rect 557398 122846 557642 122906
rect 576718 122906 576778 122982
rect 576902 122982 583402 123042
rect 583520 123028 584960 123118
rect 576902 122906 576962 122982
rect 576718 122846 576962 122906
rect 259729 122770 259795 122773
rect 259913 122770 259979 122773
rect 259729 122768 259979 122770
rect 259729 122712 259734 122768
rect 259790 122712 259918 122768
rect 259974 122712 259979 122768
rect 259729 122710 259979 122712
rect 259729 122707 259795 122710
rect 259913 122707 259979 122710
rect 462262 122708 462268 122772
rect 462332 122770 462338 122772
rect 471881 122770 471947 122773
rect 462332 122768 471947 122770
rect 462332 122712 471886 122768
rect 471942 122712 471947 122768
rect 462332 122710 471947 122712
rect 462332 122708 462338 122710
rect 471881 122707 471947 122710
rect -960 122090 480 122180
rect 2773 122090 2839 122093
rect -960 122088 2839 122090
rect -960 122032 2778 122088
rect 2834 122032 2839 122088
rect -960 122030 2839 122032
rect -960 121940 480 122030
rect 2773 122027 2839 122030
rect 393589 121680 393655 121685
rect 393589 121624 393594 121680
rect 393650 121624 393655 121680
rect 393589 121619 393655 121624
rect 393592 121549 393652 121619
rect 393589 121544 393655 121549
rect 393589 121488 393594 121544
rect 393650 121488 393655 121544
rect 393589 121483 393655 121488
rect 250161 116106 250227 116109
rect 250118 116104 250227 116106
rect 250118 116048 250166 116104
rect 250222 116048 250227 116104
rect 250118 116043 250227 116048
rect 250118 115973 250178 116043
rect 236269 115970 236335 115973
rect 236453 115970 236519 115973
rect 236269 115968 236519 115970
rect 236269 115912 236274 115968
rect 236330 115912 236458 115968
rect 236514 115912 236519 115968
rect 236269 115910 236519 115912
rect 236269 115907 236335 115910
rect 236453 115907 236519 115910
rect 250069 115968 250178 115973
rect 250069 115912 250074 115968
rect 250130 115912 250178 115968
rect 250069 115910 250178 115912
rect 250069 115907 250135 115910
rect 327165 113386 327231 113389
rect 327165 113384 327274 113386
rect 327165 113328 327170 113384
rect 327226 113328 327274 113384
rect 327165 113323 327274 113328
rect 327214 113253 327274 113323
rect 327165 113248 327274 113253
rect 327165 113192 327170 113248
rect 327226 113192 327274 113248
rect 327165 113190 327274 113192
rect 327165 113187 327231 113190
rect 583520 111482 584960 111572
rect 583342 111422 584960 111482
rect 296662 111012 296668 111076
rect 296732 111074 296738 111076
rect 304942 111074 304948 111076
rect 296732 111014 304948 111074
rect 296732 111012 296738 111014
rect 304942 111012 304948 111014
rect 305012 111012 305018 111076
rect 315982 111012 315988 111076
rect 316052 111074 316058 111076
rect 325601 111074 325667 111077
rect 316052 111072 325667 111074
rect 316052 111016 325606 111072
rect 325662 111016 325667 111072
rect 316052 111014 325667 111016
rect 316052 111012 316058 111014
rect 325601 111011 325667 111014
rect 325734 110876 325740 110940
rect 325804 110876 325810 110940
rect 405406 110938 405412 110940
rect 336782 110878 341810 110938
rect 244038 110740 244044 110804
rect 244108 110802 244114 110804
rect 248413 110802 248479 110805
rect 244108 110800 248479 110802
rect 244108 110744 248418 110800
rect 248474 110744 248479 110800
rect 244108 110742 248479 110744
rect 244108 110740 244114 110742
rect 248413 110739 248479 110742
rect 296662 110740 296668 110804
rect 296732 110740 296738 110804
rect 304942 110740 304948 110804
rect 305012 110802 305018 110804
rect 306281 110802 306347 110805
rect 305012 110800 306347 110802
rect 305012 110744 306286 110800
rect 306342 110744 306347 110800
rect 305012 110742 306347 110744
rect 305012 110740 305018 110742
rect 254117 110666 254183 110669
rect 259361 110666 259427 110669
rect 254117 110664 259427 110666
rect 254117 110608 254122 110664
rect 254178 110608 259366 110664
rect 259422 110608 259427 110664
rect 254117 110606 259427 110608
rect 254117 110603 254183 110606
rect 259361 110603 259427 110606
rect 285622 110604 285628 110668
rect 285692 110666 285698 110668
rect 296670 110666 296730 110740
rect 306281 110739 306347 110742
rect 315941 110804 316007 110805
rect 315941 110800 315988 110804
rect 316052 110802 316058 110804
rect 325601 110802 325667 110805
rect 325742 110802 325802 110876
rect 315941 110744 315946 110800
rect 315941 110740 315988 110744
rect 316052 110742 316134 110802
rect 325601 110800 325802 110802
rect 325601 110744 325606 110800
rect 325662 110744 325802 110800
rect 325601 110742 325802 110744
rect 335169 110802 335235 110805
rect 336782 110802 336842 110878
rect 335169 110800 336842 110802
rect 335169 110744 335174 110800
rect 335230 110744 336842 110800
rect 335169 110742 336842 110744
rect 316052 110740 316058 110742
rect 315941 110739 316007 110740
rect 325601 110739 325667 110742
rect 335169 110739 335235 110742
rect 285692 110606 296730 110666
rect 285692 110604 285698 110606
rect 325734 110604 325740 110668
rect 325804 110666 325810 110668
rect 335169 110666 335235 110669
rect 325804 110664 335235 110666
rect 325804 110608 335174 110664
rect 335230 110608 335235 110664
rect 325804 110606 335235 110608
rect 325804 110604 325810 110606
rect 335169 110603 335235 110606
rect 267641 110530 267707 110533
rect 277342 110530 277348 110532
rect 267641 110528 277348 110530
rect 267641 110472 267646 110528
rect 267702 110472 277348 110528
rect 267641 110470 277348 110472
rect 267641 110467 267707 110470
rect 277342 110468 277348 110470
rect 277412 110468 277418 110532
rect 341750 110530 341810 110878
rect 398606 110878 405412 110938
rect 369718 110742 379530 110802
rect 357382 110666 357388 110668
rect 350582 110606 357388 110666
rect 350582 110530 350642 110606
rect 357382 110604 357388 110606
rect 357452 110604 357458 110668
rect 341750 110470 350642 110530
rect 357566 110468 357572 110532
rect 357636 110530 357642 110532
rect 369718 110530 369778 110742
rect 357636 110470 369778 110530
rect 379470 110530 379530 110742
rect 398606 110666 398666 110878
rect 405406 110876 405412 110878
rect 405476 110876 405482 110940
rect 487797 110938 487863 110941
rect 483062 110936 487863 110938
rect 483062 110880 487802 110936
rect 487858 110880 487863 110936
rect 483062 110878 487863 110880
rect 456517 110802 456583 110805
rect 447182 110800 456583 110802
rect 447182 110744 456522 110800
rect 456578 110744 456583 110800
rect 447182 110742 456583 110744
rect 417877 110666 417943 110669
rect 389222 110606 398666 110666
rect 408542 110664 417943 110666
rect 408542 110608 417882 110664
rect 417938 110608 417943 110664
rect 408542 110606 417943 110608
rect 389222 110530 389282 110606
rect 379470 110470 389282 110530
rect 357636 110468 357642 110470
rect 405590 110468 405596 110532
rect 405660 110530 405666 110532
rect 408542 110530 408602 110606
rect 417877 110603 417943 110606
rect 418153 110666 418219 110669
rect 437197 110666 437263 110669
rect 418153 110664 424978 110666
rect 418153 110608 418158 110664
rect 418214 110608 424978 110664
rect 418153 110606 424978 110608
rect 418153 110603 418219 110606
rect 405660 110470 408602 110530
rect 424918 110530 424978 110606
rect 427862 110664 437263 110666
rect 427862 110608 437202 110664
rect 437258 110608 437263 110664
rect 427862 110606 437263 110608
rect 427862 110530 427922 110606
rect 437197 110603 437263 110606
rect 437473 110666 437539 110669
rect 437473 110664 444298 110666
rect 437473 110608 437478 110664
rect 437534 110608 444298 110664
rect 437473 110606 444298 110608
rect 437473 110603 437539 110606
rect 424918 110470 427922 110530
rect 444238 110530 444298 110606
rect 447182 110530 447242 110742
rect 456517 110739 456583 110742
rect 471881 110802 471947 110805
rect 476021 110802 476087 110805
rect 471881 110800 476087 110802
rect 471881 110744 471886 110800
rect 471942 110744 476026 110800
rect 476082 110744 476087 110800
rect 471881 110742 476087 110744
rect 471881 110739 471947 110742
rect 476021 110739 476087 110742
rect 457437 110666 457503 110669
rect 462262 110666 462268 110668
rect 457437 110664 462268 110666
rect 457437 110608 457442 110664
rect 457498 110608 462268 110664
rect 457437 110606 462268 110608
rect 457437 110603 457503 110606
rect 462262 110604 462268 110606
rect 462332 110604 462338 110668
rect 476205 110666 476271 110669
rect 483062 110666 483122 110878
rect 487797 110875 487863 110878
rect 492622 110740 492628 110804
rect 492692 110802 492698 110804
rect 492692 110742 509250 110802
rect 492692 110740 492698 110742
rect 476205 110664 483122 110666
rect 476205 110608 476210 110664
rect 476266 110608 483122 110664
rect 476205 110606 483122 110608
rect 509190 110666 509250 110742
rect 518942 110742 528570 110802
rect 509190 110606 518818 110666
rect 476205 110603 476271 110606
rect 444238 110470 447242 110530
rect 487797 110530 487863 110533
rect 492622 110530 492628 110532
rect 487797 110528 492628 110530
rect 487797 110472 487802 110528
rect 487858 110472 492628 110528
rect 487797 110470 492628 110472
rect 405660 110468 405666 110470
rect 487797 110467 487863 110470
rect 492622 110468 492628 110470
rect 492692 110468 492698 110532
rect 518758 110530 518818 110606
rect 518942 110530 519002 110742
rect 528510 110666 528570 110742
rect 538262 110742 547890 110802
rect 528510 110606 538138 110666
rect 518758 110470 519002 110530
rect 538078 110530 538138 110606
rect 538262 110530 538322 110742
rect 547830 110666 547890 110742
rect 557582 110742 567210 110802
rect 547830 110606 557458 110666
rect 538078 110470 538322 110530
rect 557398 110530 557458 110606
rect 557582 110530 557642 110742
rect 567150 110666 567210 110742
rect 583342 110666 583402 111422
rect 583520 111332 584960 111422
rect 567150 110606 576778 110666
rect 557398 110470 557642 110530
rect 576718 110530 576778 110606
rect 576902 110606 583402 110666
rect 576902 110530 576962 110606
rect 576718 110470 576962 110530
rect 462262 110332 462268 110396
rect 462332 110394 462338 110396
rect 471881 110394 471947 110397
rect 462332 110392 471947 110394
rect 462332 110336 471886 110392
rect 471942 110336 471947 110392
rect 462332 110334 471947 110336
rect 462332 110332 462338 110334
rect 471881 110331 471947 110334
rect 277342 110196 277348 110260
rect 277412 110258 277418 110260
rect 285622 110258 285628 110260
rect 277412 110198 285628 110258
rect 277412 110196 277418 110198
rect 285622 110196 285628 110198
rect 285692 110196 285698 110260
rect -960 107674 480 107764
rect 3509 107674 3575 107677
rect -960 107672 3575 107674
rect -960 107616 3514 107672
rect 3570 107616 3575 107672
rect -960 107614 3575 107616
rect -960 107524 480 107614
rect 3509 107611 3575 107614
rect 366725 106314 366791 106317
rect 367001 106314 367067 106317
rect 366725 106312 367067 106314
rect 366725 106256 366730 106312
rect 366786 106256 367006 106312
rect 367062 106256 367067 106312
rect 366725 106254 367067 106256
rect 366725 106251 366791 106254
rect 367001 106251 367067 106254
rect 583520 99636 584960 99876
rect 236269 96658 236335 96661
rect 236453 96658 236519 96661
rect 236269 96656 236519 96658
rect 236269 96600 236274 96656
rect 236330 96600 236458 96656
rect 236514 96600 236519 96656
rect 236269 96598 236519 96600
rect 236269 96595 236335 96598
rect 236453 96595 236519 96598
rect 459921 96658 459987 96661
rect 460105 96658 460171 96661
rect 459921 96656 460171 96658
rect 459921 96600 459926 96656
rect 459982 96600 460110 96656
rect 460166 96600 460171 96656
rect 459921 96598 460171 96600
rect 459921 96595 459987 96598
rect 460105 96595 460171 96598
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 299422 87348 299428 87412
rect 299492 87410 299498 87412
rect 331857 87410 331923 87413
rect 299492 87350 302066 87410
rect 299492 87348 299498 87350
rect 239990 87212 239996 87276
rect 240060 87274 240066 87276
rect 286225 87274 286291 87277
rect 240060 87214 249810 87274
rect 240060 87212 240066 87214
rect 249750 87138 249810 87214
rect 273854 87272 286291 87274
rect 273854 87216 286230 87272
rect 286286 87216 286291 87272
rect 273854 87214 286291 87216
rect 273069 87138 273135 87141
rect 249750 87136 273135 87138
rect 249750 87080 273074 87136
rect 273130 87080 273135 87136
rect 249750 87078 273135 87080
rect 273069 87075 273135 87078
rect 273253 87138 273319 87141
rect 273854 87138 273914 87214
rect 286225 87211 286291 87214
rect 299422 87138 299428 87140
rect 273253 87136 273914 87138
rect 273253 87080 273258 87136
rect 273314 87080 273914 87136
rect 273253 87078 273914 87080
rect 289494 87078 299428 87138
rect 273253 87075 273319 87078
rect 286225 87002 286291 87005
rect 289494 87002 289554 87078
rect 299422 87076 299428 87078
rect 299492 87076 299498 87140
rect 302006 87138 302066 87350
rect 322246 87408 331923 87410
rect 322246 87352 331862 87408
rect 331918 87352 331923 87408
rect 322246 87350 331923 87352
rect 322246 87138 322306 87350
rect 331857 87347 331923 87350
rect 481582 87348 481588 87412
rect 481652 87410 481658 87412
rect 491201 87410 491267 87413
rect 481652 87408 491267 87410
rect 481652 87352 491206 87408
rect 491262 87352 491267 87408
rect 481652 87350 491267 87352
rect 481652 87348 481658 87350
rect 491201 87347 491267 87350
rect 367001 87274 367067 87277
rect 454033 87274 454099 87277
rect 366958 87272 367067 87274
rect 366958 87216 367006 87272
rect 367062 87216 367067 87272
rect 366958 87211 367067 87216
rect 447182 87272 454099 87274
rect 447182 87216 454038 87272
rect 454094 87216 454099 87272
rect 447182 87214 454099 87216
rect 366958 87141 367018 87211
rect 302006 87078 311818 87138
rect 286225 87000 289554 87002
rect 286225 86944 286230 87000
rect 286286 86944 289554 87000
rect 286225 86942 289554 86944
rect 311758 87002 311818 87078
rect 311942 87078 322306 87138
rect 331857 87138 331923 87141
rect 336733 87138 336799 87141
rect 331857 87136 336799 87138
rect 331857 87080 331862 87136
rect 331918 87080 336738 87136
rect 336794 87080 336799 87136
rect 331857 87078 336799 87080
rect 311942 87002 312002 87078
rect 331857 87075 331923 87078
rect 336733 87075 336799 87078
rect 350582 87078 360210 87138
rect 366958 87136 367067 87141
rect 379053 87138 379119 87141
rect 396073 87138 396139 87141
rect 417877 87138 417943 87141
rect 366958 87080 367006 87136
rect 367062 87080 367067 87136
rect 366958 87078 367067 87080
rect 311758 86942 312002 87002
rect 346301 87002 346367 87005
rect 350582 87002 350642 87078
rect 346301 87000 350642 87002
rect 346301 86944 346306 87000
rect 346362 86944 350642 87000
rect 346301 86942 350642 86944
rect 360150 87002 360210 87078
rect 367001 87075 367067 87078
rect 369902 87136 379119 87138
rect 369902 87080 379058 87136
rect 379114 87080 379119 87136
rect 369902 87078 379119 87080
rect 369902 87002 369962 87078
rect 379053 87075 379119 87078
rect 389222 87136 396139 87138
rect 389222 87080 396078 87136
rect 396134 87080 396139 87136
rect 389222 87078 396139 87080
rect 360150 86942 369962 87002
rect 386321 87002 386387 87005
rect 389222 87002 389282 87078
rect 396073 87075 396139 87078
rect 408542 87136 417943 87138
rect 408542 87080 417882 87136
rect 417938 87080 417943 87136
rect 408542 87078 417943 87080
rect 386321 87000 389282 87002
rect 386321 86944 386326 87000
rect 386382 86944 389282 87000
rect 386321 86942 389282 86944
rect 405549 87002 405615 87005
rect 408542 87002 408602 87078
rect 417877 87075 417943 87078
rect 418613 87138 418679 87141
rect 437197 87138 437263 87141
rect 418613 87136 424978 87138
rect 418613 87080 418618 87136
rect 418674 87080 424978 87136
rect 418613 87078 424978 87080
rect 418613 87075 418679 87078
rect 405549 87000 408602 87002
rect 405549 86944 405554 87000
rect 405610 86944 408602 87000
rect 405549 86942 408602 86944
rect 424918 87002 424978 87078
rect 427862 87136 437263 87138
rect 427862 87080 437202 87136
rect 437258 87080 437263 87136
rect 427862 87078 437263 87080
rect 427862 87002 427922 87078
rect 437197 87075 437263 87078
rect 437473 87138 437539 87141
rect 437473 87136 444298 87138
rect 437473 87080 437478 87136
rect 437534 87080 444298 87136
rect 437473 87078 444298 87080
rect 437473 87075 437539 87078
rect 424918 86942 427922 87002
rect 444238 87002 444298 87078
rect 447182 87002 447242 87214
rect 454033 87211 454099 87214
rect 467925 87274 467991 87277
rect 476021 87274 476087 87277
rect 467925 87272 476087 87274
rect 467925 87216 467930 87272
rect 467986 87216 476026 87272
rect 476082 87216 476087 87272
rect 467925 87214 476087 87216
rect 467925 87211 467991 87214
rect 476021 87211 476087 87214
rect 502241 87274 502307 87277
rect 502241 87272 509250 87274
rect 502241 87216 502246 87272
rect 502302 87216 509250 87272
rect 502241 87214 509250 87216
rect 502241 87211 502307 87214
rect 463417 87172 463483 87175
rect 463417 87170 463618 87172
rect 463417 87114 463422 87170
rect 463478 87138 463618 87170
rect 463693 87138 463759 87141
rect 463478 87136 463759 87138
rect 463478 87114 463698 87136
rect 463417 87112 463698 87114
rect 463417 87109 463483 87112
rect 463558 87080 463698 87112
rect 463754 87080 463759 87136
rect 463558 87078 463759 87080
rect 463693 87075 463759 87078
rect 476205 87138 476271 87141
rect 481582 87138 481588 87140
rect 476205 87136 481588 87138
rect 476205 87080 476210 87136
rect 476266 87080 481588 87136
rect 476205 87078 481588 87080
rect 476205 87075 476271 87078
rect 481582 87076 481588 87078
rect 481652 87076 481658 87140
rect 509190 87138 509250 87214
rect 518942 87214 528570 87274
rect 509190 87078 518818 87138
rect 444238 86942 447242 87002
rect 491201 87002 491267 87005
rect 494605 87002 494671 87005
rect 491201 87000 494671 87002
rect 491201 86944 491206 87000
rect 491262 86944 494610 87000
rect 494666 86944 494671 87000
rect 491201 86942 494671 86944
rect 518758 87002 518818 87078
rect 518942 87002 519002 87214
rect 528510 87138 528570 87214
rect 538262 87214 547890 87274
rect 528510 87078 538138 87138
rect 518758 86942 519002 87002
rect 538078 87002 538138 87078
rect 538262 87002 538322 87214
rect 547830 87138 547890 87214
rect 557582 87214 567210 87274
rect 547830 87078 557458 87138
rect 538078 86942 538322 87002
rect 557398 87002 557458 87078
rect 557582 87002 557642 87214
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 557398 86942 557642 87002
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 286225 86939 286291 86942
rect 346301 86939 346367 86942
rect 386321 86939 386387 86942
rect 405549 86939 405615 86942
rect 491201 86939 491267 86942
rect 494605 86939 494671 86942
rect -960 78978 480 79068
rect 2773 78978 2839 78981
rect -960 78976 2839 78978
rect -960 78920 2778 78976
rect 2834 78920 2839 78976
rect -960 78918 2839 78920
rect -960 78828 480 78918
rect 2773 78915 2839 78918
rect 251449 77346 251515 77349
rect 251633 77346 251699 77349
rect 251449 77344 251699 77346
rect 251449 77288 251454 77344
rect 251510 77288 251638 77344
rect 251694 77288 251699 77344
rect 251449 77286 251699 77288
rect 251449 77283 251515 77286
rect 251633 77283 251699 77286
rect 473302 76468 473308 76532
rect 473372 76530 473378 76532
rect 482921 76530 482987 76533
rect 473372 76528 482987 76530
rect 473372 76472 482926 76528
rect 482982 76472 482987 76528
rect 473372 76470 482987 76472
rect 473372 76468 473378 76470
rect 482921 76467 482987 76470
rect 487797 76394 487863 76397
rect 398606 76334 405658 76394
rect 299422 76196 299428 76260
rect 299492 76258 299498 76260
rect 307702 76258 307708 76260
rect 299492 76198 307708 76258
rect 299492 76196 299498 76198
rect 307702 76196 307708 76198
rect 307772 76196 307778 76260
rect 378225 76258 378291 76261
rect 331078 76198 340890 76258
rect 241278 76060 241284 76124
rect 241348 76122 241354 76124
rect 251173 76122 251239 76125
rect 241348 76120 251239 76122
rect 241348 76064 251178 76120
rect 251234 76064 251239 76120
rect 241348 76062 251239 76064
rect 241348 76060 241354 76062
rect 251173 76059 251239 76062
rect 275369 76122 275435 76125
rect 284661 76122 284727 76125
rect 275369 76120 284727 76122
rect 275369 76064 275374 76120
rect 275430 76064 284666 76120
rect 284722 76064 284727 76120
rect 275369 76062 284727 76064
rect 275369 76059 275435 76062
rect 284661 76059 284727 76062
rect 260782 75924 260788 75988
rect 260852 75986 260858 75988
rect 270493 75986 270559 75989
rect 260852 75984 270559 75986
rect 260852 75928 270498 75984
rect 270554 75928 270559 75984
rect 260852 75926 270559 75928
rect 260852 75924 260858 75926
rect 270493 75923 270559 75926
rect 284753 75986 284819 75989
rect 299422 75986 299428 75988
rect 284753 75984 284954 75986
rect 284753 75928 284758 75984
rect 284814 75928 284954 75984
rect 284753 75926 284954 75928
rect 284753 75923 284819 75926
rect 251173 75714 251239 75717
rect 260782 75714 260788 75716
rect 251173 75712 260788 75714
rect 251173 75656 251178 75712
rect 251234 75656 260788 75712
rect 251173 75654 260788 75656
rect 251173 75651 251239 75654
rect 260782 75652 260788 75654
rect 260852 75652 260858 75716
rect 284894 75714 284954 75926
rect 288206 75926 299428 75986
rect 288206 75714 288266 75926
rect 299422 75924 299428 75926
rect 299492 75924 299498 75988
rect 307702 75924 307708 75988
rect 307772 75986 307778 75988
rect 331078 75986 331138 76198
rect 307772 75926 331138 75986
rect 340830 75986 340890 76198
rect 369902 76256 378291 76258
rect 369902 76200 378230 76256
rect 378286 76200 378291 76256
rect 369902 76198 378291 76200
rect 360101 76122 360167 76125
rect 350582 76120 360167 76122
rect 350582 76064 360106 76120
rect 360162 76064 360167 76120
rect 350582 76062 360167 76064
rect 350582 75986 350642 76062
rect 360101 76059 360167 76062
rect 360285 76122 360351 76125
rect 360285 76120 369778 76122
rect 360285 76064 360290 76120
rect 360346 76064 369778 76120
rect 360285 76062 369778 76064
rect 360285 76059 360351 76062
rect 340830 75926 350642 75986
rect 369718 75986 369778 76062
rect 369902 75986 369962 76198
rect 378225 76195 378291 76198
rect 386321 76258 386387 76261
rect 386321 76256 389098 76258
rect 386321 76200 386326 76256
rect 386382 76200 389098 76256
rect 386321 76198 389098 76200
rect 386321 76195 386387 76198
rect 369718 75926 369962 75986
rect 389038 75986 389098 76198
rect 398606 76122 398666 76334
rect 389222 76062 398666 76122
rect 389222 75986 389282 76062
rect 389038 75926 389282 75986
rect 405598 75986 405658 76334
rect 483062 76392 487863 76394
rect 483062 76336 487802 76392
rect 487858 76336 487863 76392
rect 483062 76334 487863 76336
rect 467925 76258 467991 76261
rect 473302 76258 473308 76260
rect 447182 76198 456626 76258
rect 417877 76122 417943 76125
rect 408542 76120 417943 76122
rect 408542 76064 417882 76120
rect 417938 76064 417943 76120
rect 408542 76062 417943 76064
rect 408542 75986 408602 76062
rect 417877 76059 417943 76062
rect 419349 76122 419415 76125
rect 434713 76122 434779 76125
rect 419349 76120 424978 76122
rect 419349 76064 419354 76120
rect 419410 76064 424978 76120
rect 419349 76062 424978 76064
rect 419349 76059 419415 76062
rect 405598 75926 408602 75986
rect 424918 75986 424978 76062
rect 427862 76120 434779 76122
rect 427862 76064 434718 76120
rect 434774 76064 434779 76120
rect 427862 76062 434779 76064
rect 427862 75986 427922 76062
rect 434713 76059 434779 76062
rect 437473 76122 437539 76125
rect 437473 76120 444298 76122
rect 437473 76064 437478 76120
rect 437534 76064 444298 76120
rect 437473 76062 444298 76064
rect 437473 76059 437539 76062
rect 424918 75926 427922 75986
rect 444238 75986 444298 76062
rect 447182 75986 447242 76198
rect 456566 76122 456626 76198
rect 467925 76256 473308 76258
rect 467925 76200 467930 76256
rect 467986 76200 473308 76256
rect 467925 76198 473308 76200
rect 467925 76195 467991 76198
rect 473302 76196 473308 76198
rect 473372 76196 473378 76260
rect 463693 76122 463759 76125
rect 456566 76120 463759 76122
rect 456566 76064 463698 76120
rect 463754 76064 463759 76120
rect 456566 76062 463759 76064
rect 463693 76059 463759 76062
rect 482921 76122 482987 76125
rect 483062 76122 483122 76334
rect 487797 76331 487863 76334
rect 492622 76196 492628 76260
rect 492692 76258 492698 76260
rect 583520 76258 584960 76348
rect 492692 76198 509250 76258
rect 492692 76196 492698 76198
rect 482921 76120 483122 76122
rect 482921 76064 482926 76120
rect 482982 76064 483122 76120
rect 482921 76062 483122 76064
rect 509190 76122 509250 76198
rect 518942 76198 528570 76258
rect 509190 76062 518818 76122
rect 482921 76059 482987 76062
rect 444238 75926 447242 75986
rect 487797 75986 487863 75989
rect 492622 75986 492628 75988
rect 487797 75984 492628 75986
rect 487797 75928 487802 75984
rect 487858 75928 492628 75984
rect 487797 75926 492628 75928
rect 307772 75924 307778 75926
rect 487797 75923 487863 75926
rect 492622 75924 492628 75926
rect 492692 75924 492698 75988
rect 518758 75986 518818 76062
rect 518942 75986 519002 76198
rect 528510 76122 528570 76198
rect 538262 76198 547890 76258
rect 528510 76062 538138 76122
rect 518758 75926 519002 75986
rect 538078 75986 538138 76062
rect 538262 75986 538322 76198
rect 547830 76122 547890 76198
rect 557582 76198 567210 76258
rect 547830 76062 557458 76122
rect 538078 75926 538322 75986
rect 557398 75986 557458 76062
rect 557582 75986 557642 76198
rect 567150 76122 567210 76198
rect 583342 76198 584960 76258
rect 583342 76122 583402 76198
rect 567150 76062 576778 76122
rect 557398 75926 557642 75986
rect 576718 75986 576778 76062
rect 576902 76062 583402 76122
rect 583520 76108 584960 76198
rect 576902 75986 576962 76062
rect 576718 75926 576962 75986
rect 310421 75850 310487 75853
rect 310789 75850 310855 75853
rect 310421 75848 310855 75850
rect 310421 75792 310426 75848
rect 310482 75792 310794 75848
rect 310850 75792 310855 75848
rect 310421 75790 310855 75792
rect 310421 75787 310487 75790
rect 310789 75787 310855 75790
rect 284894 75654 288266 75714
rect 244549 66466 244615 66469
rect 244230 66464 244615 66466
rect 244230 66408 244554 66464
rect 244610 66408 244615 66464
rect 244230 66406 244615 66408
rect 244230 66330 244290 66406
rect 244549 66403 244615 66406
rect 244365 66330 244431 66333
rect 244230 66328 244431 66330
rect 244230 66272 244370 66328
rect 244426 66272 244431 66328
rect 244230 66270 244431 66272
rect 244365 66267 244431 66270
rect 310421 66330 310487 66333
rect 310789 66330 310855 66333
rect 310421 66328 310855 66330
rect 310421 66272 310426 66328
rect 310482 66272 310794 66328
rect 310850 66272 310855 66328
rect 310421 66270 310855 66272
rect 310421 66267 310487 66270
rect 310789 66267 310855 66270
rect 262673 66194 262739 66197
rect 262949 66194 263015 66197
rect 331397 66194 331463 66197
rect 262673 66192 263015 66194
rect 262673 66136 262678 66192
rect 262734 66136 262954 66192
rect 263010 66136 263015 66192
rect 262673 66134 263015 66136
rect 262673 66131 262739 66134
rect 262949 66131 263015 66134
rect 331262 66192 331463 66194
rect 331262 66136 331402 66192
rect 331458 66136 331463 66192
rect 331262 66134 331463 66136
rect 331262 66058 331322 66134
rect 331397 66131 331463 66134
rect 331581 66058 331647 66061
rect 331262 66056 331647 66058
rect 331262 66000 331586 66056
rect 331642 66000 331647 66056
rect 331262 65998 331647 66000
rect 331581 65995 331647 65998
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect 583520 64562 584960 64652
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 583342 64502 584960 64562
rect 317270 64018 317276 64020
rect 307710 63958 317276 64018
rect 280102 63882 280108 63884
rect 275326 63822 280108 63882
rect 237230 63684 237236 63748
rect 237300 63746 237306 63748
rect 237300 63686 256066 63746
rect 237300 63684 237306 63686
rect 256006 63610 256066 63686
rect 275326 63610 275386 63822
rect 280102 63820 280108 63822
rect 280172 63820 280178 63884
rect 288566 63684 288572 63748
rect 288636 63746 288642 63748
rect 307710 63746 307770 63958
rect 317270 63956 317276 63958
rect 317340 63956 317346 64020
rect 405406 64018 405412 64020
rect 398606 63958 405412 64018
rect 327022 63820 327028 63884
rect 327092 63882 327098 63884
rect 378225 63882 378291 63885
rect 327092 63822 340890 63882
rect 327092 63820 327098 63822
rect 288636 63686 307770 63746
rect 288636 63684 288642 63686
rect 256006 63550 275386 63610
rect 280102 63548 280108 63612
rect 280172 63610 280178 63612
rect 288382 63610 288388 63612
rect 280172 63550 288388 63610
rect 280172 63548 280178 63550
rect 288382 63548 288388 63550
rect 288452 63548 288458 63612
rect 317270 63548 317276 63612
rect 317340 63610 317346 63612
rect 327022 63610 327028 63612
rect 317340 63550 327028 63610
rect 317340 63548 317346 63550
rect 327022 63548 327028 63550
rect 327092 63548 327098 63612
rect 340830 63610 340890 63822
rect 369902 63880 378291 63882
rect 369902 63824 378230 63880
rect 378286 63824 378291 63880
rect 369902 63822 378291 63824
rect 360101 63746 360167 63749
rect 350582 63744 360167 63746
rect 350582 63688 360106 63744
rect 360162 63688 360167 63744
rect 350582 63686 360167 63688
rect 350582 63610 350642 63686
rect 360101 63683 360167 63686
rect 360285 63746 360351 63749
rect 360285 63744 369778 63746
rect 360285 63688 360290 63744
rect 360346 63688 369778 63744
rect 360285 63686 369778 63688
rect 360285 63683 360351 63686
rect 340830 63550 350642 63610
rect 369718 63610 369778 63686
rect 369902 63610 369962 63822
rect 378225 63819 378291 63822
rect 386321 63882 386387 63885
rect 386321 63880 389098 63882
rect 386321 63824 386326 63880
rect 386382 63824 389098 63880
rect 386321 63822 389098 63824
rect 386321 63819 386387 63822
rect 369718 63550 369962 63610
rect 389038 63610 389098 63822
rect 398606 63746 398666 63958
rect 405406 63956 405412 63958
rect 405476 63956 405482 64020
rect 470550 63822 480178 63882
rect 417877 63746 417943 63749
rect 389222 63686 398666 63746
rect 408542 63744 417943 63746
rect 408542 63688 417882 63744
rect 417938 63688 417943 63744
rect 408542 63686 417943 63688
rect 389222 63610 389282 63686
rect 389038 63550 389282 63610
rect 405590 63548 405596 63612
rect 405660 63610 405666 63612
rect 408542 63610 408602 63686
rect 417877 63683 417943 63686
rect 418153 63746 418219 63749
rect 437197 63746 437263 63749
rect 418153 63744 424978 63746
rect 418153 63688 418158 63744
rect 418214 63688 424978 63744
rect 418153 63686 424978 63688
rect 418153 63683 418219 63686
rect 405660 63550 408602 63610
rect 424918 63610 424978 63686
rect 427862 63744 437263 63746
rect 427862 63688 437202 63744
rect 437258 63688 437263 63744
rect 427862 63686 437263 63688
rect 427862 63610 427922 63686
rect 437197 63683 437263 63686
rect 437473 63746 437539 63749
rect 456517 63746 456583 63749
rect 437473 63744 444298 63746
rect 437473 63688 437478 63744
rect 437534 63688 444298 63744
rect 437473 63686 444298 63688
rect 437473 63683 437539 63686
rect 424918 63550 427922 63610
rect 444238 63610 444298 63686
rect 447182 63744 456583 63746
rect 447182 63688 456522 63744
rect 456578 63688 456583 63744
rect 447182 63686 456583 63688
rect 447182 63610 447242 63686
rect 456517 63683 456583 63686
rect 456885 63746 456951 63749
rect 456885 63744 466378 63746
rect 456885 63688 456890 63744
rect 456946 63688 466378 63744
rect 456885 63686 466378 63688
rect 456885 63683 456951 63686
rect 444238 63550 447242 63610
rect 466318 63610 466378 63686
rect 470550 63610 470610 63822
rect 466318 63550 470610 63610
rect 480118 63610 480178 63822
rect 480302 63822 489930 63882
rect 480302 63610 480362 63822
rect 489870 63746 489930 63822
rect 499622 63822 509250 63882
rect 489870 63686 499498 63746
rect 480118 63550 480362 63610
rect 499438 63610 499498 63686
rect 499622 63610 499682 63822
rect 509190 63746 509250 63822
rect 518942 63822 528570 63882
rect 509190 63686 518818 63746
rect 499438 63550 499682 63610
rect 518758 63610 518818 63686
rect 518942 63610 519002 63822
rect 528510 63746 528570 63822
rect 538262 63822 547890 63882
rect 528510 63686 538138 63746
rect 518758 63550 519002 63610
rect 538078 63610 538138 63686
rect 538262 63610 538322 63822
rect 547830 63746 547890 63822
rect 557582 63822 567210 63882
rect 547830 63686 557458 63746
rect 538078 63550 538322 63610
rect 557398 63610 557458 63686
rect 557582 63610 557642 63822
rect 567150 63746 567210 63822
rect 583342 63746 583402 64502
rect 583520 64412 584960 64502
rect 567150 63686 576778 63746
rect 557398 63550 557642 63610
rect 576718 63610 576778 63686
rect 576902 63686 583402 63746
rect 576902 63610 576962 63686
rect 576718 63550 576962 63610
rect 405660 63548 405666 63550
rect 289997 60754 290063 60757
rect 290181 60754 290247 60757
rect 289997 60752 290247 60754
rect 289997 60696 290002 60752
rect 290058 60696 290186 60752
rect 290242 60696 290247 60752
rect 289997 60694 290247 60696
rect 289997 60691 290063 60694
rect 290181 60691 290247 60694
rect 286041 56674 286107 56677
rect 286225 56674 286291 56677
rect 286041 56672 286291 56674
rect 286041 56616 286046 56672
rect 286102 56616 286230 56672
rect 286286 56616 286291 56672
rect 286041 56614 286291 56616
rect 286041 56611 286107 56614
rect 286225 56611 286291 56614
rect 393497 55178 393563 55181
rect 393681 55178 393747 55181
rect 393497 55176 393747 55178
rect 393497 55120 393502 55176
rect 393558 55120 393686 55176
rect 393742 55120 393747 55176
rect 393497 55118 393747 55120
rect 393497 55115 393563 55118
rect 393681 55115 393747 55118
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 2773 50146 2839 50149
rect -960 50144 2839 50146
rect -960 50088 2778 50144
rect 2834 50088 2839 50144
rect -960 50086 2839 50088
rect -960 49996 480 50086
rect 2773 50083 2839 50086
rect 366909 48514 366975 48517
rect 366909 48512 367018 48514
rect 366909 48456 366914 48512
rect 366970 48456 367018 48512
rect 366909 48451 367018 48456
rect 366958 48381 367018 48451
rect 245929 48378 245995 48381
rect 245702 48376 245995 48378
rect 245702 48320 245934 48376
rect 245990 48320 245995 48376
rect 245702 48318 245995 48320
rect 245561 48242 245627 48245
rect 245702 48242 245762 48318
rect 245929 48315 245995 48318
rect 267733 48378 267799 48381
rect 330293 48378 330359 48381
rect 331581 48378 331647 48381
rect 267733 48376 267842 48378
rect 267733 48320 267738 48376
rect 267794 48320 267842 48376
rect 267733 48315 267842 48320
rect 245561 48240 245762 48242
rect 245561 48184 245566 48240
rect 245622 48184 245762 48240
rect 245561 48182 245762 48184
rect 267782 48242 267842 48315
rect 329974 48376 330359 48378
rect 329974 48320 330298 48376
rect 330354 48320 330359 48376
rect 329974 48318 330359 48320
rect 329974 48245 330034 48318
rect 330293 48315 330359 48318
rect 331262 48376 331647 48378
rect 331262 48320 331586 48376
rect 331642 48320 331647 48376
rect 331262 48318 331647 48320
rect 267917 48242 267983 48245
rect 267782 48240 267983 48242
rect 267782 48184 267922 48240
rect 267978 48184 267983 48240
rect 267782 48182 267983 48184
rect 245561 48179 245627 48182
rect 267917 48179 267983 48182
rect 329925 48240 330034 48245
rect 329925 48184 329930 48240
rect 329986 48184 330034 48240
rect 329925 48182 330034 48184
rect 331121 48242 331187 48245
rect 331262 48242 331322 48318
rect 331581 48315 331647 48318
rect 366909 48376 367018 48381
rect 366909 48320 366914 48376
rect 366970 48320 367018 48376
rect 366909 48318 367018 48320
rect 366909 48315 366975 48318
rect 331121 48240 331322 48242
rect 331121 48184 331126 48240
rect 331182 48184 331322 48240
rect 331121 48182 331322 48184
rect 329925 48179 329991 48182
rect 331121 48179 331187 48182
rect 303981 45794 304047 45797
rect 303662 45792 304047 45794
rect 303662 45736 303986 45792
rect 304042 45736 304047 45792
rect 303662 45734 304047 45736
rect 303662 45658 303722 45734
rect 303981 45731 304047 45734
rect 303797 45658 303863 45661
rect 303662 45656 303863 45658
rect 303662 45600 303802 45656
rect 303858 45600 303863 45656
rect 303662 45598 303863 45600
rect 303797 45595 303863 45598
rect 294086 45460 294092 45524
rect 294156 45522 294162 45524
rect 294229 45522 294295 45525
rect 294156 45520 294295 45522
rect 294156 45464 294234 45520
rect 294290 45464 294295 45520
rect 294156 45462 294295 45464
rect 294156 45460 294162 45462
rect 294229 45459 294295 45462
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 396030 40430 405658 40490
rect 270542 40294 275570 40354
rect 270401 40218 270467 40221
rect 270542 40218 270602 40294
rect 234662 40158 254042 40218
rect 232998 40020 233004 40084
rect 233068 40082 233074 40084
rect 234662 40082 234722 40158
rect 233068 40022 234722 40082
rect 253982 40082 254042 40158
rect 270401 40216 270602 40218
rect 270401 40160 270406 40216
rect 270462 40160 270602 40216
rect 270401 40158 270602 40160
rect 275510 40218 275570 40294
rect 331078 40294 340890 40354
rect 275510 40158 312002 40218
rect 270401 40155 270467 40158
rect 270401 40082 270467 40085
rect 253982 40080 270467 40082
rect 253982 40024 270406 40080
rect 270462 40024 270467 40080
rect 253982 40022 270467 40024
rect 311942 40082 312002 40158
rect 331078 40082 331138 40294
rect 311942 40022 331138 40082
rect 340830 40082 340890 40294
rect 369902 40294 389834 40354
rect 360101 40218 360167 40221
rect 350582 40216 360167 40218
rect 350582 40160 360106 40216
rect 360162 40160 360167 40216
rect 350582 40158 360167 40160
rect 350582 40082 350642 40158
rect 360101 40155 360167 40158
rect 360285 40218 360351 40221
rect 360285 40216 369778 40218
rect 360285 40160 360290 40216
rect 360346 40160 369778 40216
rect 360285 40158 369778 40160
rect 360285 40155 360351 40158
rect 340830 40022 350642 40082
rect 369718 40082 369778 40158
rect 369902 40082 369962 40294
rect 389774 40218 389834 40294
rect 396030 40218 396090 40430
rect 405598 40356 405658 40430
rect 405590 40292 405596 40356
rect 405660 40292 405666 40356
rect 470550 40294 480178 40354
rect 417877 40218 417943 40221
rect 389774 40158 396090 40218
rect 408542 40216 417943 40218
rect 408542 40160 417882 40216
rect 417938 40160 417943 40216
rect 408542 40158 417943 40160
rect 369718 40022 369962 40082
rect 233068 40020 233074 40022
rect 270401 40019 270467 40022
rect 405590 40020 405596 40084
rect 405660 40082 405666 40084
rect 408542 40082 408602 40158
rect 417877 40155 417943 40158
rect 418153 40218 418219 40221
rect 437197 40218 437263 40221
rect 418153 40216 424978 40218
rect 418153 40160 418158 40216
rect 418214 40160 424978 40216
rect 418153 40158 424978 40160
rect 418153 40155 418219 40158
rect 405660 40022 408602 40082
rect 424918 40082 424978 40158
rect 427862 40216 437263 40218
rect 427862 40160 437202 40216
rect 437258 40160 437263 40216
rect 427862 40158 437263 40160
rect 427862 40082 427922 40158
rect 437197 40155 437263 40158
rect 437565 40218 437631 40221
rect 456517 40218 456583 40221
rect 437565 40216 444298 40218
rect 437565 40160 437570 40216
rect 437626 40160 444298 40216
rect 437565 40158 444298 40160
rect 437565 40155 437631 40158
rect 424918 40022 427922 40082
rect 444238 40082 444298 40158
rect 447182 40216 456583 40218
rect 447182 40160 456522 40216
rect 456578 40160 456583 40216
rect 447182 40158 456583 40160
rect 447182 40082 447242 40158
rect 456517 40155 456583 40158
rect 456885 40218 456951 40221
rect 456885 40216 466378 40218
rect 456885 40160 456890 40216
rect 456946 40160 466378 40216
rect 456885 40158 466378 40160
rect 456885 40155 456951 40158
rect 444238 40022 447242 40082
rect 466318 40082 466378 40158
rect 470550 40082 470610 40294
rect 466318 40022 470610 40082
rect 480118 40082 480178 40294
rect 480302 40294 489930 40354
rect 480302 40082 480362 40294
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 480118 40022 480362 40082
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576902 40158 583402 40218
rect 576902 40082 576962 40158
rect 576718 40022 576962 40082
rect 405660 40020 405666 40022
rect 393405 37362 393471 37365
rect 393589 37362 393655 37365
rect 393405 37360 393655 37362
rect 393405 37304 393410 37360
rect 393466 37304 393594 37360
rect 393650 37304 393655 37360
rect 393405 37302 393655 37304
rect 393405 37299 393471 37302
rect 393589 37299 393655 37302
rect 294137 36004 294203 36005
rect -960 35866 480 35956
rect 294086 35940 294092 36004
rect 294156 36002 294203 36004
rect 294156 36000 294248 36002
rect 294198 35944 294248 36000
rect 294156 35942 294248 35944
rect 294156 35940 294203 35942
rect 294137 35939 294203 35940
rect 3141 35866 3207 35869
rect -960 35864 3207 35866
rect -960 35808 3146 35864
rect 3202 35808 3207 35864
rect -960 35806 3207 35808
rect -960 35716 480 35806
rect 3141 35803 3207 35806
rect 405590 29474 405596 29476
rect 398606 29414 405596 29474
rect 235758 29276 235764 29340
rect 235828 29338 235834 29340
rect 253105 29338 253171 29341
rect 326981 29340 327047 29341
rect 326981 29338 327028 29340
rect 235828 29336 253171 29338
rect 235828 29280 253110 29336
rect 253166 29280 253171 29336
rect 235828 29278 253171 29280
rect 235828 29276 235834 29278
rect 253105 29275 253171 29278
rect 273854 29278 278882 29338
rect 326940 29336 327028 29338
rect 326940 29280 326986 29336
rect 326940 29278 327028 29280
rect 257981 29202 258047 29205
rect 273069 29202 273135 29205
rect 257981 29200 273135 29202
rect 257981 29144 257986 29200
rect 258042 29144 273074 29200
rect 273130 29144 273135 29200
rect 257981 29142 273135 29144
rect 257981 29139 258047 29142
rect 273069 29139 273135 29142
rect 273253 29202 273319 29205
rect 273854 29202 273914 29278
rect 273253 29200 273914 29202
rect 273253 29144 273258 29200
rect 273314 29144 273914 29200
rect 273253 29142 273914 29144
rect 278822 29202 278882 29278
rect 326981 29276 327028 29278
rect 327092 29276 327098 29340
rect 336641 29338 336707 29341
rect 336641 29336 340890 29338
rect 336641 29280 336646 29336
rect 336702 29280 340890 29336
rect 336641 29278 340890 29280
rect 326981 29275 327047 29276
rect 336641 29275 336707 29278
rect 287094 29202 287100 29204
rect 278822 29142 287100 29202
rect 273253 29139 273319 29142
rect 287094 29140 287100 29142
rect 287164 29140 287170 29204
rect 325601 29202 325667 29205
rect 316174 29200 325667 29202
rect 316174 29144 325606 29200
rect 325662 29144 325667 29200
rect 316174 29142 325667 29144
rect 316174 28964 316234 29142
rect 325601 29139 325667 29142
rect 327022 29004 327028 29068
rect 327092 29066 327098 29068
rect 336641 29066 336707 29069
rect 327092 29064 336707 29066
rect 327092 29008 336646 29064
rect 336702 29008 336707 29064
rect 327092 29006 336707 29008
rect 340830 29066 340890 29278
rect 367142 29278 379530 29338
rect 367142 29205 367202 29278
rect 350582 29142 362234 29202
rect 350582 29066 350642 29142
rect 340830 29006 350642 29066
rect 362174 29066 362234 29142
rect 367093 29200 367202 29205
rect 367093 29144 367098 29200
rect 367154 29144 367202 29200
rect 367093 29142 367202 29144
rect 367093 29139 367159 29142
rect 367093 29066 367159 29069
rect 362174 29064 367159 29066
rect 362174 29008 367098 29064
rect 367154 29008 367159 29064
rect 362174 29006 367159 29008
rect 379470 29066 379530 29278
rect 398606 29202 398666 29414
rect 405590 29412 405596 29414
rect 405660 29412 405666 29476
rect 481582 29412 481588 29476
rect 481652 29474 481658 29476
rect 491201 29474 491267 29477
rect 481652 29472 491267 29474
rect 481652 29416 491206 29472
rect 491262 29416 491267 29472
rect 481652 29414 491267 29416
rect 481652 29412 481658 29414
rect 491201 29411 491267 29414
rect 467925 29338 467991 29341
rect 476021 29338 476087 29341
rect 447182 29278 463618 29338
rect 417877 29202 417943 29205
rect 389222 29142 398666 29202
rect 408542 29200 417943 29202
rect 408542 29144 417882 29200
rect 417938 29144 417943 29200
rect 408542 29142 417943 29144
rect 389222 29066 389282 29142
rect 379470 29006 389282 29066
rect 327092 29004 327098 29006
rect 336641 29003 336707 29006
rect 367093 29003 367159 29006
rect 405590 29004 405596 29068
rect 405660 29066 405666 29068
rect 408542 29066 408602 29142
rect 417877 29139 417943 29142
rect 418153 29202 418219 29205
rect 437197 29202 437263 29205
rect 418153 29200 424978 29202
rect 418153 29144 418158 29200
rect 418214 29144 424978 29200
rect 418153 29142 424978 29144
rect 418153 29139 418219 29142
rect 405660 29006 408602 29066
rect 424918 29066 424978 29142
rect 427862 29200 437263 29202
rect 427862 29144 437202 29200
rect 437258 29144 437263 29200
rect 427862 29142 437263 29144
rect 427862 29066 427922 29142
rect 437197 29139 437263 29142
rect 437473 29202 437539 29205
rect 437473 29200 444298 29202
rect 437473 29144 437478 29200
rect 437534 29144 444298 29200
rect 437473 29142 444298 29144
rect 437473 29139 437539 29142
rect 424918 29006 427922 29066
rect 444238 29066 444298 29142
rect 447182 29066 447242 29278
rect 463558 29202 463618 29278
rect 467925 29336 476087 29338
rect 467925 29280 467930 29336
rect 467986 29280 476026 29336
rect 476082 29280 476087 29336
rect 467925 29278 476087 29280
rect 467925 29275 467991 29278
rect 476021 29275 476087 29278
rect 502241 29338 502307 29341
rect 583520 29338 584960 29428
rect 502241 29336 509250 29338
rect 502241 29280 502246 29336
rect 502302 29280 509250 29336
rect 502241 29278 509250 29280
rect 502241 29275 502307 29278
rect 465257 29202 465323 29205
rect 463558 29200 465323 29202
rect 463558 29144 465262 29200
rect 465318 29144 465323 29200
rect 463558 29142 465323 29144
rect 465257 29139 465323 29142
rect 476205 29202 476271 29205
rect 481582 29202 481588 29204
rect 476205 29200 481588 29202
rect 476205 29144 476210 29200
rect 476266 29144 481588 29200
rect 476205 29142 481588 29144
rect 476205 29139 476271 29142
rect 481582 29140 481588 29142
rect 481652 29140 481658 29204
rect 509190 29202 509250 29278
rect 518942 29278 528570 29338
rect 509190 29142 518818 29202
rect 444238 29006 447242 29066
rect 491201 29066 491267 29069
rect 492765 29066 492831 29069
rect 491201 29064 492831 29066
rect 491201 29008 491206 29064
rect 491262 29008 492770 29064
rect 492826 29008 492831 29064
rect 491201 29006 492831 29008
rect 518758 29066 518818 29142
rect 518942 29066 519002 29278
rect 528510 29202 528570 29278
rect 538262 29278 547890 29338
rect 528510 29142 538138 29202
rect 518758 29006 519002 29066
rect 538078 29066 538138 29142
rect 538262 29066 538322 29278
rect 547830 29202 547890 29278
rect 557582 29278 567210 29338
rect 547830 29142 557458 29202
rect 538078 29006 538322 29066
rect 557398 29066 557458 29142
rect 557582 29066 557642 29278
rect 567150 29202 567210 29278
rect 583342 29278 584960 29338
rect 583342 29202 583402 29278
rect 567150 29142 576778 29202
rect 557398 29006 557642 29066
rect 576718 29066 576778 29142
rect 576902 29142 583402 29202
rect 583520 29188 584960 29278
rect 576902 29066 576962 29142
rect 576718 29006 576962 29066
rect 405660 29004 405666 29006
rect 491201 29003 491267 29006
rect 492765 29003 492831 29006
rect 287278 28868 287284 28932
rect 287348 28930 287354 28932
rect 306281 28930 306347 28933
rect 287348 28928 306347 28930
rect 287348 28872 306286 28928
rect 306342 28872 306347 28928
rect 287348 28870 306347 28872
rect 287348 28868 287354 28870
rect 306281 28867 306347 28870
rect 314561 28930 314627 28933
rect 315990 28930 316234 28964
rect 314561 28928 316234 28930
rect 314561 28872 314566 28928
rect 314622 28904 316234 28928
rect 325601 28930 325667 28933
rect 326981 28930 327047 28933
rect 325601 28928 327047 28930
rect 314622 28872 316050 28904
rect 314561 28870 316050 28872
rect 325601 28872 325606 28928
rect 325662 28872 326986 28928
rect 327042 28872 327047 28928
rect 325601 28870 327047 28872
rect 314561 28867 314627 28870
rect 325601 28867 325667 28870
rect 326981 28867 327047 28870
rect 341149 28930 341215 28933
rect 341333 28930 341399 28933
rect 341149 28928 341399 28930
rect 341149 28872 341154 28928
rect 341210 28872 341338 28928
rect 341394 28872 341399 28928
rect 341149 28870 341399 28872
rect 341149 28867 341215 28870
rect 341333 28867 341399 28870
rect 331489 27842 331555 27845
rect 331262 27840 331555 27842
rect 331262 27784 331494 27840
rect 331550 27784 331555 27840
rect 331262 27782 331555 27784
rect 331262 27706 331322 27782
rect 331489 27779 331555 27782
rect 331397 27706 331463 27709
rect 331262 27704 331463 27706
rect 331262 27648 331402 27704
rect 331458 27648 331463 27704
rect 331262 27646 331463 27648
rect 331397 27643 331463 27646
rect 306649 24850 306715 24853
rect 307017 24850 307083 24853
rect 306649 24848 307083 24850
rect 306649 24792 306654 24848
rect 306710 24792 307022 24848
rect 307078 24792 307083 24848
rect 306649 24790 307083 24792
rect 306649 24787 306715 24790
rect 307017 24787 307083 24790
rect 467782 21994 467788 21996
rect 614 21934 467788 21994
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 467782 21932 467788 21934
rect 467852 21932 467858 21996
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 251357 19274 251423 19277
rect 251222 19272 251423 19274
rect 251222 19216 251362 19272
rect 251418 19216 251423 19272
rect 251222 19214 251423 19216
rect 251222 19138 251282 19214
rect 251357 19211 251423 19214
rect 251633 19138 251699 19141
rect 251222 19136 251699 19138
rect 251222 19080 251638 19136
rect 251694 19080 251699 19136
rect 251222 19078 251699 19080
rect 251633 19075 251699 19078
rect 583520 17642 584960 17732
rect 583342 17582 584960 17642
rect 473302 17172 473308 17236
rect 473372 17234 473378 17236
rect 482921 17234 482987 17237
rect 473372 17232 482987 17234
rect 473372 17176 482926 17232
rect 482982 17176 482987 17232
rect 473372 17174 482987 17176
rect 473372 17172 473378 17174
rect 482921 17171 482987 17174
rect 311157 17098 311223 17101
rect 317321 17098 317387 17101
rect 336641 17098 336707 17101
rect 405406 17098 405412 17100
rect 311157 17096 317387 17098
rect 311157 17040 311162 17096
rect 311218 17040 317326 17096
rect 317382 17040 317387 17096
rect 311157 17038 317387 17040
rect 311157 17035 311223 17038
rect 317321 17035 317387 17038
rect 327030 17096 336707 17098
rect 327030 17040 336646 17096
rect 336702 17040 336707 17096
rect 327030 17038 336707 17040
rect 265617 16962 265683 16965
rect 288341 16962 288407 16965
rect 265617 16960 270418 16962
rect 265617 16904 265622 16960
rect 265678 16904 270418 16960
rect 265617 16902 270418 16904
rect 265617 16899 265683 16902
rect 231710 16764 231716 16828
rect 231780 16826 231786 16828
rect 231780 16766 245026 16826
rect 231780 16764 231786 16766
rect 244966 16690 245026 16766
rect 244966 16630 249994 16690
rect 249934 16418 249994 16630
rect 270358 16554 270418 16902
rect 288341 16960 289738 16962
rect 288341 16904 288346 16960
rect 288402 16904 289738 16960
rect 288341 16902 289738 16904
rect 288341 16899 288407 16902
rect 288341 16826 288407 16829
rect 278822 16824 288407 16826
rect 278822 16768 288346 16824
rect 288402 16768 288407 16824
rect 278822 16766 288407 16768
rect 289678 16826 289738 16902
rect 299381 16826 299447 16829
rect 289678 16824 299447 16826
rect 289678 16768 299386 16824
rect 299442 16768 299447 16824
rect 289678 16766 299447 16768
rect 278822 16690 278882 16766
rect 288341 16763 288407 16766
rect 299381 16763 299447 16766
rect 322197 16826 322263 16829
rect 327030 16826 327090 17038
rect 336641 17035 336707 17038
rect 398606 17038 405412 17098
rect 322197 16824 327090 16826
rect 322197 16768 322202 16824
rect 322258 16768 327090 16824
rect 322197 16766 327090 16768
rect 340830 16902 360210 16962
rect 322197 16763 322263 16766
rect 273302 16630 278882 16690
rect 317321 16690 317387 16693
rect 336641 16690 336707 16693
rect 340830 16690 340890 16902
rect 360150 16826 360210 16902
rect 398606 16826 398666 17038
rect 405406 17036 405412 17038
rect 405476 17036 405482 17100
rect 463366 17098 463372 17100
rect 456566 17038 463372 17098
rect 417877 16826 417943 16829
rect 360150 16766 369778 16826
rect 317321 16688 317522 16690
rect 317321 16632 317326 16688
rect 317382 16632 317522 16688
rect 317321 16630 317522 16632
rect 273302 16554 273362 16630
rect 317321 16627 317387 16630
rect 270358 16494 273362 16554
rect 265617 16418 265683 16421
rect 249934 16416 265683 16418
rect 249934 16360 265622 16416
rect 265678 16360 265683 16416
rect 249934 16358 265683 16360
rect 317462 16418 317522 16630
rect 336641 16688 340890 16690
rect 336641 16632 336646 16688
rect 336702 16632 340890 16688
rect 336641 16630 340890 16632
rect 369718 16690 369778 16766
rect 388486 16766 398666 16826
rect 408542 16824 417943 16826
rect 408542 16768 417882 16824
rect 417938 16768 417943 16824
rect 408542 16766 417943 16768
rect 388486 16690 388546 16766
rect 369718 16630 388546 16690
rect 336641 16627 336707 16630
rect 405590 16628 405596 16692
rect 405660 16690 405666 16692
rect 408542 16690 408602 16766
rect 417877 16763 417943 16766
rect 418153 16826 418219 16829
rect 437197 16826 437263 16829
rect 418153 16824 424978 16826
rect 418153 16768 418158 16824
rect 418214 16768 424978 16824
rect 418153 16766 424978 16768
rect 418153 16763 418219 16766
rect 405660 16630 408602 16690
rect 424918 16690 424978 16766
rect 427862 16824 437263 16826
rect 427862 16768 437202 16824
rect 437258 16768 437263 16824
rect 427862 16766 437263 16768
rect 427862 16690 427922 16766
rect 437197 16763 437263 16766
rect 437473 16826 437539 16829
rect 456566 16826 456626 17038
rect 463366 17036 463372 17038
rect 463436 17036 463442 17100
rect 487797 17098 487863 17101
rect 483062 17096 487863 17098
rect 483062 17040 487802 17096
rect 487858 17040 487863 17096
rect 483062 17038 487863 17040
rect 466545 16962 466611 16965
rect 473302 16962 473308 16964
rect 466545 16960 473308 16962
rect 466545 16904 466550 16960
rect 466606 16904 473308 16960
rect 466545 16902 473308 16904
rect 466545 16899 466611 16902
rect 473302 16900 473308 16902
rect 473372 16900 473378 16964
rect 437473 16824 444298 16826
rect 437473 16768 437478 16824
rect 437534 16768 444298 16824
rect 437473 16766 444298 16768
rect 437473 16763 437539 16766
rect 424918 16630 427922 16690
rect 444238 16690 444298 16766
rect 447182 16766 456626 16826
rect 482921 16826 482987 16829
rect 483062 16826 483122 17038
rect 487797 17035 487863 17038
rect 492622 16900 492628 16964
rect 492692 16962 492698 16964
rect 492692 16902 509250 16962
rect 492692 16900 492698 16902
rect 482921 16824 483122 16826
rect 482921 16768 482926 16824
rect 482982 16768 483122 16824
rect 482921 16766 483122 16768
rect 509190 16826 509250 16902
rect 518942 16902 528570 16962
rect 509190 16766 518818 16826
rect 447182 16690 447242 16766
rect 482921 16763 482987 16766
rect 444238 16630 447242 16690
rect 405660 16628 405666 16630
rect 463550 16628 463556 16692
rect 463620 16690 463626 16692
rect 463785 16690 463851 16693
rect 463620 16688 463851 16690
rect 463620 16632 463790 16688
rect 463846 16632 463851 16688
rect 463620 16630 463851 16632
rect 463620 16628 463626 16630
rect 463785 16627 463851 16630
rect 487797 16690 487863 16693
rect 492622 16690 492628 16692
rect 487797 16688 492628 16690
rect 487797 16632 487802 16688
rect 487858 16632 492628 16688
rect 487797 16630 492628 16632
rect 487797 16627 487863 16630
rect 492622 16628 492628 16630
rect 492692 16628 492698 16692
rect 518758 16690 518818 16766
rect 518942 16690 519002 16902
rect 528510 16826 528570 16902
rect 538262 16902 547890 16962
rect 528510 16766 538138 16826
rect 518758 16630 519002 16690
rect 538078 16690 538138 16766
rect 538262 16690 538322 16902
rect 547830 16826 547890 16902
rect 557582 16902 567210 16962
rect 547830 16766 557458 16826
rect 538078 16630 538322 16690
rect 557398 16690 557458 16766
rect 557582 16690 557642 16902
rect 567150 16826 567210 16902
rect 583342 16826 583402 17582
rect 583520 17492 584960 17582
rect 567150 16766 576778 16826
rect 557398 16630 557642 16690
rect 576718 16690 576778 16766
rect 576902 16766 583402 16826
rect 576902 16690 576962 16766
rect 576718 16630 576962 16690
rect 389357 16554 389423 16557
rect 389541 16554 389607 16557
rect 389357 16552 389607 16554
rect 389357 16496 389362 16552
rect 389418 16496 389546 16552
rect 389602 16496 389607 16552
rect 389357 16494 389607 16496
rect 389357 16491 389423 16494
rect 389541 16491 389607 16494
rect 322197 16418 322263 16421
rect 317462 16416 322263 16418
rect 317462 16360 322202 16416
rect 322258 16360 322263 16416
rect 317462 16358 322263 16360
rect 265617 16355 265683 16358
rect 322197 16355 322263 16358
rect 3141 11658 3207 11661
rect 466494 11658 466500 11660
rect 3141 11656 466500 11658
rect 3141 11600 3146 11656
rect 3202 11600 466500 11656
rect 3141 11598 466500 11600
rect 3141 11595 3207 11598
rect 466494 11596 466500 11598
rect 466564 11596 466570 11660
rect 251449 9754 251515 9757
rect 251633 9754 251699 9757
rect 251449 9752 251699 9754
rect 251449 9696 251454 9752
rect 251510 9696 251638 9752
rect 251694 9696 251699 9752
rect 251449 9694 251699 9696
rect 251449 9691 251515 9694
rect 251633 9691 251699 9694
rect 132585 8938 132651 8941
rect 284477 8938 284543 8941
rect 132585 8936 284543 8938
rect 132585 8880 132590 8936
rect 132646 8880 284482 8936
rect 284538 8880 284543 8936
rect 132585 8878 284543 8880
rect 132585 8875 132651 8878
rect 284477 8875 284543 8878
rect 264973 8394 265039 8397
rect 265157 8394 265223 8397
rect 264973 8392 265223 8394
rect 264973 8336 264978 8392
rect 265034 8336 265162 8392
rect 265218 8336 265223 8392
rect 264973 8334 265223 8336
rect 264973 8331 265039 8334
rect 265157 8331 265223 8334
rect 128997 7578 129063 7581
rect 283097 7578 283163 7581
rect 128997 7576 283163 7578
rect 128997 7520 129002 7576
rect 129058 7520 283102 7576
rect 283158 7520 283163 7576
rect 128997 7518 283163 7520
rect 128997 7515 129063 7518
rect 283097 7515 283163 7518
rect -960 7170 480 7260
rect 3141 7170 3207 7173
rect -960 7168 3207 7170
rect -960 7112 3146 7168
rect 3202 7112 3207 7168
rect -960 7110 3207 7112
rect -960 7020 480 7110
rect 3141 7107 3207 7110
rect 51625 6218 51691 6221
rect 249977 6218 250043 6221
rect 51625 6216 250043 6218
rect 51625 6160 51630 6216
rect 51686 6160 249982 6216
rect 250038 6160 250043 6216
rect 51625 6158 250043 6160
rect 51625 6155 51691 6158
rect 249977 6155 250043 6158
rect 583520 5796 584960 6036
rect 245745 5538 245811 5541
rect 245745 5536 245946 5538
rect 245745 5480 245750 5536
rect 245806 5480 245946 5536
rect 245745 5478 245946 5480
rect 245745 5475 245811 5478
rect 238109 5402 238175 5405
rect 245886 5402 245946 5478
rect 238109 5400 245946 5402
rect 238109 5344 238114 5400
rect 238170 5344 245946 5400
rect 238109 5342 245946 5344
rect 238109 5339 238175 5342
rect 208669 4858 208735 4861
rect 314653 4858 314719 4861
rect 208669 4856 314719 4858
rect 208669 4800 208674 4856
rect 208730 4800 314658 4856
rect 314714 4800 314719 4856
rect 208669 4798 314719 4800
rect 208669 4795 208735 4798
rect 314653 4795 314719 4798
rect 467741 4858 467807 4861
rect 576209 4858 576275 4861
rect 467741 4856 576275 4858
rect 467741 4800 467746 4856
rect 467802 4800 576214 4856
rect 576270 4800 576275 4856
rect 467741 4798 576275 4800
rect 467741 4795 467807 4798
rect 576209 4795 576275 4798
rect 6453 3362 6519 3365
rect 232037 3362 232103 3365
rect 6453 3360 232103 3362
rect 6453 3304 6458 3360
rect 6514 3304 232042 3360
rect 232098 3304 232103 3360
rect 6453 3302 232103 3304
rect 6453 3299 6519 3302
rect 232037 3299 232103 3302
rect 307385 3362 307451 3365
rect 356237 3362 356303 3365
rect 307385 3360 356303 3362
rect 307385 3304 307390 3360
rect 307446 3304 356242 3360
rect 356298 3304 356303 3360
rect 307385 3302 356303 3304
rect 307385 3299 307451 3302
rect 356237 3299 356303 3302
rect 468845 3362 468911 3365
rect 580993 3362 581059 3365
rect 468845 3360 581059 3362
rect 468845 3304 468850 3360
rect 468906 3304 580998 3360
rect 581054 3304 581059 3360
rect 468845 3302 581059 3304
rect 468845 3299 468911 3302
rect 580993 3299 581059 3302
rect 340873 3090 340939 3093
rect 345749 3090 345815 3093
rect 340873 3088 345815 3090
rect 340873 3032 340878 3088
rect 340934 3032 345754 3088
rect 345810 3032 345815 3088
rect 340873 3030 345815 3032
rect 340873 3027 340939 3030
rect 345749 3027 345815 3030
<< via3 >>
rect 465764 583204 465828 583268
rect 465580 583068 465644 583132
rect 247908 582932 247972 582996
rect 247724 582796 247788 582860
rect 247540 582660 247604 582724
rect 231716 579260 231780 579324
rect 233004 579320 233068 579324
rect 233004 579264 233018 579320
rect 233018 579264 233068 579320
rect 233004 579260 233068 579264
rect 235764 579260 235828 579324
rect 237236 579320 237300 579324
rect 237236 579264 237250 579320
rect 237250 579264 237300 579320
rect 237236 579260 237300 579264
rect 239996 579260 240060 579324
rect 241284 579260 241348 579324
rect 244044 579260 244108 579324
rect 245332 579320 245396 579324
rect 245332 579264 245382 579320
rect 245382 579264 245396 579320
rect 245332 579260 245396 579264
rect 248276 579260 248340 579324
rect 249012 579260 249076 579324
rect 466500 579320 466564 579324
rect 466500 579264 466514 579320
rect 466514 579264 466564 579320
rect 466500 579260 466564 579264
rect 467788 579260 467852 579324
rect 465764 533020 465828 533084
rect 465948 486100 466012 486164
rect 247908 337996 247972 338060
rect 251404 307668 251468 307732
rect 341380 299372 341444 299436
rect 251404 298148 251468 298212
rect 341380 289852 341444 289916
rect 341380 280060 341444 280124
rect 341380 270540 341444 270604
rect 341380 260748 341444 260812
rect 247724 252452 247788 252516
rect 341380 251228 341444 251292
rect 460060 241496 460124 241500
rect 460060 241440 460074 241496
rect 460074 241440 460124 241496
rect 460060 241436 460124 241440
rect 460060 234560 460124 234564
rect 460060 234504 460110 234560
rect 460110 234504 460124 234560
rect 460060 234500 460124 234504
rect 247172 220764 247236 220828
rect 247172 211168 247236 211172
rect 247172 211112 247222 211168
rect 247222 211112 247236 211168
rect 247172 211108 247236 211112
rect 366956 173904 367020 173908
rect 366956 173848 367006 173904
rect 367006 173848 367020 173904
rect 366956 173844 367020 173848
rect 247540 165548 247604 165612
rect 366956 164248 367020 164252
rect 366956 164192 367006 164248
rect 367006 164192 367020 164248
rect 366956 164188 367020 164192
rect 249012 157524 249076 157588
rect 405412 157796 405476 157860
rect 405596 157388 405660 157452
rect 258028 134540 258092 134604
rect 245332 134132 245396 134196
rect 258028 134132 258092 134196
rect 405596 134132 405660 134196
rect 405596 133860 405660 133924
rect 492628 134132 492692 134196
rect 492628 133860 492692 133924
rect 315988 123524 316052 123588
rect 267780 123252 267844 123316
rect 315988 123252 316052 123316
rect 248276 123116 248340 123180
rect 267780 122980 267844 123044
rect 462268 122980 462332 123044
rect 492628 123116 492692 123180
rect 492628 122844 492692 122908
rect 462268 122708 462332 122772
rect 296668 111012 296732 111076
rect 304948 111012 305012 111076
rect 315988 111012 316052 111076
rect 325740 110876 325804 110940
rect 244044 110740 244108 110804
rect 296668 110740 296732 110804
rect 304948 110740 305012 110804
rect 285628 110604 285692 110668
rect 315988 110800 316052 110804
rect 315988 110744 316002 110800
rect 316002 110744 316052 110800
rect 315988 110740 316052 110744
rect 325740 110604 325804 110668
rect 277348 110468 277412 110532
rect 357388 110604 357452 110668
rect 357572 110468 357636 110532
rect 405412 110876 405476 110940
rect 405596 110468 405660 110532
rect 462268 110604 462332 110668
rect 492628 110740 492692 110804
rect 492628 110468 492692 110532
rect 462268 110332 462332 110396
rect 277348 110196 277412 110260
rect 285628 110196 285692 110260
rect 299428 87348 299492 87412
rect 239996 87212 240060 87276
rect 299428 87076 299492 87140
rect 481588 87348 481652 87412
rect 481588 87076 481652 87140
rect 473308 76468 473372 76532
rect 299428 76196 299492 76260
rect 307708 76196 307772 76260
rect 241284 76060 241348 76124
rect 260788 75924 260852 75988
rect 260788 75652 260852 75716
rect 299428 75924 299492 75988
rect 307708 75924 307772 75988
rect 473308 76196 473372 76260
rect 492628 76196 492692 76260
rect 492628 75924 492692 75988
rect 237236 63684 237300 63748
rect 280108 63820 280172 63884
rect 288572 63684 288636 63748
rect 317276 63956 317340 64020
rect 327028 63820 327092 63884
rect 280108 63548 280172 63612
rect 288388 63548 288452 63612
rect 317276 63548 317340 63612
rect 327028 63548 327092 63612
rect 405412 63956 405476 64020
rect 405596 63548 405660 63612
rect 294092 45460 294156 45524
rect 233004 40020 233068 40084
rect 405596 40292 405660 40356
rect 405596 40020 405660 40084
rect 294092 36000 294156 36004
rect 294092 35944 294142 36000
rect 294142 35944 294156 36000
rect 294092 35940 294156 35944
rect 235764 29276 235828 29340
rect 327028 29336 327092 29340
rect 327028 29280 327042 29336
rect 327042 29280 327092 29336
rect 327028 29276 327092 29280
rect 287100 29140 287164 29204
rect 327028 29004 327092 29068
rect 405596 29412 405660 29476
rect 481588 29412 481652 29476
rect 405596 29004 405660 29068
rect 481588 29140 481652 29204
rect 287284 28868 287348 28932
rect 467788 21932 467852 21996
rect 473308 17172 473372 17236
rect 231716 16764 231780 16828
rect 405412 17036 405476 17100
rect 405596 16628 405660 16692
rect 463372 17036 463436 17100
rect 473308 16900 473372 16964
rect 492628 16900 492692 16964
rect 463556 16628 463620 16692
rect 492628 16628 492692 16692
rect 466500 11596 466564 11660
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 231715 579324 231781 579325
rect 231715 579260 231716 579324
rect 231780 579260 231781 579324
rect 231715 579259 231781 579260
rect 233003 579324 233069 579325
rect 233003 579260 233004 579324
rect 233068 579260 233069 579324
rect 233003 579259 233069 579260
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 231718 16829 231778 579259
rect 233006 40085 233066 579259
rect 234804 560454 235404 595898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 235763 579324 235829 579325
rect 235763 579260 235764 579324
rect 235828 579260 235829 579324
rect 235763 579259 235829 579260
rect 237235 579324 237301 579325
rect 237235 579260 237236 579324
rect 237300 579260 237301 579324
rect 237235 579259 237301 579260
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 233003 40084 233069 40085
rect 233003 40020 233004 40084
rect 233068 40020 233069 40084
rect 233003 40019 233069 40020
rect 234804 20454 235404 55898
rect 235766 29341 235826 579259
rect 237238 63749 237298 579259
rect 238404 564054 239004 599498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 239995 579324 240061 579325
rect 239995 579260 239996 579324
rect 240060 579260 240061 579324
rect 239995 579259 240061 579260
rect 241283 579324 241349 579325
rect 241283 579260 241284 579324
rect 241348 579260 241349 579324
rect 241283 579259 241349 579260
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 237235 63748 237301 63749
rect 237235 63684 237236 63748
rect 237300 63684 237301 63748
rect 237235 63683 237301 63684
rect 238404 60054 239004 95498
rect 239998 87277 240058 579259
rect 239995 87276 240061 87277
rect 239995 87212 239996 87276
rect 240060 87212 240061 87276
rect 239995 87211 240061 87212
rect 241286 76125 241346 579259
rect 242004 567654 242604 603098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 244043 579324 244109 579325
rect 244043 579260 244044 579324
rect 244108 579260 244109 579324
rect 244043 579259 244109 579260
rect 245331 579324 245397 579325
rect 245331 579260 245332 579324
rect 245396 579260 245397 579324
rect 245331 579259 245397 579260
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 244046 110805 244106 579259
rect 245334 134197 245394 579259
rect 245604 571254 246204 606698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 247907 582996 247973 582997
rect 247907 582932 247908 582996
rect 247972 582932 247973 582996
rect 247907 582931 247973 582932
rect 247723 582860 247789 582861
rect 247723 582796 247724 582860
rect 247788 582796 247789 582860
rect 247723 582795 247789 582796
rect 247539 582724 247605 582725
rect 247539 582660 247540 582724
rect 247604 582660 247605 582724
rect 247539 582659 247605 582660
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 247171 220828 247237 220829
rect 247171 220764 247172 220828
rect 247236 220764 247237 220828
rect 247171 220763 247237 220764
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 247174 211173 247234 220763
rect 247171 211172 247237 211173
rect 247171 211108 247172 211172
rect 247236 211108 247237 211172
rect 247171 211107 247237 211108
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 247542 165613 247602 582659
rect 247726 252517 247786 582795
rect 247910 338061 247970 582931
rect 248275 579324 248341 579325
rect 248275 579260 248276 579324
rect 248340 579260 248341 579324
rect 248275 579259 248341 579260
rect 249011 579324 249077 579325
rect 249011 579260 249012 579324
rect 249076 579260 249077 579324
rect 249011 579259 249077 579260
rect 247907 338060 247973 338061
rect 247907 337996 247908 338060
rect 247972 337996 247973 338060
rect 247907 337995 247973 337996
rect 247723 252516 247789 252517
rect 247723 252452 247724 252516
rect 247788 252452 247789 252516
rect 247723 252451 247789 252452
rect 247539 165612 247605 165613
rect 247539 165548 247540 165612
rect 247604 165548 247605 165612
rect 247539 165547 247605 165548
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245331 134196 245397 134197
rect 245331 134132 245332 134196
rect 245396 134132 245397 134196
rect 245331 134131 245397 134132
rect 244043 110804 244109 110805
rect 244043 110740 244044 110804
rect 244108 110740 244109 110804
rect 244043 110739 244109 110740
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 241283 76124 241349 76125
rect 241283 76060 241284 76124
rect 241348 76060 241349 76124
rect 241283 76059 241349 76060
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 235763 29340 235829 29341
rect 235763 29276 235764 29340
rect 235828 29276 235829 29340
rect 235763 29275 235829 29276
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 231715 16828 231781 16829
rect 231715 16764 231716 16828
rect 231780 16764 231781 16828
rect 231715 16763 231781 16764
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 103254 246204 138698
rect 248278 123181 248338 579259
rect 249014 157589 249074 579259
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 251403 307732 251469 307733
rect 251403 307668 251404 307732
rect 251468 307668 251469 307732
rect 251403 307667 251469 307668
rect 251406 298213 251466 307667
rect 251403 298212 251469 298213
rect 251403 298148 251404 298212
rect 251468 298148 251469 298212
rect 251403 298147 251469 298148
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 249011 157588 249077 157589
rect 249011 157524 249012 157588
rect 249076 157524 249077 157588
rect 249011 157523 249077 157524
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 248275 123180 248341 123181
rect 248275 123116 248276 123180
rect 248340 123116 248341 123180
rect 248275 123115 248341 123116
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 258027 134604 258093 134605
rect 258027 134540 258028 134604
rect 258092 134540 258093 134604
rect 258027 134539 258093 134540
rect 258030 134197 258090 134539
rect 258027 134196 258093 134197
rect 258027 134132 258028 134196
rect 258092 134132 258093 134196
rect 258027 134131 258093 134132
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 267779 123316 267845 123317
rect 267779 123252 267780 123316
rect 267844 123252 267845 123316
rect 267779 123251 267845 123252
rect 267782 123045 267842 123251
rect 267779 123044 267845 123045
rect 267779 122980 267780 123044
rect 267844 122980 267845 123044
rect 267779 122979 267845 122980
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 260787 75988 260853 75989
rect 260787 75924 260788 75988
rect 260852 75924 260853 75988
rect 260787 75923 260853 75924
rect 260790 75717 260850 75923
rect 260787 75716 260853 75717
rect 260787 75652 260788 75716
rect 260852 75652 260853 75716
rect 260787 75651 260853 75652
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 277347 110532 277413 110533
rect 277347 110468 277348 110532
rect 277412 110468 277413 110532
rect 277347 110467 277413 110468
rect 277350 110261 277410 110467
rect 277347 110260 277413 110261
rect 277347 110196 277348 110260
rect 277412 110196 277413 110260
rect 277347 110195 277413 110196
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 285627 110668 285693 110669
rect 285627 110604 285628 110668
rect 285692 110604 285693 110668
rect 285627 110603 285693 110604
rect 285630 110261 285690 110603
rect 288804 110454 289404 145898
rect 285627 110260 285693 110261
rect 285627 110196 285628 110260
rect 285692 110196 285693 110260
rect 285627 110195 285693 110196
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 280107 63884 280173 63885
rect 280107 63820 280108 63884
rect 280172 63820 280173 63884
rect 280107 63819 280173 63820
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 280110 63613 280170 63819
rect 280107 63612 280173 63613
rect 280107 63548 280108 63612
rect 280172 63548 280173 63612
rect 280107 63547 280173 63548
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 31254 282204 66698
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288571 63748 288637 63749
rect 288571 63684 288572 63748
rect 288636 63684 288637 63748
rect 288571 63683 288637 63684
rect 288387 63612 288453 63613
rect 288387 63548 288388 63612
rect 288452 63610 288453 63612
rect 288574 63610 288634 63683
rect 288452 63550 288634 63610
rect 288452 63548 288453 63550
rect 288387 63547 288453 63548
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 287102 29550 287346 29610
rect 287102 29205 287162 29550
rect 287099 29204 287165 29205
rect 287099 29140 287100 29204
rect 287164 29140 287165 29204
rect 287099 29139 287165 29140
rect 287286 28933 287346 29550
rect 287283 28932 287349 28933
rect 287283 28868 287284 28932
rect 287348 28868 287349 28932
rect 287283 28867 287349 28868
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 296667 111076 296733 111077
rect 296667 111012 296668 111076
rect 296732 111012 296733 111076
rect 296667 111011 296733 111012
rect 296670 110805 296730 111011
rect 296667 110804 296733 110805
rect 296667 110740 296668 110804
rect 296732 110740 296733 110804
rect 296667 110739 296733 110740
rect 299427 87412 299493 87413
rect 299427 87348 299428 87412
rect 299492 87348 299493 87412
rect 299427 87347 299493 87348
rect 299430 87141 299490 87347
rect 299427 87140 299493 87141
rect 299427 87076 299428 87140
rect 299492 87076 299493 87140
rect 299427 87075 299493 87076
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 299604 85254 300204 120698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 304947 111076 305013 111077
rect 304947 111012 304948 111076
rect 305012 111012 305013 111076
rect 304947 111011 305013 111012
rect 304950 110805 305010 111011
rect 304947 110804 305013 110805
rect 304947 110740 304948 110804
rect 305012 110740 305013 110804
rect 304947 110739 305013 110740
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299427 76260 299493 76261
rect 299427 76196 299428 76260
rect 299492 76196 299493 76260
rect 299427 76195 299493 76196
rect 299430 75989 299490 76195
rect 299427 75988 299493 75989
rect 299427 75924 299428 75988
rect 299492 75924 299493 75988
rect 299427 75923 299493 75924
rect 294091 45524 294157 45525
rect 294091 45460 294092 45524
rect 294156 45460 294157 45524
rect 294091 45459 294157 45460
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 294094 36005 294154 45459
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 294091 36004 294157 36005
rect 294091 35940 294092 36004
rect 294156 35940 294157 36004
rect 294091 35939 294157 35940
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 307707 76260 307773 76261
rect 307707 76196 307708 76260
rect 307772 76196 307773 76260
rect 307707 76195 307773 76196
rect 307710 75989 307770 76195
rect 307707 75988 307773 75989
rect 307707 75924 307708 75988
rect 307772 75924 307773 75988
rect 307707 75923 307773 75924
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 315987 123588 316053 123589
rect 315987 123524 315988 123588
rect 316052 123524 316053 123588
rect 315987 123523 316053 123524
rect 315990 123317 316050 123523
rect 315987 123316 316053 123317
rect 315987 123252 315988 123316
rect 316052 123252 316053 123316
rect 315987 123251 316053 123252
rect 315987 111076 316053 111077
rect 315987 111012 315988 111076
rect 316052 111012 316053 111076
rect 315987 111011 316053 111012
rect 315990 110805 316050 111011
rect 315987 110804 316053 110805
rect 315987 110740 315988 110804
rect 316052 110740 316053 110804
rect 315987 110739 316053 110740
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317275 64020 317341 64021
rect 317275 63956 317276 64020
rect 317340 63956 317341 64020
rect 317275 63955 317341 63956
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 317278 63613 317338 63955
rect 317275 63612 317341 63613
rect 317275 63548 317276 63612
rect 317340 63548 317341 63612
rect 317275 63547 317341 63548
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 325739 110940 325805 110941
rect 325739 110876 325740 110940
rect 325804 110876 325805 110940
rect 325739 110875 325805 110876
rect 325742 110669 325802 110875
rect 325739 110668 325805 110669
rect 325739 110604 325740 110668
rect 325804 110604 325805 110668
rect 325739 110603 325805 110604
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 327027 63884 327093 63885
rect 327027 63820 327028 63884
rect 327092 63820 327093 63884
rect 327027 63819 327093 63820
rect 327030 63613 327090 63819
rect 327027 63612 327093 63613
rect 327027 63548 327028 63612
rect 327092 63548 327093 63612
rect 327027 63547 327093 63548
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 327027 29340 327093 29341
rect 327027 29276 327028 29340
rect 327092 29276 327093 29340
rect 327027 29275 327093 29276
rect 327030 29069 327090 29275
rect 327027 29068 327093 29069
rect 327027 29004 327028 29068
rect 327092 29004 327093 29068
rect 327027 29003 327093 29004
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 341379 299436 341445 299437
rect 341379 299372 341380 299436
rect 341444 299372 341445 299436
rect 341379 299371 341445 299372
rect 341382 289917 341442 299371
rect 341379 289916 341445 289917
rect 341379 289852 341380 289916
rect 341444 289852 341445 289916
rect 341379 289851 341445 289852
rect 341379 280124 341445 280125
rect 341379 280060 341380 280124
rect 341444 280060 341445 280124
rect 341379 280059 341445 280060
rect 341382 270605 341442 280059
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 341379 270604 341445 270605
rect 341379 270540 341380 270604
rect 341444 270540 341445 270604
rect 341379 270539 341445 270540
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 341379 260812 341445 260813
rect 341379 260748 341380 260812
rect 341444 260748 341445 260812
rect 341379 260747 341445 260748
rect 341382 251293 341442 260747
rect 341379 251292 341445 251293
rect 341379 251228 341380 251292
rect 341444 251228 341445 251292
rect 341379 251227 341445 251228
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 357387 110668 357453 110669
rect 357387 110604 357388 110668
rect 357452 110604 357453 110668
rect 357387 110603 357453 110604
rect 357390 110530 357450 110603
rect 357571 110532 357637 110533
rect 357571 110530 357572 110532
rect 357390 110470 357572 110530
rect 357571 110468 357572 110470
rect 357636 110468 357637 110532
rect 357571 110467 357637 110468
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 366955 173908 367021 173909
rect 366955 173844 366956 173908
rect 367020 173844 367021 173908
rect 366955 173843 367021 173844
rect 366958 164253 367018 173843
rect 366955 164252 367021 164253
rect 366955 164188 366956 164252
rect 367020 164188 367021 164252
rect 366955 164187 367021 164188
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 405411 157860 405477 157861
rect 405411 157796 405412 157860
rect 405476 157796 405477 157860
rect 405411 157795 405477 157796
rect 405414 157450 405474 157795
rect 405595 157452 405661 157453
rect 405595 157450 405596 157452
rect 405414 157390 405596 157450
rect 405595 157388 405596 157390
rect 405660 157388 405661 157452
rect 405595 157387 405661 157388
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 405595 134196 405661 134197
rect 405595 134132 405596 134196
rect 405660 134132 405661 134196
rect 405595 134131 405661 134132
rect 405598 133925 405658 134131
rect 405595 133924 405661 133925
rect 405595 133860 405596 133924
rect 405660 133860 405661 133924
rect 405595 133859 405661 133860
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 405411 110940 405477 110941
rect 405411 110876 405412 110940
rect 405476 110876 405477 110940
rect 405411 110875 405477 110876
rect 405414 110530 405474 110875
rect 405595 110532 405661 110533
rect 405595 110530 405596 110532
rect 405414 110470 405596 110530
rect 405595 110468 405596 110470
rect 405660 110468 405661 110532
rect 405595 110467 405661 110468
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 405411 64020 405477 64021
rect 405411 63956 405412 64020
rect 405476 63956 405477 64020
rect 405411 63955 405477 63956
rect 405414 63610 405474 63955
rect 405595 63612 405661 63613
rect 405595 63610 405596 63612
rect 405414 63550 405596 63610
rect 405595 63548 405596 63550
rect 405660 63548 405661 63612
rect 405595 63547 405661 63548
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 405595 40356 405661 40357
rect 405595 40292 405596 40356
rect 405660 40292 405661 40356
rect 405595 40291 405661 40292
rect 405598 40085 405658 40291
rect 405595 40084 405661 40085
rect 405595 40020 405596 40084
rect 405660 40020 405661 40084
rect 405595 40019 405661 40020
rect 405595 29476 405661 29477
rect 405595 29412 405596 29476
rect 405660 29412 405661 29476
rect 405595 29411 405661 29412
rect 405598 29069 405658 29411
rect 405595 29068 405661 29069
rect 405595 29004 405596 29068
rect 405660 29004 405661 29068
rect 405595 29003 405661 29004
rect 405411 17100 405477 17101
rect 405411 17036 405412 17100
rect 405476 17036 405477 17100
rect 405411 17035 405477 17036
rect 405414 16690 405474 17035
rect 405595 16692 405661 16693
rect 405595 16690 405596 16692
rect 405414 16630 405596 16690
rect 405595 16628 405596 16630
rect 405660 16628 405661 16692
rect 405595 16627 405661 16628
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 465763 583268 465829 583269
rect 465763 583204 465764 583268
rect 465828 583204 465829 583268
rect 465763 583203 465829 583204
rect 465579 583132 465645 583133
rect 465579 583068 465580 583132
rect 465644 583068 465645 583132
rect 465579 583067 465645 583068
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 465582 487930 465642 583067
rect 465766 533085 465826 583203
rect 466499 579324 466565 579325
rect 466499 579260 466500 579324
rect 466564 579260 466565 579324
rect 466499 579259 466565 579260
rect 467787 579324 467853 579325
rect 467787 579260 467788 579324
rect 467852 579260 467853 579324
rect 467787 579259 467853 579260
rect 465763 533084 465829 533085
rect 465763 533020 465764 533084
rect 465828 533020 465829 533084
rect 465763 533019 465829 533020
rect 465582 487870 466010 487930
rect 465950 486165 466010 487870
rect 465947 486164 466013 486165
rect 465947 486100 465948 486164
rect 466012 486100 466013 486164
rect 465947 486099 466013 486100
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 460059 241500 460125 241501
rect 460059 241436 460060 241500
rect 460124 241436 460125 241500
rect 460059 241435 460125 241436
rect 460062 234565 460122 241435
rect 460059 234564 460125 234565
rect 460059 234500 460060 234564
rect 460124 234500 460125 234564
rect 460059 234499 460125 234500
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 462267 123044 462333 123045
rect 462267 122980 462268 123044
rect 462332 122980 462333 123044
rect 462267 122979 462333 122980
rect 462270 122773 462330 122979
rect 462267 122772 462333 122773
rect 462267 122708 462268 122772
rect 462332 122708 462333 122772
rect 462267 122707 462333 122708
rect 462267 110668 462333 110669
rect 462267 110604 462268 110668
rect 462332 110604 462333 110668
rect 462267 110603 462333 110604
rect 462270 110397 462330 110603
rect 462267 110396 462333 110397
rect 462267 110332 462268 110396
rect 462332 110332 462333 110396
rect 462267 110331 462333 110332
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 463371 17100 463437 17101
rect 463371 17036 463372 17100
rect 463436 17036 463437 17100
rect 463371 17035 463437 17036
rect 463374 16690 463434 17035
rect 463555 16692 463621 16693
rect 463555 16690 463556 16692
rect 463374 16630 463556 16690
rect 463555 16628 463556 16630
rect 463620 16628 463621 16692
rect 463555 16627 463621 16628
rect 466502 11661 466562 579259
rect 467790 21997 467850 579259
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 467787 21996 467853 21997
rect 467787 21932 467788 21996
rect 467852 21932 467853 21996
rect 467787 21931 467853 21932
rect 466499 11660 466565 11661
rect 466499 11596 466500 11660
rect 466564 11596 466565 11660
rect 466499 11595 466565 11596
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 473307 76532 473373 76533
rect 473307 76468 473308 76532
rect 473372 76468 473373 76532
rect 473307 76467 473373 76468
rect 473310 76261 473370 76467
rect 473307 76260 473373 76261
rect 473307 76196 473308 76260
rect 473372 76196 473373 76260
rect 473307 76195 473373 76196
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 473307 17236 473373 17237
rect 473307 17172 473308 17236
rect 473372 17172 473373 17236
rect 473307 17171 473373 17172
rect 473310 16965 473370 17171
rect 473307 16964 473373 16965
rect 473307 16900 473308 16964
rect 473372 16900 473373 16964
rect 473307 16899 473373 16900
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 481587 87412 481653 87413
rect 481587 87348 481588 87412
rect 481652 87348 481653 87412
rect 481587 87347 481653 87348
rect 481590 87141 481650 87347
rect 481587 87140 481653 87141
rect 481587 87076 481588 87140
rect 481652 87076 481653 87140
rect 481587 87075 481653 87076
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 481587 29476 481653 29477
rect 481587 29412 481588 29476
rect 481652 29412 481653 29476
rect 481587 29411 481653 29412
rect 481590 29205 481650 29411
rect 481587 29204 481653 29205
rect 481587 29140 481588 29204
rect 481652 29140 481653 29204
rect 481587 29139 481653 29140
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 492627 134196 492693 134197
rect 492627 134132 492628 134196
rect 492692 134132 492693 134196
rect 492627 134131 492693 134132
rect 492630 133925 492690 134131
rect 492627 133924 492693 133925
rect 492627 133860 492628 133924
rect 492692 133860 492693 133924
rect 492627 133859 492693 133860
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 492627 123180 492693 123181
rect 492627 123116 492628 123180
rect 492692 123116 492693 123180
rect 492627 123115 492693 123116
rect 492630 122909 492690 123115
rect 492627 122908 492693 122909
rect 492627 122844 492628 122908
rect 492692 122844 492693 122908
rect 492627 122843 492693 122844
rect 492627 110804 492693 110805
rect 492627 110740 492628 110804
rect 492692 110740 492693 110804
rect 492627 110739 492693 110740
rect 492630 110533 492690 110739
rect 492627 110532 492693 110533
rect 492627 110468 492628 110532
rect 492692 110468 492693 110532
rect 492627 110467 492693 110468
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 492627 76260 492693 76261
rect 492627 76196 492628 76260
rect 492692 76196 492693 76260
rect 492627 76195 492693 76196
rect 492630 75989 492690 76195
rect 492627 75988 492693 75989
rect 492627 75924 492628 75988
rect 492692 75924 492693 75988
rect 492627 75923 492693 75924
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 492627 16964 492693 16965
rect 492627 16900 492628 16964
rect 492692 16900 492693 16964
rect 492627 16899 492693 16900
rect 492630 16693 492690 16899
rect 492627 16692 492693 16693
rect 492627 16628 492628 16692
rect 492692 16628 492693 16692
rect 492627 16627 492693 16628
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use user_proj_example  mprj
timestamp 1608085893
transform 1 0 229999 0 1 340000
box 1 0 239542 240000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
