magic
tech sky130A
magscale 1 2
timestamp 1608417145
<< obsli1 >>
rect 906 1445 218670 217617
<< obsm1 >>
rect 0 1096 219576 219156
<< metal2 >>
rect 740 219200 796 220000
rect 2580 219200 2636 220000
rect 4512 219200 4568 220000
rect 6444 219200 6500 220000
rect 8376 219200 8432 220000
rect 10308 219200 10364 220000
rect 12240 219200 12296 220000
rect 14172 219200 14228 220000
rect 16104 219200 16160 220000
rect 18036 219200 18092 220000
rect 19968 219200 20024 220000
rect 21900 219200 21956 220000
rect 23832 219200 23888 220000
rect 25764 219200 25820 220000
rect 27696 219200 27752 220000
rect 29628 219200 29684 220000
rect 31560 219200 31616 220000
rect 33492 219200 33548 220000
rect 35424 219200 35480 220000
rect 37356 219200 37412 220000
rect 39288 219200 39344 220000
rect 41220 219200 41276 220000
rect 43152 219200 43208 220000
rect 45084 219200 45140 220000
rect 47016 219200 47072 220000
rect 48948 219200 49004 220000
rect 50880 219200 50936 220000
rect 52812 219200 52868 220000
rect 54744 219200 54800 220000
rect 56676 219200 56732 220000
rect 58608 219200 58664 220000
rect 60540 219200 60596 220000
rect 62472 219200 62528 220000
rect 64404 219200 64460 220000
rect 66336 219200 66392 220000
rect 68268 219200 68324 220000
rect 70200 219200 70256 220000
rect 72132 219200 72188 220000
rect 74064 219200 74120 220000
rect 75904 219200 75960 220000
rect 77836 219200 77892 220000
rect 79768 219200 79824 220000
rect 81700 219200 81756 220000
rect 83632 219200 83688 220000
rect 85564 219200 85620 220000
rect 87496 219200 87552 220000
rect 89428 219200 89484 220000
rect 91360 219200 91416 220000
rect 93292 219200 93348 220000
rect 95224 219200 95280 220000
rect 97156 219200 97212 220000
rect 99088 219200 99144 220000
rect 101020 219200 101076 220000
rect 102952 219200 103008 220000
rect 104884 219200 104940 220000
rect 106816 219200 106872 220000
rect 108748 219200 108804 220000
rect 110680 219200 110736 220000
rect 112612 219200 112668 220000
rect 114544 219200 114600 220000
rect 116476 219200 116532 220000
rect 118408 219200 118464 220000
rect 120340 219200 120396 220000
rect 122272 219200 122328 220000
rect 124204 219200 124260 220000
rect 126136 219200 126192 220000
rect 128068 219200 128124 220000
rect 130000 219200 130056 220000
rect 131932 219200 131988 220000
rect 133864 219200 133920 220000
rect 135796 219200 135852 220000
rect 137728 219200 137784 220000
rect 139660 219200 139716 220000
rect 141592 219200 141648 220000
rect 143524 219200 143580 220000
rect 145456 219200 145512 220000
rect 147388 219200 147444 220000
rect 149228 219200 149284 220000
rect 151160 219200 151216 220000
rect 153092 219200 153148 220000
rect 155024 219200 155080 220000
rect 156956 219200 157012 220000
rect 158888 219200 158944 220000
rect 160820 219200 160876 220000
rect 162752 219200 162808 220000
rect 164684 219200 164740 220000
rect 166616 219200 166672 220000
rect 168548 219200 168604 220000
rect 170480 219200 170536 220000
rect 172412 219200 172468 220000
rect 174344 219200 174400 220000
rect 176276 219200 176332 220000
rect 178208 219200 178264 220000
rect 180140 219200 180196 220000
rect 182072 219200 182128 220000
rect 184004 219200 184060 220000
rect 185936 219200 185992 220000
rect 187868 219200 187924 220000
rect 189800 219200 189856 220000
rect 191732 219200 191788 220000
rect 193664 219200 193720 220000
rect 195596 219200 195652 220000
rect 197528 219200 197584 220000
rect 199460 219200 199516 220000
rect 201392 219200 201448 220000
rect 203324 219200 203380 220000
rect 205256 219200 205312 220000
rect 207188 219200 207244 220000
rect 209120 219200 209176 220000
rect 211052 219200 211108 220000
rect 212984 219200 213040 220000
rect 214916 219200 214972 220000
rect 216848 219200 216904 220000
rect 218780 219200 218836 220000
rect 4 0 60 800
rect 372 0 428 800
rect 832 0 888 800
rect 1292 0 1348 800
rect 1752 0 1808 800
rect 2212 0 2268 800
rect 2672 0 2728 800
rect 3132 0 3188 800
rect 3592 0 3648 800
rect 3960 0 4016 800
rect 4420 0 4476 800
rect 4880 0 4936 800
rect 5340 0 5396 800
rect 5800 0 5856 800
rect 6260 0 6316 800
rect 6720 0 6776 800
rect 7180 0 7236 800
rect 7548 0 7604 800
rect 8008 0 8064 800
rect 8468 0 8524 800
rect 8928 0 8984 800
rect 9388 0 9444 800
rect 9848 0 9904 800
rect 10308 0 10364 800
rect 10768 0 10824 800
rect 11136 0 11192 800
rect 11596 0 11652 800
rect 12056 0 12112 800
rect 12516 0 12572 800
rect 12976 0 13032 800
rect 13436 0 13492 800
rect 13896 0 13952 800
rect 14356 0 14412 800
rect 14816 0 14872 800
rect 15184 0 15240 800
rect 15644 0 15700 800
rect 16104 0 16160 800
rect 16564 0 16620 800
rect 17024 0 17080 800
rect 17484 0 17540 800
rect 17944 0 18000 800
rect 18404 0 18460 800
rect 18772 0 18828 800
rect 19232 0 19288 800
rect 19692 0 19748 800
rect 20152 0 20208 800
rect 20612 0 20668 800
rect 21072 0 21128 800
rect 21532 0 21588 800
rect 21992 0 22048 800
rect 22360 0 22416 800
rect 22820 0 22876 800
rect 23280 0 23336 800
rect 23740 0 23796 800
rect 24200 0 24256 800
rect 24660 0 24716 800
rect 25120 0 25176 800
rect 25580 0 25636 800
rect 26040 0 26096 800
rect 26408 0 26464 800
rect 26868 0 26924 800
rect 27328 0 27384 800
rect 27788 0 27844 800
rect 28248 0 28304 800
rect 28708 0 28764 800
rect 29168 0 29224 800
rect 29628 0 29684 800
rect 29996 0 30052 800
rect 30456 0 30512 800
rect 30916 0 30972 800
rect 31376 0 31432 800
rect 31836 0 31892 800
rect 32296 0 32352 800
rect 32756 0 32812 800
rect 33216 0 33272 800
rect 33584 0 33640 800
rect 34044 0 34100 800
rect 34504 0 34560 800
rect 34964 0 35020 800
rect 35424 0 35480 800
rect 35884 0 35940 800
rect 36344 0 36400 800
rect 36804 0 36860 800
rect 37264 0 37320 800
rect 37632 0 37688 800
rect 38092 0 38148 800
rect 38552 0 38608 800
rect 39012 0 39068 800
rect 39472 0 39528 800
rect 39932 0 39988 800
rect 40392 0 40448 800
rect 40852 0 40908 800
rect 41220 0 41276 800
rect 41680 0 41736 800
rect 42140 0 42196 800
rect 42600 0 42656 800
rect 43060 0 43116 800
rect 43520 0 43576 800
rect 43980 0 44036 800
rect 44440 0 44496 800
rect 44808 0 44864 800
rect 45268 0 45324 800
rect 45728 0 45784 800
rect 46188 0 46244 800
rect 46648 0 46704 800
rect 47108 0 47164 800
rect 47568 0 47624 800
rect 48028 0 48084 800
rect 48396 0 48452 800
rect 48856 0 48912 800
rect 49316 0 49372 800
rect 49776 0 49832 800
rect 50236 0 50292 800
rect 50696 0 50752 800
rect 51156 0 51212 800
rect 51616 0 51672 800
rect 52076 0 52132 800
rect 52444 0 52500 800
rect 52904 0 52960 800
rect 53364 0 53420 800
rect 53824 0 53880 800
rect 54284 0 54340 800
rect 54744 0 54800 800
rect 55204 0 55260 800
rect 55664 0 55720 800
rect 56032 0 56088 800
rect 56492 0 56548 800
rect 56952 0 57008 800
rect 57412 0 57468 800
rect 57872 0 57928 800
rect 58332 0 58388 800
rect 58792 0 58848 800
rect 59252 0 59308 800
rect 59620 0 59676 800
rect 60080 0 60136 800
rect 60540 0 60596 800
rect 61000 0 61056 800
rect 61460 0 61516 800
rect 61920 0 61976 800
rect 62380 0 62436 800
rect 62840 0 62896 800
rect 63300 0 63356 800
rect 63668 0 63724 800
rect 64128 0 64184 800
rect 64588 0 64644 800
rect 65048 0 65104 800
rect 65508 0 65564 800
rect 65968 0 66024 800
rect 66428 0 66484 800
rect 66888 0 66944 800
rect 67256 0 67312 800
rect 67716 0 67772 800
rect 68176 0 68232 800
rect 68636 0 68692 800
rect 69096 0 69152 800
rect 69556 0 69612 800
rect 70016 0 70072 800
rect 70476 0 70532 800
rect 70844 0 70900 800
rect 71304 0 71360 800
rect 71764 0 71820 800
rect 72224 0 72280 800
rect 72684 0 72740 800
rect 73144 0 73200 800
rect 73604 0 73660 800
rect 74064 0 74120 800
rect 74524 0 74580 800
rect 74892 0 74948 800
rect 75352 0 75408 800
rect 75812 0 75868 800
rect 76272 0 76328 800
rect 76732 0 76788 800
rect 77192 0 77248 800
rect 77652 0 77708 800
rect 78112 0 78168 800
rect 78480 0 78536 800
rect 78940 0 78996 800
rect 79400 0 79456 800
rect 79860 0 79916 800
rect 80320 0 80376 800
rect 80780 0 80836 800
rect 81240 0 81296 800
rect 81700 0 81756 800
rect 82068 0 82124 800
rect 82528 0 82584 800
rect 82988 0 83044 800
rect 83448 0 83504 800
rect 83908 0 83964 800
rect 84368 0 84424 800
rect 84828 0 84884 800
rect 85288 0 85344 800
rect 85748 0 85804 800
rect 86116 0 86172 800
rect 86576 0 86632 800
rect 87036 0 87092 800
rect 87496 0 87552 800
rect 87956 0 88012 800
rect 88416 0 88472 800
rect 88876 0 88932 800
rect 89336 0 89392 800
rect 89704 0 89760 800
rect 90164 0 90220 800
rect 90624 0 90680 800
rect 91084 0 91140 800
rect 91544 0 91600 800
rect 92004 0 92060 800
rect 92464 0 92520 800
rect 92924 0 92980 800
rect 93292 0 93348 800
rect 93752 0 93808 800
rect 94212 0 94268 800
rect 94672 0 94728 800
rect 95132 0 95188 800
rect 95592 0 95648 800
rect 96052 0 96108 800
rect 96512 0 96568 800
rect 96880 0 96936 800
rect 97340 0 97396 800
rect 97800 0 97856 800
rect 98260 0 98316 800
rect 98720 0 98776 800
rect 99180 0 99236 800
rect 99640 0 99696 800
rect 100100 0 100156 800
rect 100560 0 100616 800
rect 100928 0 100984 800
rect 101388 0 101444 800
rect 101848 0 101904 800
rect 102308 0 102364 800
rect 102768 0 102824 800
rect 103228 0 103284 800
rect 103688 0 103744 800
rect 104148 0 104204 800
rect 104516 0 104572 800
rect 104976 0 105032 800
rect 105436 0 105492 800
rect 105896 0 105952 800
rect 106356 0 106412 800
rect 106816 0 106872 800
rect 107276 0 107332 800
rect 107736 0 107792 800
rect 108104 0 108160 800
rect 108564 0 108620 800
rect 109024 0 109080 800
rect 109484 0 109540 800
rect 109944 0 110000 800
rect 110404 0 110460 800
rect 110864 0 110920 800
rect 111324 0 111380 800
rect 111784 0 111840 800
rect 112152 0 112208 800
rect 112612 0 112668 800
rect 113072 0 113128 800
rect 113532 0 113588 800
rect 113992 0 114048 800
rect 114452 0 114508 800
rect 114912 0 114968 800
rect 115372 0 115428 800
rect 115740 0 115796 800
rect 116200 0 116256 800
rect 116660 0 116716 800
rect 117120 0 117176 800
rect 117580 0 117636 800
rect 118040 0 118096 800
rect 118500 0 118556 800
rect 118960 0 119016 800
rect 119328 0 119384 800
rect 119788 0 119844 800
rect 120248 0 120304 800
rect 120708 0 120764 800
rect 121168 0 121224 800
rect 121628 0 121684 800
rect 122088 0 122144 800
rect 122548 0 122604 800
rect 123008 0 123064 800
rect 123376 0 123432 800
rect 123836 0 123892 800
rect 124296 0 124352 800
rect 124756 0 124812 800
rect 125216 0 125272 800
rect 125676 0 125732 800
rect 126136 0 126192 800
rect 126596 0 126652 800
rect 126964 0 127020 800
rect 127424 0 127480 800
rect 127884 0 127940 800
rect 128344 0 128400 800
rect 128804 0 128860 800
rect 129264 0 129320 800
rect 129724 0 129780 800
rect 130184 0 130240 800
rect 130552 0 130608 800
rect 131012 0 131068 800
rect 131472 0 131528 800
rect 131932 0 131988 800
rect 132392 0 132448 800
rect 132852 0 132908 800
rect 133312 0 133368 800
rect 133772 0 133828 800
rect 134140 0 134196 800
rect 134600 0 134656 800
rect 135060 0 135116 800
rect 135520 0 135576 800
rect 135980 0 136036 800
rect 136440 0 136496 800
rect 136900 0 136956 800
rect 137360 0 137416 800
rect 137820 0 137876 800
rect 138188 0 138244 800
rect 138648 0 138704 800
rect 139108 0 139164 800
rect 139568 0 139624 800
rect 140028 0 140084 800
rect 140488 0 140544 800
rect 140948 0 141004 800
rect 141408 0 141464 800
rect 141776 0 141832 800
rect 142236 0 142292 800
rect 142696 0 142752 800
rect 143156 0 143212 800
rect 143616 0 143672 800
rect 144076 0 144132 800
rect 144536 0 144592 800
rect 144996 0 145052 800
rect 145364 0 145420 800
rect 145824 0 145880 800
rect 146284 0 146340 800
rect 146744 0 146800 800
rect 147204 0 147260 800
rect 147664 0 147720 800
rect 148124 0 148180 800
rect 148584 0 148640 800
rect 149044 0 149100 800
rect 149412 0 149468 800
rect 149872 0 149928 800
rect 150332 0 150388 800
rect 150792 0 150848 800
rect 151252 0 151308 800
rect 151712 0 151768 800
rect 152172 0 152228 800
rect 152632 0 152688 800
rect 153000 0 153056 800
rect 153460 0 153516 800
rect 153920 0 153976 800
rect 154380 0 154436 800
rect 154840 0 154896 800
rect 155300 0 155356 800
rect 155760 0 155816 800
rect 156220 0 156276 800
rect 156588 0 156644 800
rect 157048 0 157104 800
rect 157508 0 157564 800
rect 157968 0 158024 800
rect 158428 0 158484 800
rect 158888 0 158944 800
rect 159348 0 159404 800
rect 159808 0 159864 800
rect 160268 0 160324 800
rect 160636 0 160692 800
rect 161096 0 161152 800
rect 161556 0 161612 800
rect 162016 0 162072 800
rect 162476 0 162532 800
rect 162936 0 162992 800
rect 163396 0 163452 800
rect 163856 0 163912 800
rect 164224 0 164280 800
rect 164684 0 164740 800
rect 165144 0 165200 800
rect 165604 0 165660 800
rect 166064 0 166120 800
rect 166524 0 166580 800
rect 166984 0 167040 800
rect 167444 0 167500 800
rect 167812 0 167868 800
rect 168272 0 168328 800
rect 168732 0 168788 800
rect 169192 0 169248 800
rect 169652 0 169708 800
rect 170112 0 170168 800
rect 170572 0 170628 800
rect 171032 0 171088 800
rect 171492 0 171548 800
rect 171860 0 171916 800
rect 172320 0 172376 800
rect 172780 0 172836 800
rect 173240 0 173296 800
rect 173700 0 173756 800
rect 174160 0 174216 800
rect 174620 0 174676 800
rect 175080 0 175136 800
rect 175448 0 175504 800
rect 175908 0 175964 800
rect 176368 0 176424 800
rect 176828 0 176884 800
rect 177288 0 177344 800
rect 177748 0 177804 800
rect 178208 0 178264 800
rect 178668 0 178724 800
rect 179036 0 179092 800
rect 179496 0 179552 800
rect 179956 0 180012 800
rect 180416 0 180472 800
rect 180876 0 180932 800
rect 181336 0 181392 800
rect 181796 0 181852 800
rect 182256 0 182312 800
rect 182624 0 182680 800
rect 183084 0 183140 800
rect 183544 0 183600 800
rect 184004 0 184060 800
rect 184464 0 184520 800
rect 184924 0 184980 800
rect 185384 0 185440 800
rect 185844 0 185900 800
rect 186304 0 186360 800
rect 186672 0 186728 800
rect 187132 0 187188 800
rect 187592 0 187648 800
rect 188052 0 188108 800
rect 188512 0 188568 800
rect 188972 0 189028 800
rect 189432 0 189488 800
rect 189892 0 189948 800
rect 190260 0 190316 800
rect 190720 0 190776 800
rect 191180 0 191236 800
rect 191640 0 191696 800
rect 192100 0 192156 800
rect 192560 0 192616 800
rect 193020 0 193076 800
rect 193480 0 193536 800
rect 193848 0 193904 800
rect 194308 0 194364 800
rect 194768 0 194824 800
rect 195228 0 195284 800
rect 195688 0 195744 800
rect 196148 0 196204 800
rect 196608 0 196664 800
rect 197068 0 197124 800
rect 197528 0 197584 800
rect 197896 0 197952 800
rect 198356 0 198412 800
rect 198816 0 198872 800
rect 199276 0 199332 800
rect 199736 0 199792 800
rect 200196 0 200252 800
rect 200656 0 200712 800
rect 201116 0 201172 800
rect 201484 0 201540 800
rect 201944 0 202000 800
rect 202404 0 202460 800
rect 202864 0 202920 800
rect 203324 0 203380 800
rect 203784 0 203840 800
rect 204244 0 204300 800
rect 204704 0 204760 800
rect 205072 0 205128 800
rect 205532 0 205588 800
rect 205992 0 206048 800
rect 206452 0 206508 800
rect 206912 0 206968 800
rect 207372 0 207428 800
rect 207832 0 207888 800
rect 208292 0 208348 800
rect 208752 0 208808 800
rect 209120 0 209176 800
rect 209580 0 209636 800
rect 210040 0 210096 800
rect 210500 0 210556 800
rect 210960 0 211016 800
rect 211420 0 211476 800
rect 211880 0 211936 800
rect 212340 0 212396 800
rect 212708 0 212764 800
rect 213168 0 213224 800
rect 213628 0 213684 800
rect 214088 0 214144 800
rect 214548 0 214604 800
rect 215008 0 215064 800
rect 215468 0 215524 800
rect 215928 0 215984 800
rect 216296 0 216352 800
rect 216756 0 216812 800
rect 217216 0 217272 800
rect 217676 0 217732 800
rect 218136 0 218192 800
rect 218596 0 218652 800
rect 219056 0 219112 800
rect 219516 0 219572 800
<< obsm2 >>
rect 6 219144 684 219200
rect 852 219144 2524 219200
rect 2692 219144 4456 219200
rect 4624 219144 6388 219200
rect 6556 219144 8320 219200
rect 8488 219144 10252 219200
rect 10420 219144 12184 219200
rect 12352 219144 14116 219200
rect 14284 219144 16048 219200
rect 16216 219144 17980 219200
rect 18148 219144 19912 219200
rect 20080 219144 21844 219200
rect 22012 219144 23776 219200
rect 23944 219144 25708 219200
rect 25876 219144 27640 219200
rect 27808 219144 29572 219200
rect 29740 219144 31504 219200
rect 31672 219144 33436 219200
rect 33604 219144 35368 219200
rect 35536 219144 37300 219200
rect 37468 219144 39232 219200
rect 39400 219144 41164 219200
rect 41332 219144 43096 219200
rect 43264 219144 45028 219200
rect 45196 219144 46960 219200
rect 47128 219144 48892 219200
rect 49060 219144 50824 219200
rect 50992 219144 52756 219200
rect 52924 219144 54688 219200
rect 54856 219144 56620 219200
rect 56788 219144 58552 219200
rect 58720 219144 60484 219200
rect 60652 219144 62416 219200
rect 62584 219144 64348 219200
rect 64516 219144 66280 219200
rect 66448 219144 68212 219200
rect 68380 219144 70144 219200
rect 70312 219144 72076 219200
rect 72244 219144 74008 219200
rect 74176 219144 75848 219200
rect 76016 219144 77780 219200
rect 77948 219144 79712 219200
rect 79880 219144 81644 219200
rect 81812 219144 83576 219200
rect 83744 219144 85508 219200
rect 85676 219144 87440 219200
rect 87608 219144 89372 219200
rect 89540 219144 91304 219200
rect 91472 219144 93236 219200
rect 93404 219144 95168 219200
rect 95336 219144 97100 219200
rect 97268 219144 99032 219200
rect 99200 219144 100964 219200
rect 101132 219144 102896 219200
rect 103064 219144 104828 219200
rect 104996 219144 106760 219200
rect 106928 219144 108692 219200
rect 108860 219144 110624 219200
rect 110792 219144 112556 219200
rect 112724 219144 114488 219200
rect 114656 219144 116420 219200
rect 116588 219144 118352 219200
rect 118520 219144 120284 219200
rect 120452 219144 122216 219200
rect 122384 219144 124148 219200
rect 124316 219144 126080 219200
rect 126248 219144 128012 219200
rect 128180 219144 129944 219200
rect 130112 219144 131876 219200
rect 132044 219144 133808 219200
rect 133976 219144 135740 219200
rect 135908 219144 137672 219200
rect 137840 219144 139604 219200
rect 139772 219144 141536 219200
rect 141704 219144 143468 219200
rect 143636 219144 145400 219200
rect 145568 219144 147332 219200
rect 147500 219144 149172 219200
rect 149340 219144 151104 219200
rect 151272 219144 153036 219200
rect 153204 219144 154968 219200
rect 155136 219144 156900 219200
rect 157068 219144 158832 219200
rect 159000 219144 160764 219200
rect 160932 219144 162696 219200
rect 162864 219144 164628 219200
rect 164796 219144 166560 219200
rect 166728 219144 168492 219200
rect 168660 219144 170424 219200
rect 170592 219144 172356 219200
rect 172524 219144 174288 219200
rect 174456 219144 176220 219200
rect 176388 219144 178152 219200
rect 178320 219144 180084 219200
rect 180252 219144 182016 219200
rect 182184 219144 183948 219200
rect 184116 219144 185880 219200
rect 186048 219144 187812 219200
rect 187980 219144 189744 219200
rect 189912 219144 191676 219200
rect 191844 219144 193608 219200
rect 193776 219144 195540 219200
rect 195708 219144 197472 219200
rect 197640 219144 199404 219200
rect 199572 219144 201336 219200
rect 201504 219144 203268 219200
rect 203436 219144 205200 219200
rect 205368 219144 207132 219200
rect 207300 219144 209064 219200
rect 209232 219144 210996 219200
rect 211164 219144 212928 219200
rect 213096 219144 214860 219200
rect 215028 219144 216792 219200
rect 216960 219144 218724 219200
rect 218892 219144 219570 219200
rect 6 856 219570 219144
rect 116 800 316 856
rect 484 800 776 856
rect 944 800 1236 856
rect 1404 800 1696 856
rect 1864 800 2156 856
rect 2324 800 2616 856
rect 2784 800 3076 856
rect 3244 800 3536 856
rect 3704 800 3904 856
rect 4072 800 4364 856
rect 4532 800 4824 856
rect 4992 800 5284 856
rect 5452 800 5744 856
rect 5912 800 6204 856
rect 6372 800 6664 856
rect 6832 800 7124 856
rect 7292 800 7492 856
rect 7660 800 7952 856
rect 8120 800 8412 856
rect 8580 800 8872 856
rect 9040 800 9332 856
rect 9500 800 9792 856
rect 9960 800 10252 856
rect 10420 800 10712 856
rect 10880 800 11080 856
rect 11248 800 11540 856
rect 11708 800 12000 856
rect 12168 800 12460 856
rect 12628 800 12920 856
rect 13088 800 13380 856
rect 13548 800 13840 856
rect 14008 800 14300 856
rect 14468 800 14760 856
rect 14928 800 15128 856
rect 15296 800 15588 856
rect 15756 800 16048 856
rect 16216 800 16508 856
rect 16676 800 16968 856
rect 17136 800 17428 856
rect 17596 800 17888 856
rect 18056 800 18348 856
rect 18516 800 18716 856
rect 18884 800 19176 856
rect 19344 800 19636 856
rect 19804 800 20096 856
rect 20264 800 20556 856
rect 20724 800 21016 856
rect 21184 800 21476 856
rect 21644 800 21936 856
rect 22104 800 22304 856
rect 22472 800 22764 856
rect 22932 800 23224 856
rect 23392 800 23684 856
rect 23852 800 24144 856
rect 24312 800 24604 856
rect 24772 800 25064 856
rect 25232 800 25524 856
rect 25692 800 25984 856
rect 26152 800 26352 856
rect 26520 800 26812 856
rect 26980 800 27272 856
rect 27440 800 27732 856
rect 27900 800 28192 856
rect 28360 800 28652 856
rect 28820 800 29112 856
rect 29280 800 29572 856
rect 29740 800 29940 856
rect 30108 800 30400 856
rect 30568 800 30860 856
rect 31028 800 31320 856
rect 31488 800 31780 856
rect 31948 800 32240 856
rect 32408 800 32700 856
rect 32868 800 33160 856
rect 33328 800 33528 856
rect 33696 800 33988 856
rect 34156 800 34448 856
rect 34616 800 34908 856
rect 35076 800 35368 856
rect 35536 800 35828 856
rect 35996 800 36288 856
rect 36456 800 36748 856
rect 36916 800 37208 856
rect 37376 800 37576 856
rect 37744 800 38036 856
rect 38204 800 38496 856
rect 38664 800 38956 856
rect 39124 800 39416 856
rect 39584 800 39876 856
rect 40044 800 40336 856
rect 40504 800 40796 856
rect 40964 800 41164 856
rect 41332 800 41624 856
rect 41792 800 42084 856
rect 42252 800 42544 856
rect 42712 800 43004 856
rect 43172 800 43464 856
rect 43632 800 43924 856
rect 44092 800 44384 856
rect 44552 800 44752 856
rect 44920 800 45212 856
rect 45380 800 45672 856
rect 45840 800 46132 856
rect 46300 800 46592 856
rect 46760 800 47052 856
rect 47220 800 47512 856
rect 47680 800 47972 856
rect 48140 800 48340 856
rect 48508 800 48800 856
rect 48968 800 49260 856
rect 49428 800 49720 856
rect 49888 800 50180 856
rect 50348 800 50640 856
rect 50808 800 51100 856
rect 51268 800 51560 856
rect 51728 800 52020 856
rect 52188 800 52388 856
rect 52556 800 52848 856
rect 53016 800 53308 856
rect 53476 800 53768 856
rect 53936 800 54228 856
rect 54396 800 54688 856
rect 54856 800 55148 856
rect 55316 800 55608 856
rect 55776 800 55976 856
rect 56144 800 56436 856
rect 56604 800 56896 856
rect 57064 800 57356 856
rect 57524 800 57816 856
rect 57984 800 58276 856
rect 58444 800 58736 856
rect 58904 800 59196 856
rect 59364 800 59564 856
rect 59732 800 60024 856
rect 60192 800 60484 856
rect 60652 800 60944 856
rect 61112 800 61404 856
rect 61572 800 61864 856
rect 62032 800 62324 856
rect 62492 800 62784 856
rect 62952 800 63244 856
rect 63412 800 63612 856
rect 63780 800 64072 856
rect 64240 800 64532 856
rect 64700 800 64992 856
rect 65160 800 65452 856
rect 65620 800 65912 856
rect 66080 800 66372 856
rect 66540 800 66832 856
rect 67000 800 67200 856
rect 67368 800 67660 856
rect 67828 800 68120 856
rect 68288 800 68580 856
rect 68748 800 69040 856
rect 69208 800 69500 856
rect 69668 800 69960 856
rect 70128 800 70420 856
rect 70588 800 70788 856
rect 70956 800 71248 856
rect 71416 800 71708 856
rect 71876 800 72168 856
rect 72336 800 72628 856
rect 72796 800 73088 856
rect 73256 800 73548 856
rect 73716 800 74008 856
rect 74176 800 74468 856
rect 74636 800 74836 856
rect 75004 800 75296 856
rect 75464 800 75756 856
rect 75924 800 76216 856
rect 76384 800 76676 856
rect 76844 800 77136 856
rect 77304 800 77596 856
rect 77764 800 78056 856
rect 78224 800 78424 856
rect 78592 800 78884 856
rect 79052 800 79344 856
rect 79512 800 79804 856
rect 79972 800 80264 856
rect 80432 800 80724 856
rect 80892 800 81184 856
rect 81352 800 81644 856
rect 81812 800 82012 856
rect 82180 800 82472 856
rect 82640 800 82932 856
rect 83100 800 83392 856
rect 83560 800 83852 856
rect 84020 800 84312 856
rect 84480 800 84772 856
rect 84940 800 85232 856
rect 85400 800 85692 856
rect 85860 800 86060 856
rect 86228 800 86520 856
rect 86688 800 86980 856
rect 87148 800 87440 856
rect 87608 800 87900 856
rect 88068 800 88360 856
rect 88528 800 88820 856
rect 88988 800 89280 856
rect 89448 800 89648 856
rect 89816 800 90108 856
rect 90276 800 90568 856
rect 90736 800 91028 856
rect 91196 800 91488 856
rect 91656 800 91948 856
rect 92116 800 92408 856
rect 92576 800 92868 856
rect 93036 800 93236 856
rect 93404 800 93696 856
rect 93864 800 94156 856
rect 94324 800 94616 856
rect 94784 800 95076 856
rect 95244 800 95536 856
rect 95704 800 95996 856
rect 96164 800 96456 856
rect 96624 800 96824 856
rect 96992 800 97284 856
rect 97452 800 97744 856
rect 97912 800 98204 856
rect 98372 800 98664 856
rect 98832 800 99124 856
rect 99292 800 99584 856
rect 99752 800 100044 856
rect 100212 800 100504 856
rect 100672 800 100872 856
rect 101040 800 101332 856
rect 101500 800 101792 856
rect 101960 800 102252 856
rect 102420 800 102712 856
rect 102880 800 103172 856
rect 103340 800 103632 856
rect 103800 800 104092 856
rect 104260 800 104460 856
rect 104628 800 104920 856
rect 105088 800 105380 856
rect 105548 800 105840 856
rect 106008 800 106300 856
rect 106468 800 106760 856
rect 106928 800 107220 856
rect 107388 800 107680 856
rect 107848 800 108048 856
rect 108216 800 108508 856
rect 108676 800 108968 856
rect 109136 800 109428 856
rect 109596 800 109888 856
rect 110056 800 110348 856
rect 110516 800 110808 856
rect 110976 800 111268 856
rect 111436 800 111728 856
rect 111896 800 112096 856
rect 112264 800 112556 856
rect 112724 800 113016 856
rect 113184 800 113476 856
rect 113644 800 113936 856
rect 114104 800 114396 856
rect 114564 800 114856 856
rect 115024 800 115316 856
rect 115484 800 115684 856
rect 115852 800 116144 856
rect 116312 800 116604 856
rect 116772 800 117064 856
rect 117232 800 117524 856
rect 117692 800 117984 856
rect 118152 800 118444 856
rect 118612 800 118904 856
rect 119072 800 119272 856
rect 119440 800 119732 856
rect 119900 800 120192 856
rect 120360 800 120652 856
rect 120820 800 121112 856
rect 121280 800 121572 856
rect 121740 800 122032 856
rect 122200 800 122492 856
rect 122660 800 122952 856
rect 123120 800 123320 856
rect 123488 800 123780 856
rect 123948 800 124240 856
rect 124408 800 124700 856
rect 124868 800 125160 856
rect 125328 800 125620 856
rect 125788 800 126080 856
rect 126248 800 126540 856
rect 126708 800 126908 856
rect 127076 800 127368 856
rect 127536 800 127828 856
rect 127996 800 128288 856
rect 128456 800 128748 856
rect 128916 800 129208 856
rect 129376 800 129668 856
rect 129836 800 130128 856
rect 130296 800 130496 856
rect 130664 800 130956 856
rect 131124 800 131416 856
rect 131584 800 131876 856
rect 132044 800 132336 856
rect 132504 800 132796 856
rect 132964 800 133256 856
rect 133424 800 133716 856
rect 133884 800 134084 856
rect 134252 800 134544 856
rect 134712 800 135004 856
rect 135172 800 135464 856
rect 135632 800 135924 856
rect 136092 800 136384 856
rect 136552 800 136844 856
rect 137012 800 137304 856
rect 137472 800 137764 856
rect 137932 800 138132 856
rect 138300 800 138592 856
rect 138760 800 139052 856
rect 139220 800 139512 856
rect 139680 800 139972 856
rect 140140 800 140432 856
rect 140600 800 140892 856
rect 141060 800 141352 856
rect 141520 800 141720 856
rect 141888 800 142180 856
rect 142348 800 142640 856
rect 142808 800 143100 856
rect 143268 800 143560 856
rect 143728 800 144020 856
rect 144188 800 144480 856
rect 144648 800 144940 856
rect 145108 800 145308 856
rect 145476 800 145768 856
rect 145936 800 146228 856
rect 146396 800 146688 856
rect 146856 800 147148 856
rect 147316 800 147608 856
rect 147776 800 148068 856
rect 148236 800 148528 856
rect 148696 800 148988 856
rect 149156 800 149356 856
rect 149524 800 149816 856
rect 149984 800 150276 856
rect 150444 800 150736 856
rect 150904 800 151196 856
rect 151364 800 151656 856
rect 151824 800 152116 856
rect 152284 800 152576 856
rect 152744 800 152944 856
rect 153112 800 153404 856
rect 153572 800 153864 856
rect 154032 800 154324 856
rect 154492 800 154784 856
rect 154952 800 155244 856
rect 155412 800 155704 856
rect 155872 800 156164 856
rect 156332 800 156532 856
rect 156700 800 156992 856
rect 157160 800 157452 856
rect 157620 800 157912 856
rect 158080 800 158372 856
rect 158540 800 158832 856
rect 159000 800 159292 856
rect 159460 800 159752 856
rect 159920 800 160212 856
rect 160380 800 160580 856
rect 160748 800 161040 856
rect 161208 800 161500 856
rect 161668 800 161960 856
rect 162128 800 162420 856
rect 162588 800 162880 856
rect 163048 800 163340 856
rect 163508 800 163800 856
rect 163968 800 164168 856
rect 164336 800 164628 856
rect 164796 800 165088 856
rect 165256 800 165548 856
rect 165716 800 166008 856
rect 166176 800 166468 856
rect 166636 800 166928 856
rect 167096 800 167388 856
rect 167556 800 167756 856
rect 167924 800 168216 856
rect 168384 800 168676 856
rect 168844 800 169136 856
rect 169304 800 169596 856
rect 169764 800 170056 856
rect 170224 800 170516 856
rect 170684 800 170976 856
rect 171144 800 171436 856
rect 171604 800 171804 856
rect 171972 800 172264 856
rect 172432 800 172724 856
rect 172892 800 173184 856
rect 173352 800 173644 856
rect 173812 800 174104 856
rect 174272 800 174564 856
rect 174732 800 175024 856
rect 175192 800 175392 856
rect 175560 800 175852 856
rect 176020 800 176312 856
rect 176480 800 176772 856
rect 176940 800 177232 856
rect 177400 800 177692 856
rect 177860 800 178152 856
rect 178320 800 178612 856
rect 178780 800 178980 856
rect 179148 800 179440 856
rect 179608 800 179900 856
rect 180068 800 180360 856
rect 180528 800 180820 856
rect 180988 800 181280 856
rect 181448 800 181740 856
rect 181908 800 182200 856
rect 182368 800 182568 856
rect 182736 800 183028 856
rect 183196 800 183488 856
rect 183656 800 183948 856
rect 184116 800 184408 856
rect 184576 800 184868 856
rect 185036 800 185328 856
rect 185496 800 185788 856
rect 185956 800 186248 856
rect 186416 800 186616 856
rect 186784 800 187076 856
rect 187244 800 187536 856
rect 187704 800 187996 856
rect 188164 800 188456 856
rect 188624 800 188916 856
rect 189084 800 189376 856
rect 189544 800 189836 856
rect 190004 800 190204 856
rect 190372 800 190664 856
rect 190832 800 191124 856
rect 191292 800 191584 856
rect 191752 800 192044 856
rect 192212 800 192504 856
rect 192672 800 192964 856
rect 193132 800 193424 856
rect 193592 800 193792 856
rect 193960 800 194252 856
rect 194420 800 194712 856
rect 194880 800 195172 856
rect 195340 800 195632 856
rect 195800 800 196092 856
rect 196260 800 196552 856
rect 196720 800 197012 856
rect 197180 800 197472 856
rect 197640 800 197840 856
rect 198008 800 198300 856
rect 198468 800 198760 856
rect 198928 800 199220 856
rect 199388 800 199680 856
rect 199848 800 200140 856
rect 200308 800 200600 856
rect 200768 800 201060 856
rect 201228 800 201428 856
rect 201596 800 201888 856
rect 202056 800 202348 856
rect 202516 800 202808 856
rect 202976 800 203268 856
rect 203436 800 203728 856
rect 203896 800 204188 856
rect 204356 800 204648 856
rect 204816 800 205016 856
rect 205184 800 205476 856
rect 205644 800 205936 856
rect 206104 800 206396 856
rect 206564 800 206856 856
rect 207024 800 207316 856
rect 207484 800 207776 856
rect 207944 800 208236 856
rect 208404 800 208696 856
rect 208864 800 209064 856
rect 209232 800 209524 856
rect 209692 800 209984 856
rect 210152 800 210444 856
rect 210612 800 210904 856
rect 211072 800 211364 856
rect 211532 800 211824 856
rect 211992 800 212284 856
rect 212452 800 212652 856
rect 212820 800 213112 856
rect 213280 800 213572 856
rect 213740 800 214032 856
rect 214200 800 214492 856
rect 214660 800 214952 856
rect 215120 800 215412 856
rect 215580 800 215872 856
rect 216040 800 216240 856
rect 216408 800 216700 856
rect 216868 800 217160 856
rect 217328 800 217620 856
rect 217788 800 218080 856
rect 218248 800 218540 856
rect 218708 800 219000 856
rect 219168 800 219460 856
<< obsm3 >>
rect 367 2143 217185 217633
<< metal4 >>
rect 4010 2128 4330 217648
rect 19370 2128 19690 217648
<< obsm4 >>
rect 13109 2128 19290 217648
rect 19770 2128 216495 217648
<< labels >>
rlabel metal2 s 740 219200 796 220000 6 io_in[0]
port 1 nsew default input
rlabel metal2 s 58608 219200 58664 220000 6 io_in[10]
port 2 nsew default input
rlabel metal2 s 64404 219200 64460 220000 6 io_in[11]
port 3 nsew default input
rlabel metal2 s 70200 219200 70256 220000 6 io_in[12]
port 4 nsew default input
rlabel metal2 s 75904 219200 75960 220000 6 io_in[13]
port 5 nsew default input
rlabel metal2 s 81700 219200 81756 220000 6 io_in[14]
port 6 nsew default input
rlabel metal2 s 87496 219200 87552 220000 6 io_in[15]
port 7 nsew default input
rlabel metal2 s 93292 219200 93348 220000 6 io_in[16]
port 8 nsew default input
rlabel metal2 s 99088 219200 99144 220000 6 io_in[17]
port 9 nsew default input
rlabel metal2 s 104884 219200 104940 220000 6 io_in[18]
port 10 nsew default input
rlabel metal2 s 110680 219200 110736 220000 6 io_in[19]
port 11 nsew default input
rlabel metal2 s 6444 219200 6500 220000 6 io_in[1]
port 12 nsew default input
rlabel metal2 s 116476 219200 116532 220000 6 io_in[20]
port 13 nsew default input
rlabel metal2 s 122272 219200 122328 220000 6 io_in[21]
port 14 nsew default input
rlabel metal2 s 128068 219200 128124 220000 6 io_in[22]
port 15 nsew default input
rlabel metal2 s 133864 219200 133920 220000 6 io_in[23]
port 16 nsew default input
rlabel metal2 s 139660 219200 139716 220000 6 io_in[24]
port 17 nsew default input
rlabel metal2 s 145456 219200 145512 220000 6 io_in[25]
port 18 nsew default input
rlabel metal2 s 151160 219200 151216 220000 6 io_in[26]
port 19 nsew default input
rlabel metal2 s 156956 219200 157012 220000 6 io_in[27]
port 20 nsew default input
rlabel metal2 s 162752 219200 162808 220000 6 io_in[28]
port 21 nsew default input
rlabel metal2 s 168548 219200 168604 220000 6 io_in[29]
port 22 nsew default input
rlabel metal2 s 12240 219200 12296 220000 6 io_in[2]
port 23 nsew default input
rlabel metal2 s 174344 219200 174400 220000 6 io_in[30]
port 24 nsew default input
rlabel metal2 s 180140 219200 180196 220000 6 io_in[31]
port 25 nsew default input
rlabel metal2 s 185936 219200 185992 220000 6 io_in[32]
port 26 nsew default input
rlabel metal2 s 191732 219200 191788 220000 6 io_in[33]
port 27 nsew default input
rlabel metal2 s 197528 219200 197584 220000 6 io_in[34]
port 28 nsew default input
rlabel metal2 s 203324 219200 203380 220000 6 io_in[35]
port 29 nsew default input
rlabel metal2 s 209120 219200 209176 220000 6 io_in[36]
port 30 nsew default input
rlabel metal2 s 214916 219200 214972 220000 6 io_in[37]
port 31 nsew default input
rlabel metal2 s 18036 219200 18092 220000 6 io_in[3]
port 32 nsew default input
rlabel metal2 s 23832 219200 23888 220000 6 io_in[4]
port 33 nsew default input
rlabel metal2 s 29628 219200 29684 220000 6 io_in[5]
port 34 nsew default input
rlabel metal2 s 35424 219200 35480 220000 6 io_in[6]
port 35 nsew default input
rlabel metal2 s 41220 219200 41276 220000 6 io_in[7]
port 36 nsew default input
rlabel metal2 s 47016 219200 47072 220000 6 io_in[8]
port 37 nsew default input
rlabel metal2 s 52812 219200 52868 220000 6 io_in[9]
port 38 nsew default input
rlabel metal2 s 2580 219200 2636 220000 6 io_oeb[0]
port 39 nsew default output
rlabel metal2 s 60540 219200 60596 220000 6 io_oeb[10]
port 40 nsew default output
rlabel metal2 s 66336 219200 66392 220000 6 io_oeb[11]
port 41 nsew default output
rlabel metal2 s 72132 219200 72188 220000 6 io_oeb[12]
port 42 nsew default output
rlabel metal2 s 77836 219200 77892 220000 6 io_oeb[13]
port 43 nsew default output
rlabel metal2 s 83632 219200 83688 220000 6 io_oeb[14]
port 44 nsew default output
rlabel metal2 s 89428 219200 89484 220000 6 io_oeb[15]
port 45 nsew default output
rlabel metal2 s 95224 219200 95280 220000 6 io_oeb[16]
port 46 nsew default output
rlabel metal2 s 101020 219200 101076 220000 6 io_oeb[17]
port 47 nsew default output
rlabel metal2 s 106816 219200 106872 220000 6 io_oeb[18]
port 48 nsew default output
rlabel metal2 s 112612 219200 112668 220000 6 io_oeb[19]
port 49 nsew default output
rlabel metal2 s 8376 219200 8432 220000 6 io_oeb[1]
port 50 nsew default output
rlabel metal2 s 118408 219200 118464 220000 6 io_oeb[20]
port 51 nsew default output
rlabel metal2 s 124204 219200 124260 220000 6 io_oeb[21]
port 52 nsew default output
rlabel metal2 s 130000 219200 130056 220000 6 io_oeb[22]
port 53 nsew default output
rlabel metal2 s 135796 219200 135852 220000 6 io_oeb[23]
port 54 nsew default output
rlabel metal2 s 141592 219200 141648 220000 6 io_oeb[24]
port 55 nsew default output
rlabel metal2 s 147388 219200 147444 220000 6 io_oeb[25]
port 56 nsew default output
rlabel metal2 s 153092 219200 153148 220000 6 io_oeb[26]
port 57 nsew default output
rlabel metal2 s 158888 219200 158944 220000 6 io_oeb[27]
port 58 nsew default output
rlabel metal2 s 164684 219200 164740 220000 6 io_oeb[28]
port 59 nsew default output
rlabel metal2 s 170480 219200 170536 220000 6 io_oeb[29]
port 60 nsew default output
rlabel metal2 s 14172 219200 14228 220000 6 io_oeb[2]
port 61 nsew default output
rlabel metal2 s 176276 219200 176332 220000 6 io_oeb[30]
port 62 nsew default output
rlabel metal2 s 182072 219200 182128 220000 6 io_oeb[31]
port 63 nsew default output
rlabel metal2 s 187868 219200 187924 220000 6 io_oeb[32]
port 64 nsew default output
rlabel metal2 s 193664 219200 193720 220000 6 io_oeb[33]
port 65 nsew default output
rlabel metal2 s 199460 219200 199516 220000 6 io_oeb[34]
port 66 nsew default output
rlabel metal2 s 205256 219200 205312 220000 6 io_oeb[35]
port 67 nsew default output
rlabel metal2 s 211052 219200 211108 220000 6 io_oeb[36]
port 68 nsew default output
rlabel metal2 s 216848 219200 216904 220000 6 io_oeb[37]
port 69 nsew default output
rlabel metal2 s 19968 219200 20024 220000 6 io_oeb[3]
port 70 nsew default output
rlabel metal2 s 25764 219200 25820 220000 6 io_oeb[4]
port 71 nsew default output
rlabel metal2 s 31560 219200 31616 220000 6 io_oeb[5]
port 72 nsew default output
rlabel metal2 s 37356 219200 37412 220000 6 io_oeb[6]
port 73 nsew default output
rlabel metal2 s 43152 219200 43208 220000 6 io_oeb[7]
port 74 nsew default output
rlabel metal2 s 48948 219200 49004 220000 6 io_oeb[8]
port 75 nsew default output
rlabel metal2 s 54744 219200 54800 220000 6 io_oeb[9]
port 76 nsew default output
rlabel metal2 s 4512 219200 4568 220000 6 io_out[0]
port 77 nsew default output
rlabel metal2 s 62472 219200 62528 220000 6 io_out[10]
port 78 nsew default output
rlabel metal2 s 68268 219200 68324 220000 6 io_out[11]
port 79 nsew default output
rlabel metal2 s 74064 219200 74120 220000 6 io_out[12]
port 80 nsew default output
rlabel metal2 s 79768 219200 79824 220000 6 io_out[13]
port 81 nsew default output
rlabel metal2 s 85564 219200 85620 220000 6 io_out[14]
port 82 nsew default output
rlabel metal2 s 91360 219200 91416 220000 6 io_out[15]
port 83 nsew default output
rlabel metal2 s 97156 219200 97212 220000 6 io_out[16]
port 84 nsew default output
rlabel metal2 s 102952 219200 103008 220000 6 io_out[17]
port 85 nsew default output
rlabel metal2 s 108748 219200 108804 220000 6 io_out[18]
port 86 nsew default output
rlabel metal2 s 114544 219200 114600 220000 6 io_out[19]
port 87 nsew default output
rlabel metal2 s 10308 219200 10364 220000 6 io_out[1]
port 88 nsew default output
rlabel metal2 s 120340 219200 120396 220000 6 io_out[20]
port 89 nsew default output
rlabel metal2 s 126136 219200 126192 220000 6 io_out[21]
port 90 nsew default output
rlabel metal2 s 131932 219200 131988 220000 6 io_out[22]
port 91 nsew default output
rlabel metal2 s 137728 219200 137784 220000 6 io_out[23]
port 92 nsew default output
rlabel metal2 s 143524 219200 143580 220000 6 io_out[24]
port 93 nsew default output
rlabel metal2 s 149228 219200 149284 220000 6 io_out[25]
port 94 nsew default output
rlabel metal2 s 155024 219200 155080 220000 6 io_out[26]
port 95 nsew default output
rlabel metal2 s 160820 219200 160876 220000 6 io_out[27]
port 96 nsew default output
rlabel metal2 s 166616 219200 166672 220000 6 io_out[28]
port 97 nsew default output
rlabel metal2 s 172412 219200 172468 220000 6 io_out[29]
port 98 nsew default output
rlabel metal2 s 16104 219200 16160 220000 6 io_out[2]
port 99 nsew default output
rlabel metal2 s 178208 219200 178264 220000 6 io_out[30]
port 100 nsew default output
rlabel metal2 s 184004 219200 184060 220000 6 io_out[31]
port 101 nsew default output
rlabel metal2 s 189800 219200 189856 220000 6 io_out[32]
port 102 nsew default output
rlabel metal2 s 195596 219200 195652 220000 6 io_out[33]
port 103 nsew default output
rlabel metal2 s 201392 219200 201448 220000 6 io_out[34]
port 104 nsew default output
rlabel metal2 s 207188 219200 207244 220000 6 io_out[35]
port 105 nsew default output
rlabel metal2 s 212984 219200 213040 220000 6 io_out[36]
port 106 nsew default output
rlabel metal2 s 218780 219200 218836 220000 6 io_out[37]
port 107 nsew default output
rlabel metal2 s 21900 219200 21956 220000 6 io_out[3]
port 108 nsew default output
rlabel metal2 s 27696 219200 27752 220000 6 io_out[4]
port 109 nsew default output
rlabel metal2 s 33492 219200 33548 220000 6 io_out[5]
port 110 nsew default output
rlabel metal2 s 39288 219200 39344 220000 6 io_out[6]
port 111 nsew default output
rlabel metal2 s 45084 219200 45140 220000 6 io_out[7]
port 112 nsew default output
rlabel metal2 s 50880 219200 50936 220000 6 io_out[8]
port 113 nsew default output
rlabel metal2 s 56676 219200 56732 220000 6 io_out[9]
port 114 nsew default output
rlabel metal2 s 47568 0 47624 800 6 la_data_in[0]
port 115 nsew default input
rlabel metal2 s 182256 0 182312 800 6 la_data_in[100]
port 116 nsew default input
rlabel metal2 s 183544 0 183600 800 6 la_data_in[101]
port 117 nsew default input
rlabel metal2 s 184924 0 184980 800 6 la_data_in[102]
port 118 nsew default input
rlabel metal2 s 186304 0 186360 800 6 la_data_in[103]
port 119 nsew default input
rlabel metal2 s 187592 0 187648 800 6 la_data_in[104]
port 120 nsew default input
rlabel metal2 s 188972 0 189028 800 6 la_data_in[105]
port 121 nsew default input
rlabel metal2 s 190260 0 190316 800 6 la_data_in[106]
port 122 nsew default input
rlabel metal2 s 191640 0 191696 800 6 la_data_in[107]
port 123 nsew default input
rlabel metal2 s 193020 0 193076 800 6 la_data_in[108]
port 124 nsew default input
rlabel metal2 s 194308 0 194364 800 6 la_data_in[109]
port 125 nsew default input
rlabel metal2 s 61000 0 61056 800 6 la_data_in[10]
port 126 nsew default input
rlabel metal2 s 195688 0 195744 800 6 la_data_in[110]
port 127 nsew default input
rlabel metal2 s 197068 0 197124 800 6 la_data_in[111]
port 128 nsew default input
rlabel metal2 s 198356 0 198412 800 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 199736 0 199792 800 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 201116 0 201172 800 6 la_data_in[114]
port 131 nsew default input
rlabel metal2 s 202404 0 202460 800 6 la_data_in[115]
port 132 nsew default input
rlabel metal2 s 203784 0 203840 800 6 la_data_in[116]
port 133 nsew default input
rlabel metal2 s 205072 0 205128 800 6 la_data_in[117]
port 134 nsew default input
rlabel metal2 s 206452 0 206508 800 6 la_data_in[118]
port 135 nsew default input
rlabel metal2 s 207832 0 207888 800 6 la_data_in[119]
port 136 nsew default input
rlabel metal2 s 62380 0 62436 800 6 la_data_in[11]
port 137 nsew default input
rlabel metal2 s 209120 0 209176 800 6 la_data_in[120]
port 138 nsew default input
rlabel metal2 s 210500 0 210556 800 6 la_data_in[121]
port 139 nsew default input
rlabel metal2 s 211880 0 211936 800 6 la_data_in[122]
port 140 nsew default input
rlabel metal2 s 213168 0 213224 800 6 la_data_in[123]
port 141 nsew default input
rlabel metal2 s 214548 0 214604 800 6 la_data_in[124]
port 142 nsew default input
rlabel metal2 s 215928 0 215984 800 6 la_data_in[125]
port 143 nsew default input
rlabel metal2 s 217216 0 217272 800 6 la_data_in[126]
port 144 nsew default input
rlabel metal2 s 218596 0 218652 800 6 la_data_in[127]
port 145 nsew default input
rlabel metal2 s 63668 0 63724 800 6 la_data_in[12]
port 146 nsew default input
rlabel metal2 s 65048 0 65104 800 6 la_data_in[13]
port 147 nsew default input
rlabel metal2 s 66428 0 66484 800 6 la_data_in[14]
port 148 nsew default input
rlabel metal2 s 67716 0 67772 800 6 la_data_in[15]
port 149 nsew default input
rlabel metal2 s 69096 0 69152 800 6 la_data_in[16]
port 150 nsew default input
rlabel metal2 s 70476 0 70532 800 6 la_data_in[17]
port 151 nsew default input
rlabel metal2 s 71764 0 71820 800 6 la_data_in[18]
port 152 nsew default input
rlabel metal2 s 73144 0 73200 800 6 la_data_in[19]
port 153 nsew default input
rlabel metal2 s 48856 0 48912 800 6 la_data_in[1]
port 154 nsew default input
rlabel metal2 s 74524 0 74580 800 6 la_data_in[20]
port 155 nsew default input
rlabel metal2 s 75812 0 75868 800 6 la_data_in[21]
port 156 nsew default input
rlabel metal2 s 77192 0 77248 800 6 la_data_in[22]
port 157 nsew default input
rlabel metal2 s 78480 0 78536 800 6 la_data_in[23]
port 158 nsew default input
rlabel metal2 s 79860 0 79916 800 6 la_data_in[24]
port 159 nsew default input
rlabel metal2 s 81240 0 81296 800 6 la_data_in[25]
port 160 nsew default input
rlabel metal2 s 82528 0 82584 800 6 la_data_in[26]
port 161 nsew default input
rlabel metal2 s 83908 0 83964 800 6 la_data_in[27]
port 162 nsew default input
rlabel metal2 s 85288 0 85344 800 6 la_data_in[28]
port 163 nsew default input
rlabel metal2 s 86576 0 86632 800 6 la_data_in[29]
port 164 nsew default input
rlabel metal2 s 50236 0 50292 800 6 la_data_in[2]
port 165 nsew default input
rlabel metal2 s 87956 0 88012 800 6 la_data_in[30]
port 166 nsew default input
rlabel metal2 s 89336 0 89392 800 6 la_data_in[31]
port 167 nsew default input
rlabel metal2 s 90624 0 90680 800 6 la_data_in[32]
port 168 nsew default input
rlabel metal2 s 92004 0 92060 800 6 la_data_in[33]
port 169 nsew default input
rlabel metal2 s 93292 0 93348 800 6 la_data_in[34]
port 170 nsew default input
rlabel metal2 s 94672 0 94728 800 6 la_data_in[35]
port 171 nsew default input
rlabel metal2 s 96052 0 96108 800 6 la_data_in[36]
port 172 nsew default input
rlabel metal2 s 97340 0 97396 800 6 la_data_in[37]
port 173 nsew default input
rlabel metal2 s 98720 0 98776 800 6 la_data_in[38]
port 174 nsew default input
rlabel metal2 s 100100 0 100156 800 6 la_data_in[39]
port 175 nsew default input
rlabel metal2 s 51616 0 51672 800 6 la_data_in[3]
port 176 nsew default input
rlabel metal2 s 101388 0 101444 800 6 la_data_in[40]
port 177 nsew default input
rlabel metal2 s 102768 0 102824 800 6 la_data_in[41]
port 178 nsew default input
rlabel metal2 s 104148 0 104204 800 6 la_data_in[42]
port 179 nsew default input
rlabel metal2 s 105436 0 105492 800 6 la_data_in[43]
port 180 nsew default input
rlabel metal2 s 106816 0 106872 800 6 la_data_in[44]
port 181 nsew default input
rlabel metal2 s 108104 0 108160 800 6 la_data_in[45]
port 182 nsew default input
rlabel metal2 s 109484 0 109540 800 6 la_data_in[46]
port 183 nsew default input
rlabel metal2 s 110864 0 110920 800 6 la_data_in[47]
port 184 nsew default input
rlabel metal2 s 112152 0 112208 800 6 la_data_in[48]
port 185 nsew default input
rlabel metal2 s 113532 0 113588 800 6 la_data_in[49]
port 186 nsew default input
rlabel metal2 s 52904 0 52960 800 6 la_data_in[4]
port 187 nsew default input
rlabel metal2 s 114912 0 114968 800 6 la_data_in[50]
port 188 nsew default input
rlabel metal2 s 116200 0 116256 800 6 la_data_in[51]
port 189 nsew default input
rlabel metal2 s 117580 0 117636 800 6 la_data_in[52]
port 190 nsew default input
rlabel metal2 s 118960 0 119016 800 6 la_data_in[53]
port 191 nsew default input
rlabel metal2 s 120248 0 120304 800 6 la_data_in[54]
port 192 nsew default input
rlabel metal2 s 121628 0 121684 800 6 la_data_in[55]
port 193 nsew default input
rlabel metal2 s 123008 0 123064 800 6 la_data_in[56]
port 194 nsew default input
rlabel metal2 s 124296 0 124352 800 6 la_data_in[57]
port 195 nsew default input
rlabel metal2 s 125676 0 125732 800 6 la_data_in[58]
port 196 nsew default input
rlabel metal2 s 126964 0 127020 800 6 la_data_in[59]
port 197 nsew default input
rlabel metal2 s 54284 0 54340 800 6 la_data_in[5]
port 198 nsew default input
rlabel metal2 s 128344 0 128400 800 6 la_data_in[60]
port 199 nsew default input
rlabel metal2 s 129724 0 129780 800 6 la_data_in[61]
port 200 nsew default input
rlabel metal2 s 131012 0 131068 800 6 la_data_in[62]
port 201 nsew default input
rlabel metal2 s 132392 0 132448 800 6 la_data_in[63]
port 202 nsew default input
rlabel metal2 s 133772 0 133828 800 6 la_data_in[64]
port 203 nsew default input
rlabel metal2 s 135060 0 135116 800 6 la_data_in[65]
port 204 nsew default input
rlabel metal2 s 136440 0 136496 800 6 la_data_in[66]
port 205 nsew default input
rlabel metal2 s 137820 0 137876 800 6 la_data_in[67]
port 206 nsew default input
rlabel metal2 s 139108 0 139164 800 6 la_data_in[68]
port 207 nsew default input
rlabel metal2 s 140488 0 140544 800 6 la_data_in[69]
port 208 nsew default input
rlabel metal2 s 55664 0 55720 800 6 la_data_in[6]
port 209 nsew default input
rlabel metal2 s 141776 0 141832 800 6 la_data_in[70]
port 210 nsew default input
rlabel metal2 s 143156 0 143212 800 6 la_data_in[71]
port 211 nsew default input
rlabel metal2 s 144536 0 144592 800 6 la_data_in[72]
port 212 nsew default input
rlabel metal2 s 145824 0 145880 800 6 la_data_in[73]
port 213 nsew default input
rlabel metal2 s 147204 0 147260 800 6 la_data_in[74]
port 214 nsew default input
rlabel metal2 s 148584 0 148640 800 6 la_data_in[75]
port 215 nsew default input
rlabel metal2 s 149872 0 149928 800 6 la_data_in[76]
port 216 nsew default input
rlabel metal2 s 151252 0 151308 800 6 la_data_in[77]
port 217 nsew default input
rlabel metal2 s 152632 0 152688 800 6 la_data_in[78]
port 218 nsew default input
rlabel metal2 s 153920 0 153976 800 6 la_data_in[79]
port 219 nsew default input
rlabel metal2 s 56952 0 57008 800 6 la_data_in[7]
port 220 nsew default input
rlabel metal2 s 155300 0 155356 800 6 la_data_in[80]
port 221 nsew default input
rlabel metal2 s 156588 0 156644 800 6 la_data_in[81]
port 222 nsew default input
rlabel metal2 s 157968 0 158024 800 6 la_data_in[82]
port 223 nsew default input
rlabel metal2 s 159348 0 159404 800 6 la_data_in[83]
port 224 nsew default input
rlabel metal2 s 160636 0 160692 800 6 la_data_in[84]
port 225 nsew default input
rlabel metal2 s 162016 0 162072 800 6 la_data_in[85]
port 226 nsew default input
rlabel metal2 s 163396 0 163452 800 6 la_data_in[86]
port 227 nsew default input
rlabel metal2 s 164684 0 164740 800 6 la_data_in[87]
port 228 nsew default input
rlabel metal2 s 166064 0 166120 800 6 la_data_in[88]
port 229 nsew default input
rlabel metal2 s 167444 0 167500 800 6 la_data_in[89]
port 230 nsew default input
rlabel metal2 s 58332 0 58388 800 6 la_data_in[8]
port 231 nsew default input
rlabel metal2 s 168732 0 168788 800 6 la_data_in[90]
port 232 nsew default input
rlabel metal2 s 170112 0 170168 800 6 la_data_in[91]
port 233 nsew default input
rlabel metal2 s 171492 0 171548 800 6 la_data_in[92]
port 234 nsew default input
rlabel metal2 s 172780 0 172836 800 6 la_data_in[93]
port 235 nsew default input
rlabel metal2 s 174160 0 174216 800 6 la_data_in[94]
port 236 nsew default input
rlabel metal2 s 175448 0 175504 800 6 la_data_in[95]
port 237 nsew default input
rlabel metal2 s 176828 0 176884 800 6 la_data_in[96]
port 238 nsew default input
rlabel metal2 s 178208 0 178264 800 6 la_data_in[97]
port 239 nsew default input
rlabel metal2 s 179496 0 179552 800 6 la_data_in[98]
port 240 nsew default input
rlabel metal2 s 180876 0 180932 800 6 la_data_in[99]
port 241 nsew default input
rlabel metal2 s 59620 0 59676 800 6 la_data_in[9]
port 242 nsew default input
rlabel metal2 s 48028 0 48084 800 6 la_data_out[0]
port 243 nsew default output
rlabel metal2 s 182624 0 182680 800 6 la_data_out[100]
port 244 nsew default output
rlabel metal2 s 184004 0 184060 800 6 la_data_out[101]
port 245 nsew default output
rlabel metal2 s 185384 0 185440 800 6 la_data_out[102]
port 246 nsew default output
rlabel metal2 s 186672 0 186728 800 6 la_data_out[103]
port 247 nsew default output
rlabel metal2 s 188052 0 188108 800 6 la_data_out[104]
port 248 nsew default output
rlabel metal2 s 189432 0 189488 800 6 la_data_out[105]
port 249 nsew default output
rlabel metal2 s 190720 0 190776 800 6 la_data_out[106]
port 250 nsew default output
rlabel metal2 s 192100 0 192156 800 6 la_data_out[107]
port 251 nsew default output
rlabel metal2 s 193480 0 193536 800 6 la_data_out[108]
port 252 nsew default output
rlabel metal2 s 194768 0 194824 800 6 la_data_out[109]
port 253 nsew default output
rlabel metal2 s 61460 0 61516 800 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 196148 0 196204 800 6 la_data_out[110]
port 255 nsew default output
rlabel metal2 s 197528 0 197584 800 6 la_data_out[111]
port 256 nsew default output
rlabel metal2 s 198816 0 198872 800 6 la_data_out[112]
port 257 nsew default output
rlabel metal2 s 200196 0 200252 800 6 la_data_out[113]
port 258 nsew default output
rlabel metal2 s 201484 0 201540 800 6 la_data_out[114]
port 259 nsew default output
rlabel metal2 s 202864 0 202920 800 6 la_data_out[115]
port 260 nsew default output
rlabel metal2 s 204244 0 204300 800 6 la_data_out[116]
port 261 nsew default output
rlabel metal2 s 205532 0 205588 800 6 la_data_out[117]
port 262 nsew default output
rlabel metal2 s 206912 0 206968 800 6 la_data_out[118]
port 263 nsew default output
rlabel metal2 s 208292 0 208348 800 6 la_data_out[119]
port 264 nsew default output
rlabel metal2 s 62840 0 62896 800 6 la_data_out[11]
port 265 nsew default output
rlabel metal2 s 209580 0 209636 800 6 la_data_out[120]
port 266 nsew default output
rlabel metal2 s 210960 0 211016 800 6 la_data_out[121]
port 267 nsew default output
rlabel metal2 s 212340 0 212396 800 6 la_data_out[122]
port 268 nsew default output
rlabel metal2 s 213628 0 213684 800 6 la_data_out[123]
port 269 nsew default output
rlabel metal2 s 215008 0 215064 800 6 la_data_out[124]
port 270 nsew default output
rlabel metal2 s 216296 0 216352 800 6 la_data_out[125]
port 271 nsew default output
rlabel metal2 s 217676 0 217732 800 6 la_data_out[126]
port 272 nsew default output
rlabel metal2 s 219056 0 219112 800 6 la_data_out[127]
port 273 nsew default output
rlabel metal2 s 64128 0 64184 800 6 la_data_out[12]
port 274 nsew default output
rlabel metal2 s 65508 0 65564 800 6 la_data_out[13]
port 275 nsew default output
rlabel metal2 s 66888 0 66944 800 6 la_data_out[14]
port 276 nsew default output
rlabel metal2 s 68176 0 68232 800 6 la_data_out[15]
port 277 nsew default output
rlabel metal2 s 69556 0 69612 800 6 la_data_out[16]
port 278 nsew default output
rlabel metal2 s 70844 0 70900 800 6 la_data_out[17]
port 279 nsew default output
rlabel metal2 s 72224 0 72280 800 6 la_data_out[18]
port 280 nsew default output
rlabel metal2 s 73604 0 73660 800 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 49316 0 49372 800 6 la_data_out[1]
port 282 nsew default output
rlabel metal2 s 74892 0 74948 800 6 la_data_out[20]
port 283 nsew default output
rlabel metal2 s 76272 0 76328 800 6 la_data_out[21]
port 284 nsew default output
rlabel metal2 s 77652 0 77708 800 6 la_data_out[22]
port 285 nsew default output
rlabel metal2 s 78940 0 78996 800 6 la_data_out[23]
port 286 nsew default output
rlabel metal2 s 80320 0 80376 800 6 la_data_out[24]
port 287 nsew default output
rlabel metal2 s 81700 0 81756 800 6 la_data_out[25]
port 288 nsew default output
rlabel metal2 s 82988 0 83044 800 6 la_data_out[26]
port 289 nsew default output
rlabel metal2 s 84368 0 84424 800 6 la_data_out[27]
port 290 nsew default output
rlabel metal2 s 85748 0 85804 800 6 la_data_out[28]
port 291 nsew default output
rlabel metal2 s 87036 0 87092 800 6 la_data_out[29]
port 292 nsew default output
rlabel metal2 s 50696 0 50752 800 6 la_data_out[2]
port 293 nsew default output
rlabel metal2 s 88416 0 88472 800 6 la_data_out[30]
port 294 nsew default output
rlabel metal2 s 89704 0 89760 800 6 la_data_out[31]
port 295 nsew default output
rlabel metal2 s 91084 0 91140 800 6 la_data_out[32]
port 296 nsew default output
rlabel metal2 s 92464 0 92520 800 6 la_data_out[33]
port 297 nsew default output
rlabel metal2 s 93752 0 93808 800 6 la_data_out[34]
port 298 nsew default output
rlabel metal2 s 95132 0 95188 800 6 la_data_out[35]
port 299 nsew default output
rlabel metal2 s 96512 0 96568 800 6 la_data_out[36]
port 300 nsew default output
rlabel metal2 s 97800 0 97856 800 6 la_data_out[37]
port 301 nsew default output
rlabel metal2 s 99180 0 99236 800 6 la_data_out[38]
port 302 nsew default output
rlabel metal2 s 100560 0 100616 800 6 la_data_out[39]
port 303 nsew default output
rlabel metal2 s 52076 0 52132 800 6 la_data_out[3]
port 304 nsew default output
rlabel metal2 s 101848 0 101904 800 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 103228 0 103284 800 6 la_data_out[41]
port 306 nsew default output
rlabel metal2 s 104516 0 104572 800 6 la_data_out[42]
port 307 nsew default output
rlabel metal2 s 105896 0 105952 800 6 la_data_out[43]
port 308 nsew default output
rlabel metal2 s 107276 0 107332 800 6 la_data_out[44]
port 309 nsew default output
rlabel metal2 s 108564 0 108620 800 6 la_data_out[45]
port 310 nsew default output
rlabel metal2 s 109944 0 110000 800 6 la_data_out[46]
port 311 nsew default output
rlabel metal2 s 111324 0 111380 800 6 la_data_out[47]
port 312 nsew default output
rlabel metal2 s 112612 0 112668 800 6 la_data_out[48]
port 313 nsew default output
rlabel metal2 s 113992 0 114048 800 6 la_data_out[49]
port 314 nsew default output
rlabel metal2 s 53364 0 53420 800 6 la_data_out[4]
port 315 nsew default output
rlabel metal2 s 115372 0 115428 800 6 la_data_out[50]
port 316 nsew default output
rlabel metal2 s 116660 0 116716 800 6 la_data_out[51]
port 317 nsew default output
rlabel metal2 s 118040 0 118096 800 6 la_data_out[52]
port 318 nsew default output
rlabel metal2 s 119328 0 119384 800 6 la_data_out[53]
port 319 nsew default output
rlabel metal2 s 120708 0 120764 800 6 la_data_out[54]
port 320 nsew default output
rlabel metal2 s 122088 0 122144 800 6 la_data_out[55]
port 321 nsew default output
rlabel metal2 s 123376 0 123432 800 6 la_data_out[56]
port 322 nsew default output
rlabel metal2 s 124756 0 124812 800 6 la_data_out[57]
port 323 nsew default output
rlabel metal2 s 126136 0 126192 800 6 la_data_out[58]
port 324 nsew default output
rlabel metal2 s 127424 0 127480 800 6 la_data_out[59]
port 325 nsew default output
rlabel metal2 s 54744 0 54800 800 6 la_data_out[5]
port 326 nsew default output
rlabel metal2 s 128804 0 128860 800 6 la_data_out[60]
port 327 nsew default output
rlabel metal2 s 130184 0 130240 800 6 la_data_out[61]
port 328 nsew default output
rlabel metal2 s 131472 0 131528 800 6 la_data_out[62]
port 329 nsew default output
rlabel metal2 s 132852 0 132908 800 6 la_data_out[63]
port 330 nsew default output
rlabel metal2 s 134140 0 134196 800 6 la_data_out[64]
port 331 nsew default output
rlabel metal2 s 135520 0 135576 800 6 la_data_out[65]
port 332 nsew default output
rlabel metal2 s 136900 0 136956 800 6 la_data_out[66]
port 333 nsew default output
rlabel metal2 s 138188 0 138244 800 6 la_data_out[67]
port 334 nsew default output
rlabel metal2 s 139568 0 139624 800 6 la_data_out[68]
port 335 nsew default output
rlabel metal2 s 140948 0 141004 800 6 la_data_out[69]
port 336 nsew default output
rlabel metal2 s 56032 0 56088 800 6 la_data_out[6]
port 337 nsew default output
rlabel metal2 s 142236 0 142292 800 6 la_data_out[70]
port 338 nsew default output
rlabel metal2 s 143616 0 143672 800 6 la_data_out[71]
port 339 nsew default output
rlabel metal2 s 144996 0 145052 800 6 la_data_out[72]
port 340 nsew default output
rlabel metal2 s 146284 0 146340 800 6 la_data_out[73]
port 341 nsew default output
rlabel metal2 s 147664 0 147720 800 6 la_data_out[74]
port 342 nsew default output
rlabel metal2 s 149044 0 149100 800 6 la_data_out[75]
port 343 nsew default output
rlabel metal2 s 150332 0 150388 800 6 la_data_out[76]
port 344 nsew default output
rlabel metal2 s 151712 0 151768 800 6 la_data_out[77]
port 345 nsew default output
rlabel metal2 s 153000 0 153056 800 6 la_data_out[78]
port 346 nsew default output
rlabel metal2 s 154380 0 154436 800 6 la_data_out[79]
port 347 nsew default output
rlabel metal2 s 57412 0 57468 800 6 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 155760 0 155816 800 6 la_data_out[80]
port 349 nsew default output
rlabel metal2 s 157048 0 157104 800 6 la_data_out[81]
port 350 nsew default output
rlabel metal2 s 158428 0 158484 800 6 la_data_out[82]
port 351 nsew default output
rlabel metal2 s 159808 0 159864 800 6 la_data_out[83]
port 352 nsew default output
rlabel metal2 s 161096 0 161152 800 6 la_data_out[84]
port 353 nsew default output
rlabel metal2 s 162476 0 162532 800 6 la_data_out[85]
port 354 nsew default output
rlabel metal2 s 163856 0 163912 800 6 la_data_out[86]
port 355 nsew default output
rlabel metal2 s 165144 0 165200 800 6 la_data_out[87]
port 356 nsew default output
rlabel metal2 s 166524 0 166580 800 6 la_data_out[88]
port 357 nsew default output
rlabel metal2 s 167812 0 167868 800 6 la_data_out[89]
port 358 nsew default output
rlabel metal2 s 58792 0 58848 800 6 la_data_out[8]
port 359 nsew default output
rlabel metal2 s 169192 0 169248 800 6 la_data_out[90]
port 360 nsew default output
rlabel metal2 s 170572 0 170628 800 6 la_data_out[91]
port 361 nsew default output
rlabel metal2 s 171860 0 171916 800 6 la_data_out[92]
port 362 nsew default output
rlabel metal2 s 173240 0 173296 800 6 la_data_out[93]
port 363 nsew default output
rlabel metal2 s 174620 0 174676 800 6 la_data_out[94]
port 364 nsew default output
rlabel metal2 s 175908 0 175964 800 6 la_data_out[95]
port 365 nsew default output
rlabel metal2 s 177288 0 177344 800 6 la_data_out[96]
port 366 nsew default output
rlabel metal2 s 178668 0 178724 800 6 la_data_out[97]
port 367 nsew default output
rlabel metal2 s 179956 0 180012 800 6 la_data_out[98]
port 368 nsew default output
rlabel metal2 s 181336 0 181392 800 6 la_data_out[99]
port 369 nsew default output
rlabel metal2 s 60080 0 60136 800 6 la_data_out[9]
port 370 nsew default output
rlabel metal2 s 48396 0 48452 800 6 la_oen[0]
port 371 nsew default input
rlabel metal2 s 183084 0 183140 800 6 la_oen[100]
port 372 nsew default input
rlabel metal2 s 184464 0 184520 800 6 la_oen[101]
port 373 nsew default input
rlabel metal2 s 185844 0 185900 800 6 la_oen[102]
port 374 nsew default input
rlabel metal2 s 187132 0 187188 800 6 la_oen[103]
port 375 nsew default input
rlabel metal2 s 188512 0 188568 800 6 la_oen[104]
port 376 nsew default input
rlabel metal2 s 189892 0 189948 800 6 la_oen[105]
port 377 nsew default input
rlabel metal2 s 191180 0 191236 800 6 la_oen[106]
port 378 nsew default input
rlabel metal2 s 192560 0 192616 800 6 la_oen[107]
port 379 nsew default input
rlabel metal2 s 193848 0 193904 800 6 la_oen[108]
port 380 nsew default input
rlabel metal2 s 195228 0 195284 800 6 la_oen[109]
port 381 nsew default input
rlabel metal2 s 61920 0 61976 800 6 la_oen[10]
port 382 nsew default input
rlabel metal2 s 196608 0 196664 800 6 la_oen[110]
port 383 nsew default input
rlabel metal2 s 197896 0 197952 800 6 la_oen[111]
port 384 nsew default input
rlabel metal2 s 199276 0 199332 800 6 la_oen[112]
port 385 nsew default input
rlabel metal2 s 200656 0 200712 800 6 la_oen[113]
port 386 nsew default input
rlabel metal2 s 201944 0 202000 800 6 la_oen[114]
port 387 nsew default input
rlabel metal2 s 203324 0 203380 800 6 la_oen[115]
port 388 nsew default input
rlabel metal2 s 204704 0 204760 800 6 la_oen[116]
port 389 nsew default input
rlabel metal2 s 205992 0 206048 800 6 la_oen[117]
port 390 nsew default input
rlabel metal2 s 207372 0 207428 800 6 la_oen[118]
port 391 nsew default input
rlabel metal2 s 208752 0 208808 800 6 la_oen[119]
port 392 nsew default input
rlabel metal2 s 63300 0 63356 800 6 la_oen[11]
port 393 nsew default input
rlabel metal2 s 210040 0 210096 800 6 la_oen[120]
port 394 nsew default input
rlabel metal2 s 211420 0 211476 800 6 la_oen[121]
port 395 nsew default input
rlabel metal2 s 212708 0 212764 800 6 la_oen[122]
port 396 nsew default input
rlabel metal2 s 214088 0 214144 800 6 la_oen[123]
port 397 nsew default input
rlabel metal2 s 215468 0 215524 800 6 la_oen[124]
port 398 nsew default input
rlabel metal2 s 216756 0 216812 800 6 la_oen[125]
port 399 nsew default input
rlabel metal2 s 218136 0 218192 800 6 la_oen[126]
port 400 nsew default input
rlabel metal2 s 219516 0 219572 800 6 la_oen[127]
port 401 nsew default input
rlabel metal2 s 64588 0 64644 800 6 la_oen[12]
port 402 nsew default input
rlabel metal2 s 65968 0 66024 800 6 la_oen[13]
port 403 nsew default input
rlabel metal2 s 67256 0 67312 800 6 la_oen[14]
port 404 nsew default input
rlabel metal2 s 68636 0 68692 800 6 la_oen[15]
port 405 nsew default input
rlabel metal2 s 70016 0 70072 800 6 la_oen[16]
port 406 nsew default input
rlabel metal2 s 71304 0 71360 800 6 la_oen[17]
port 407 nsew default input
rlabel metal2 s 72684 0 72740 800 6 la_oen[18]
port 408 nsew default input
rlabel metal2 s 74064 0 74120 800 6 la_oen[19]
port 409 nsew default input
rlabel metal2 s 49776 0 49832 800 6 la_oen[1]
port 410 nsew default input
rlabel metal2 s 75352 0 75408 800 6 la_oen[20]
port 411 nsew default input
rlabel metal2 s 76732 0 76788 800 6 la_oen[21]
port 412 nsew default input
rlabel metal2 s 78112 0 78168 800 6 la_oen[22]
port 413 nsew default input
rlabel metal2 s 79400 0 79456 800 6 la_oen[23]
port 414 nsew default input
rlabel metal2 s 80780 0 80836 800 6 la_oen[24]
port 415 nsew default input
rlabel metal2 s 82068 0 82124 800 6 la_oen[25]
port 416 nsew default input
rlabel metal2 s 83448 0 83504 800 6 la_oen[26]
port 417 nsew default input
rlabel metal2 s 84828 0 84884 800 6 la_oen[27]
port 418 nsew default input
rlabel metal2 s 86116 0 86172 800 6 la_oen[28]
port 419 nsew default input
rlabel metal2 s 87496 0 87552 800 6 la_oen[29]
port 420 nsew default input
rlabel metal2 s 51156 0 51212 800 6 la_oen[2]
port 421 nsew default input
rlabel metal2 s 88876 0 88932 800 6 la_oen[30]
port 422 nsew default input
rlabel metal2 s 90164 0 90220 800 6 la_oen[31]
port 423 nsew default input
rlabel metal2 s 91544 0 91600 800 6 la_oen[32]
port 424 nsew default input
rlabel metal2 s 92924 0 92980 800 6 la_oen[33]
port 425 nsew default input
rlabel metal2 s 94212 0 94268 800 6 la_oen[34]
port 426 nsew default input
rlabel metal2 s 95592 0 95648 800 6 la_oen[35]
port 427 nsew default input
rlabel metal2 s 96880 0 96936 800 6 la_oen[36]
port 428 nsew default input
rlabel metal2 s 98260 0 98316 800 6 la_oen[37]
port 429 nsew default input
rlabel metal2 s 99640 0 99696 800 6 la_oen[38]
port 430 nsew default input
rlabel metal2 s 100928 0 100984 800 6 la_oen[39]
port 431 nsew default input
rlabel metal2 s 52444 0 52500 800 6 la_oen[3]
port 432 nsew default input
rlabel metal2 s 102308 0 102364 800 6 la_oen[40]
port 433 nsew default input
rlabel metal2 s 103688 0 103744 800 6 la_oen[41]
port 434 nsew default input
rlabel metal2 s 104976 0 105032 800 6 la_oen[42]
port 435 nsew default input
rlabel metal2 s 106356 0 106412 800 6 la_oen[43]
port 436 nsew default input
rlabel metal2 s 107736 0 107792 800 6 la_oen[44]
port 437 nsew default input
rlabel metal2 s 109024 0 109080 800 6 la_oen[45]
port 438 nsew default input
rlabel metal2 s 110404 0 110460 800 6 la_oen[46]
port 439 nsew default input
rlabel metal2 s 111784 0 111840 800 6 la_oen[47]
port 440 nsew default input
rlabel metal2 s 113072 0 113128 800 6 la_oen[48]
port 441 nsew default input
rlabel metal2 s 114452 0 114508 800 6 la_oen[49]
port 442 nsew default input
rlabel metal2 s 53824 0 53880 800 6 la_oen[4]
port 443 nsew default input
rlabel metal2 s 115740 0 115796 800 6 la_oen[50]
port 444 nsew default input
rlabel metal2 s 117120 0 117176 800 6 la_oen[51]
port 445 nsew default input
rlabel metal2 s 118500 0 118556 800 6 la_oen[52]
port 446 nsew default input
rlabel metal2 s 119788 0 119844 800 6 la_oen[53]
port 447 nsew default input
rlabel metal2 s 121168 0 121224 800 6 la_oen[54]
port 448 nsew default input
rlabel metal2 s 122548 0 122604 800 6 la_oen[55]
port 449 nsew default input
rlabel metal2 s 123836 0 123892 800 6 la_oen[56]
port 450 nsew default input
rlabel metal2 s 125216 0 125272 800 6 la_oen[57]
port 451 nsew default input
rlabel metal2 s 126596 0 126652 800 6 la_oen[58]
port 452 nsew default input
rlabel metal2 s 127884 0 127940 800 6 la_oen[59]
port 453 nsew default input
rlabel metal2 s 55204 0 55260 800 6 la_oen[5]
port 454 nsew default input
rlabel metal2 s 129264 0 129320 800 6 la_oen[60]
port 455 nsew default input
rlabel metal2 s 130552 0 130608 800 6 la_oen[61]
port 456 nsew default input
rlabel metal2 s 131932 0 131988 800 6 la_oen[62]
port 457 nsew default input
rlabel metal2 s 133312 0 133368 800 6 la_oen[63]
port 458 nsew default input
rlabel metal2 s 134600 0 134656 800 6 la_oen[64]
port 459 nsew default input
rlabel metal2 s 135980 0 136036 800 6 la_oen[65]
port 460 nsew default input
rlabel metal2 s 137360 0 137416 800 6 la_oen[66]
port 461 nsew default input
rlabel metal2 s 138648 0 138704 800 6 la_oen[67]
port 462 nsew default input
rlabel metal2 s 140028 0 140084 800 6 la_oen[68]
port 463 nsew default input
rlabel metal2 s 141408 0 141464 800 6 la_oen[69]
port 464 nsew default input
rlabel metal2 s 56492 0 56548 800 6 la_oen[6]
port 465 nsew default input
rlabel metal2 s 142696 0 142752 800 6 la_oen[70]
port 466 nsew default input
rlabel metal2 s 144076 0 144132 800 6 la_oen[71]
port 467 nsew default input
rlabel metal2 s 145364 0 145420 800 6 la_oen[72]
port 468 nsew default input
rlabel metal2 s 146744 0 146800 800 6 la_oen[73]
port 469 nsew default input
rlabel metal2 s 148124 0 148180 800 6 la_oen[74]
port 470 nsew default input
rlabel metal2 s 149412 0 149468 800 6 la_oen[75]
port 471 nsew default input
rlabel metal2 s 150792 0 150848 800 6 la_oen[76]
port 472 nsew default input
rlabel metal2 s 152172 0 152228 800 6 la_oen[77]
port 473 nsew default input
rlabel metal2 s 153460 0 153516 800 6 la_oen[78]
port 474 nsew default input
rlabel metal2 s 154840 0 154896 800 6 la_oen[79]
port 475 nsew default input
rlabel metal2 s 57872 0 57928 800 6 la_oen[7]
port 476 nsew default input
rlabel metal2 s 156220 0 156276 800 6 la_oen[80]
port 477 nsew default input
rlabel metal2 s 157508 0 157564 800 6 la_oen[81]
port 478 nsew default input
rlabel metal2 s 158888 0 158944 800 6 la_oen[82]
port 479 nsew default input
rlabel metal2 s 160268 0 160324 800 6 la_oen[83]
port 480 nsew default input
rlabel metal2 s 161556 0 161612 800 6 la_oen[84]
port 481 nsew default input
rlabel metal2 s 162936 0 162992 800 6 la_oen[85]
port 482 nsew default input
rlabel metal2 s 164224 0 164280 800 6 la_oen[86]
port 483 nsew default input
rlabel metal2 s 165604 0 165660 800 6 la_oen[87]
port 484 nsew default input
rlabel metal2 s 166984 0 167040 800 6 la_oen[88]
port 485 nsew default input
rlabel metal2 s 168272 0 168328 800 6 la_oen[89]
port 486 nsew default input
rlabel metal2 s 59252 0 59308 800 6 la_oen[8]
port 487 nsew default input
rlabel metal2 s 169652 0 169708 800 6 la_oen[90]
port 488 nsew default input
rlabel metal2 s 171032 0 171088 800 6 la_oen[91]
port 489 nsew default input
rlabel metal2 s 172320 0 172376 800 6 la_oen[92]
port 490 nsew default input
rlabel metal2 s 173700 0 173756 800 6 la_oen[93]
port 491 nsew default input
rlabel metal2 s 175080 0 175136 800 6 la_oen[94]
port 492 nsew default input
rlabel metal2 s 176368 0 176424 800 6 la_oen[95]
port 493 nsew default input
rlabel metal2 s 177748 0 177804 800 6 la_oen[96]
port 494 nsew default input
rlabel metal2 s 179036 0 179092 800 6 la_oen[97]
port 495 nsew default input
rlabel metal2 s 180416 0 180472 800 6 la_oen[98]
port 496 nsew default input
rlabel metal2 s 181796 0 181852 800 6 la_oen[99]
port 497 nsew default input
rlabel metal2 s 60540 0 60596 800 6 la_oen[9]
port 498 nsew default input
rlabel metal2 s 4 0 60 800 6 wb_clk_i
port 499 nsew default input
rlabel metal2 s 372 0 428 800 6 wb_rst_i
port 500 nsew default input
rlabel metal2 s 832 0 888 800 6 wbs_ack_o
port 501 nsew default output
rlabel metal2 s 2672 0 2728 800 6 wbs_adr_i[0]
port 502 nsew default input
rlabel metal2 s 17944 0 18000 800 6 wbs_adr_i[10]
port 503 nsew default input
rlabel metal2 s 19232 0 19288 800 6 wbs_adr_i[11]
port 504 nsew default input
rlabel metal2 s 20612 0 20668 800 6 wbs_adr_i[12]
port 505 nsew default input
rlabel metal2 s 21992 0 22048 800 6 wbs_adr_i[13]
port 506 nsew default input
rlabel metal2 s 23280 0 23336 800 6 wbs_adr_i[14]
port 507 nsew default input
rlabel metal2 s 24660 0 24716 800 6 wbs_adr_i[15]
port 508 nsew default input
rlabel metal2 s 26040 0 26096 800 6 wbs_adr_i[16]
port 509 nsew default input
rlabel metal2 s 27328 0 27384 800 6 wbs_adr_i[17]
port 510 nsew default input
rlabel metal2 s 28708 0 28764 800 6 wbs_adr_i[18]
port 511 nsew default input
rlabel metal2 s 29996 0 30052 800 6 wbs_adr_i[19]
port 512 nsew default input
rlabel metal2 s 4420 0 4476 800 6 wbs_adr_i[1]
port 513 nsew default input
rlabel metal2 s 31376 0 31432 800 6 wbs_adr_i[20]
port 514 nsew default input
rlabel metal2 s 32756 0 32812 800 6 wbs_adr_i[21]
port 515 nsew default input
rlabel metal2 s 34044 0 34100 800 6 wbs_adr_i[22]
port 516 nsew default input
rlabel metal2 s 35424 0 35480 800 6 wbs_adr_i[23]
port 517 nsew default input
rlabel metal2 s 36804 0 36860 800 6 wbs_adr_i[24]
port 518 nsew default input
rlabel metal2 s 38092 0 38148 800 6 wbs_adr_i[25]
port 519 nsew default input
rlabel metal2 s 39472 0 39528 800 6 wbs_adr_i[26]
port 520 nsew default input
rlabel metal2 s 40852 0 40908 800 6 wbs_adr_i[27]
port 521 nsew default input
rlabel metal2 s 42140 0 42196 800 6 wbs_adr_i[28]
port 522 nsew default input
rlabel metal2 s 43520 0 43576 800 6 wbs_adr_i[29]
port 523 nsew default input
rlabel metal2 s 6260 0 6316 800 6 wbs_adr_i[2]
port 524 nsew default input
rlabel metal2 s 44808 0 44864 800 6 wbs_adr_i[30]
port 525 nsew default input
rlabel metal2 s 46188 0 46244 800 6 wbs_adr_i[31]
port 526 nsew default input
rlabel metal2 s 8008 0 8064 800 6 wbs_adr_i[3]
port 527 nsew default input
rlabel metal2 s 9848 0 9904 800 6 wbs_adr_i[4]
port 528 nsew default input
rlabel metal2 s 11136 0 11192 800 6 wbs_adr_i[5]
port 529 nsew default input
rlabel metal2 s 12516 0 12572 800 6 wbs_adr_i[6]
port 530 nsew default input
rlabel metal2 s 13896 0 13952 800 6 wbs_adr_i[7]
port 531 nsew default input
rlabel metal2 s 15184 0 15240 800 6 wbs_adr_i[8]
port 532 nsew default input
rlabel metal2 s 16564 0 16620 800 6 wbs_adr_i[9]
port 533 nsew default input
rlabel metal2 s 1292 0 1348 800 6 wbs_cyc_i
port 534 nsew default input
rlabel metal2 s 3132 0 3188 800 6 wbs_dat_i[0]
port 535 nsew default input
rlabel metal2 s 18404 0 18460 800 6 wbs_dat_i[10]
port 536 nsew default input
rlabel metal2 s 19692 0 19748 800 6 wbs_dat_i[11]
port 537 nsew default input
rlabel metal2 s 21072 0 21128 800 6 wbs_dat_i[12]
port 538 nsew default input
rlabel metal2 s 22360 0 22416 800 6 wbs_dat_i[13]
port 539 nsew default input
rlabel metal2 s 23740 0 23796 800 6 wbs_dat_i[14]
port 540 nsew default input
rlabel metal2 s 25120 0 25176 800 6 wbs_dat_i[15]
port 541 nsew default input
rlabel metal2 s 26408 0 26464 800 6 wbs_dat_i[16]
port 542 nsew default input
rlabel metal2 s 27788 0 27844 800 6 wbs_dat_i[17]
port 543 nsew default input
rlabel metal2 s 29168 0 29224 800 6 wbs_dat_i[18]
port 544 nsew default input
rlabel metal2 s 30456 0 30512 800 6 wbs_dat_i[19]
port 545 nsew default input
rlabel metal2 s 4880 0 4936 800 6 wbs_dat_i[1]
port 546 nsew default input
rlabel metal2 s 31836 0 31892 800 6 wbs_dat_i[20]
port 547 nsew default input
rlabel metal2 s 33216 0 33272 800 6 wbs_dat_i[21]
port 548 nsew default input
rlabel metal2 s 34504 0 34560 800 6 wbs_dat_i[22]
port 549 nsew default input
rlabel metal2 s 35884 0 35940 800 6 wbs_dat_i[23]
port 550 nsew default input
rlabel metal2 s 37264 0 37320 800 6 wbs_dat_i[24]
port 551 nsew default input
rlabel metal2 s 38552 0 38608 800 6 wbs_dat_i[25]
port 552 nsew default input
rlabel metal2 s 39932 0 39988 800 6 wbs_dat_i[26]
port 553 nsew default input
rlabel metal2 s 41220 0 41276 800 6 wbs_dat_i[27]
port 554 nsew default input
rlabel metal2 s 42600 0 42656 800 6 wbs_dat_i[28]
port 555 nsew default input
rlabel metal2 s 43980 0 44036 800 6 wbs_dat_i[29]
port 556 nsew default input
rlabel metal2 s 6720 0 6776 800 6 wbs_dat_i[2]
port 557 nsew default input
rlabel metal2 s 45268 0 45324 800 6 wbs_dat_i[30]
port 558 nsew default input
rlabel metal2 s 46648 0 46704 800 6 wbs_dat_i[31]
port 559 nsew default input
rlabel metal2 s 8468 0 8524 800 6 wbs_dat_i[3]
port 560 nsew default input
rlabel metal2 s 10308 0 10364 800 6 wbs_dat_i[4]
port 561 nsew default input
rlabel metal2 s 11596 0 11652 800 6 wbs_dat_i[5]
port 562 nsew default input
rlabel metal2 s 12976 0 13032 800 6 wbs_dat_i[6]
port 563 nsew default input
rlabel metal2 s 14356 0 14412 800 6 wbs_dat_i[7]
port 564 nsew default input
rlabel metal2 s 15644 0 15700 800 6 wbs_dat_i[8]
port 565 nsew default input
rlabel metal2 s 17024 0 17080 800 6 wbs_dat_i[9]
port 566 nsew default input
rlabel metal2 s 3592 0 3648 800 6 wbs_dat_o[0]
port 567 nsew default output
rlabel metal2 s 18772 0 18828 800 6 wbs_dat_o[10]
port 568 nsew default output
rlabel metal2 s 20152 0 20208 800 6 wbs_dat_o[11]
port 569 nsew default output
rlabel metal2 s 21532 0 21588 800 6 wbs_dat_o[12]
port 570 nsew default output
rlabel metal2 s 22820 0 22876 800 6 wbs_dat_o[13]
port 571 nsew default output
rlabel metal2 s 24200 0 24256 800 6 wbs_dat_o[14]
port 572 nsew default output
rlabel metal2 s 25580 0 25636 800 6 wbs_dat_o[15]
port 573 nsew default output
rlabel metal2 s 26868 0 26924 800 6 wbs_dat_o[16]
port 574 nsew default output
rlabel metal2 s 28248 0 28304 800 6 wbs_dat_o[17]
port 575 nsew default output
rlabel metal2 s 29628 0 29684 800 6 wbs_dat_o[18]
port 576 nsew default output
rlabel metal2 s 30916 0 30972 800 6 wbs_dat_o[19]
port 577 nsew default output
rlabel metal2 s 5340 0 5396 800 6 wbs_dat_o[1]
port 578 nsew default output
rlabel metal2 s 32296 0 32352 800 6 wbs_dat_o[20]
port 579 nsew default output
rlabel metal2 s 33584 0 33640 800 6 wbs_dat_o[21]
port 580 nsew default output
rlabel metal2 s 34964 0 35020 800 6 wbs_dat_o[22]
port 581 nsew default output
rlabel metal2 s 36344 0 36400 800 6 wbs_dat_o[23]
port 582 nsew default output
rlabel metal2 s 37632 0 37688 800 6 wbs_dat_o[24]
port 583 nsew default output
rlabel metal2 s 39012 0 39068 800 6 wbs_dat_o[25]
port 584 nsew default output
rlabel metal2 s 40392 0 40448 800 6 wbs_dat_o[26]
port 585 nsew default output
rlabel metal2 s 41680 0 41736 800 6 wbs_dat_o[27]
port 586 nsew default output
rlabel metal2 s 43060 0 43116 800 6 wbs_dat_o[28]
port 587 nsew default output
rlabel metal2 s 44440 0 44496 800 6 wbs_dat_o[29]
port 588 nsew default output
rlabel metal2 s 7180 0 7236 800 6 wbs_dat_o[2]
port 589 nsew default output
rlabel metal2 s 45728 0 45784 800 6 wbs_dat_o[30]
port 590 nsew default output
rlabel metal2 s 47108 0 47164 800 6 wbs_dat_o[31]
port 591 nsew default output
rlabel metal2 s 8928 0 8984 800 6 wbs_dat_o[3]
port 592 nsew default output
rlabel metal2 s 10768 0 10824 800 6 wbs_dat_o[4]
port 593 nsew default output
rlabel metal2 s 12056 0 12112 800 6 wbs_dat_o[5]
port 594 nsew default output
rlabel metal2 s 13436 0 13492 800 6 wbs_dat_o[6]
port 595 nsew default output
rlabel metal2 s 14816 0 14872 800 6 wbs_dat_o[7]
port 596 nsew default output
rlabel metal2 s 16104 0 16160 800 6 wbs_dat_o[8]
port 597 nsew default output
rlabel metal2 s 17484 0 17540 800 6 wbs_dat_o[9]
port 598 nsew default output
rlabel metal2 s 3960 0 4016 800 6 wbs_sel_i[0]
port 599 nsew default input
rlabel metal2 s 5800 0 5856 800 6 wbs_sel_i[1]
port 600 nsew default input
rlabel metal2 s 7548 0 7604 800 6 wbs_sel_i[2]
port 601 nsew default input
rlabel metal2 s 9388 0 9444 800 6 wbs_sel_i[3]
port 602 nsew default input
rlabel metal2 s 1752 0 1808 800 6 wbs_stb_i
port 603 nsew default input
rlabel metal2 s 2212 0 2268 800 6 wbs_we_i
port 604 nsew default input
rlabel metal4 s 4010 2128 4330 217648 6 VPWR
port 605 nsew power input
rlabel metal4 s 19370 2128 19690 217648 6 VGND
port 606 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 219576 220000
string LEFview TRUE
<< end >>
