VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1393.870 84.560 1394.190 84.620 ;
        RECT 1441.710 84.560 1442.030 84.620 ;
        RECT 1393.870 84.420 1442.030 84.560 ;
        RECT 1393.870 84.360 1394.190 84.420 ;
        RECT 1441.710 84.360 1442.030 84.420 ;
        RECT 2042.010 84.220 2042.330 84.280 ;
        RECT 2053.510 84.220 2053.830 84.280 ;
        RECT 2042.010 84.080 2053.830 84.220 ;
        RECT 2042.010 84.020 2042.330 84.080 ;
        RECT 2053.510 84.020 2053.830 84.080 ;
        RECT 2379.650 84.220 2379.970 84.280 ;
        RECT 2387.470 84.220 2387.790 84.280 ;
        RECT 2379.650 84.080 2387.790 84.220 ;
        RECT 2379.650 84.020 2379.970 84.080 ;
        RECT 2387.470 84.020 2387.790 84.080 ;
        RECT 1738.410 83.540 1738.730 83.600 ;
        RECT 1779.810 83.540 1780.130 83.600 ;
        RECT 1738.410 83.400 1780.130 83.540 ;
        RECT 1738.410 83.340 1738.730 83.400 ;
        RECT 1779.810 83.340 1780.130 83.400 ;
        RECT 2608.270 83.540 2608.590 83.600 ;
        RECT 2622.530 83.540 2622.850 83.600 ;
        RECT 2608.270 83.400 2622.850 83.540 ;
        RECT 2608.270 83.340 2608.590 83.400 ;
        RECT 2622.530 83.340 2622.850 83.400 ;
      LAYER via ;
        RECT 1393.900 84.360 1394.160 84.620 ;
        RECT 1441.740 84.360 1442.000 84.620 ;
        RECT 2042.040 84.020 2042.300 84.280 ;
        RECT 2053.540 84.020 2053.800 84.280 ;
        RECT 2379.680 84.020 2379.940 84.280 ;
        RECT 2387.500 84.020 2387.760 84.280 ;
        RECT 1738.440 83.340 1738.700 83.600 ;
        RECT 1779.840 83.340 1780.100 83.600 ;
        RECT 2608.300 83.340 2608.560 83.600 ;
        RECT 2622.560 83.340 2622.820 83.600 ;
      LAYER met2 ;
        RECT 1155.080 3199.810 1155.360 3200.000 ;
        RECT 1156.990 3199.810 1157.270 3199.925 ;
        RECT 1155.080 3199.670 1157.270 3199.810 ;
        RECT 1155.080 3197.600 1155.360 3199.670 ;
        RECT 1156.990 3199.555 1157.270 3199.670 ;
        RECT 2801.030 86.515 2801.310 86.885 ;
        RECT 1345.130 85.835 1345.410 86.205 ;
        RECT 1676.330 85.835 1676.610 86.205 ;
        RECT 2704.430 85.835 2704.710 86.205 ;
        RECT 1345.200 84.165 1345.340 85.835 ;
        RECT 1393.890 84.475 1394.170 84.845 ;
        RECT 1617.910 84.730 1618.190 84.845 ;
        RECT 1393.900 84.330 1394.160 84.475 ;
        RECT 1441.740 84.330 1442.000 84.650 ;
        RECT 1617.520 84.590 1618.190 84.730 ;
        RECT 1220.930 84.050 1221.210 84.165 ;
        RECT 1221.850 84.050 1222.130 84.165 ;
        RECT 1220.930 83.910 1222.130 84.050 ;
        RECT 1220.930 83.795 1221.210 83.910 ;
        RECT 1221.850 83.795 1222.130 83.910 ;
        RECT 1345.130 83.795 1345.410 84.165 ;
        RECT 1441.800 83.485 1441.940 84.330 ;
        RECT 1617.520 84.165 1617.660 84.590 ;
        RECT 1617.910 84.475 1618.190 84.590 ;
        RECT 1676.400 84.165 1676.540 85.835 ;
        RECT 2053.530 85.155 2053.810 85.525 ;
        RECT 2090.330 85.155 2090.610 85.525 ;
        RECT 1779.830 84.475 1780.110 84.845 ;
        RECT 1545.230 83.795 1545.510 84.165 ;
        RECT 1617.450 83.795 1617.730 84.165 ;
        RECT 1676.330 83.795 1676.610 84.165 ;
        RECT 1441.730 83.115 1442.010 83.485 ;
        RECT 1496.470 83.115 1496.750 83.485 ;
        RECT 1496.540 82.805 1496.680 83.115 ;
        RECT 1496.470 82.435 1496.750 82.805 ;
        RECT 1545.300 82.125 1545.440 83.795 ;
        RECT 1779.900 83.630 1780.040 84.475 ;
        RECT 2053.600 84.310 2053.740 85.155 ;
        RECT 2090.400 84.730 2090.540 85.155 ;
        RECT 2091.250 84.730 2091.530 84.845 ;
        RECT 2090.400 84.590 2091.530 84.730 ;
        RECT 2091.250 84.475 2091.530 84.590 ;
        RECT 2283.990 84.475 2284.270 84.845 ;
        RECT 2622.550 84.475 2622.830 84.845 ;
        RECT 2042.040 84.165 2042.300 84.310 ;
        RECT 1852.510 83.795 1852.790 84.165 ;
        RECT 1932.550 83.795 1932.830 84.165 ;
        RECT 1994.650 83.795 1994.930 84.165 ;
        RECT 2042.030 83.795 2042.310 84.165 ;
        RECT 2053.540 83.990 2053.800 84.310 ;
        RECT 2283.530 84.050 2283.810 84.165 ;
        RECT 2284.060 84.050 2284.200 84.475 ;
        RECT 2379.680 84.165 2379.940 84.310 ;
        RECT 2387.500 84.165 2387.760 84.310 ;
        RECT 2283.530 83.910 2284.200 84.050 ;
        RECT 2283.530 83.795 2283.810 83.910 ;
        RECT 2379.670 83.795 2379.950 84.165 ;
        RECT 2387.490 83.795 2387.770 84.165 ;
        RECT 2572.870 83.795 2573.150 84.165 ;
        RECT 1738.440 83.485 1738.700 83.630 ;
        RECT 1731.070 83.115 1731.350 83.485 ;
        RECT 1738.430 83.115 1738.710 83.485 ;
        RECT 1779.840 83.310 1780.100 83.630 ;
        RECT 1731.140 82.805 1731.280 83.115 ;
        RECT 1731.070 82.435 1731.350 82.805 ;
        RECT 1852.580 82.125 1852.720 83.795 ;
        RECT 1932.620 82.805 1932.760 83.795 ;
        RECT 1994.720 82.805 1994.860 83.795 ;
        RECT 1932.550 82.435 1932.830 82.805 ;
        RECT 1994.650 82.435 1994.930 82.805 ;
        RECT 2572.940 82.125 2573.080 83.795 ;
        RECT 2622.620 83.630 2622.760 84.475 ;
        RECT 2704.500 84.165 2704.640 85.835 ;
        RECT 2801.100 84.845 2801.240 86.515 ;
        RECT 2801.030 84.475 2801.310 84.845 ;
        RECT 2704.430 83.795 2704.710 84.165 ;
        RECT 2863.130 83.795 2863.410 84.165 ;
        RECT 2608.300 83.485 2608.560 83.630 ;
        RECT 2608.290 83.115 2608.570 83.485 ;
        RECT 2622.560 83.310 2622.820 83.630 ;
        RECT 2863.200 83.370 2863.340 83.795 ;
        RECT 2863.590 83.370 2863.870 83.485 ;
        RECT 2863.200 83.230 2863.870 83.370 ;
        RECT 2863.590 83.115 2863.870 83.230 ;
        RECT 1545.230 81.755 1545.510 82.125 ;
        RECT 1852.510 81.755 1852.790 82.125 ;
        RECT 2572.870 81.755 2573.150 82.125 ;
      LAYER via2 ;
        RECT 1156.990 3199.600 1157.270 3199.880 ;
        RECT 2801.030 86.560 2801.310 86.840 ;
        RECT 1345.130 85.880 1345.410 86.160 ;
        RECT 1676.330 85.880 1676.610 86.160 ;
        RECT 2704.430 85.880 2704.710 86.160 ;
        RECT 1393.890 84.520 1394.170 84.800 ;
        RECT 1220.930 83.840 1221.210 84.120 ;
        RECT 1221.850 83.840 1222.130 84.120 ;
        RECT 1345.130 83.840 1345.410 84.120 ;
        RECT 1617.910 84.520 1618.190 84.800 ;
        RECT 2053.530 85.200 2053.810 85.480 ;
        RECT 2090.330 85.200 2090.610 85.480 ;
        RECT 1779.830 84.520 1780.110 84.800 ;
        RECT 1545.230 83.840 1545.510 84.120 ;
        RECT 1617.450 83.840 1617.730 84.120 ;
        RECT 1676.330 83.840 1676.610 84.120 ;
        RECT 1441.730 83.160 1442.010 83.440 ;
        RECT 1496.470 83.160 1496.750 83.440 ;
        RECT 1496.470 82.480 1496.750 82.760 ;
        RECT 2091.250 84.520 2091.530 84.800 ;
        RECT 2283.990 84.520 2284.270 84.800 ;
        RECT 2622.550 84.520 2622.830 84.800 ;
        RECT 1852.510 83.840 1852.790 84.120 ;
        RECT 1932.550 83.840 1932.830 84.120 ;
        RECT 1994.650 83.840 1994.930 84.120 ;
        RECT 2042.030 83.840 2042.310 84.120 ;
        RECT 2283.530 83.840 2283.810 84.120 ;
        RECT 2379.670 83.840 2379.950 84.120 ;
        RECT 2387.490 83.840 2387.770 84.120 ;
        RECT 2572.870 83.840 2573.150 84.120 ;
        RECT 1731.070 83.160 1731.350 83.440 ;
        RECT 1738.430 83.160 1738.710 83.440 ;
        RECT 1731.070 82.480 1731.350 82.760 ;
        RECT 1932.550 82.480 1932.830 82.760 ;
        RECT 1994.650 82.480 1994.930 82.760 ;
        RECT 2801.030 84.520 2801.310 84.800 ;
        RECT 2704.430 83.840 2704.710 84.120 ;
        RECT 2863.130 83.840 2863.410 84.120 ;
        RECT 2608.290 83.160 2608.570 83.440 ;
        RECT 2863.590 83.160 2863.870 83.440 ;
        RECT 1545.230 81.800 1545.510 82.080 ;
        RECT 1852.510 81.800 1852.790 82.080 ;
        RECT 2572.870 81.800 2573.150 82.080 ;
      LAYER met3 ;
        RECT 1156.965 3199.890 1157.295 3199.905 ;
        RECT 1158.550 3199.890 1158.930 3199.900 ;
        RECT 1156.965 3199.590 1158.930 3199.890 ;
        RECT 1156.965 3199.575 1157.295 3199.590 ;
        RECT 1158.550 3199.580 1158.930 3199.590 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2916.710 87.910 2924.800 88.210 ;
        RECT 2752.910 86.850 2753.290 86.860 ;
        RECT 2801.005 86.850 2801.335 86.865 ;
        RECT 2752.910 86.550 2801.335 86.850 ;
        RECT 2752.910 86.540 2753.290 86.550 ;
        RECT 2801.005 86.535 2801.335 86.550 ;
        RECT 1297.470 86.170 1297.850 86.180 ;
        RECT 1345.105 86.170 1345.435 86.185 ;
        RECT 1297.470 85.870 1345.435 86.170 ;
        RECT 1297.470 85.860 1297.850 85.870 ;
        RECT 1345.105 85.855 1345.435 85.870 ;
        RECT 1628.670 86.170 1629.050 86.180 ;
        RECT 1676.305 86.170 1676.635 86.185 ;
        RECT 1628.670 85.870 1676.635 86.170 ;
        RECT 1628.670 85.860 1629.050 85.870 ;
        RECT 1676.305 85.855 1676.635 85.870 ;
        RECT 2656.310 86.170 2656.690 86.180 ;
        RECT 2704.405 86.170 2704.735 86.185 ;
        RECT 2656.310 85.870 2704.735 86.170 ;
        RECT 2656.310 85.860 2656.690 85.870 ;
        RECT 2704.405 85.855 2704.735 85.870 ;
        RECT 2053.505 85.490 2053.835 85.505 ;
        RECT 2090.305 85.490 2090.635 85.505 ;
        RECT 2510.030 85.490 2510.410 85.500 ;
        RECT 2752.910 85.490 2753.290 85.500 ;
        RECT 2053.505 85.190 2090.635 85.490 ;
        RECT 2053.505 85.175 2053.835 85.190 ;
        RECT 2090.305 85.175 2090.635 85.190 ;
        RECT 2476.030 85.190 2510.410 85.490 ;
        RECT 1297.470 84.810 1297.850 84.820 ;
        RECT 1393.865 84.810 1394.195 84.825 ;
        RECT 1255.190 84.510 1297.850 84.810 ;
        RECT 1158.550 84.130 1158.930 84.140 ;
        RECT 1220.905 84.130 1221.235 84.145 ;
        RECT 1158.550 83.830 1221.235 84.130 ;
        RECT 1158.550 83.820 1158.930 83.830 ;
        RECT 1220.905 83.815 1221.235 83.830 ;
        RECT 1221.825 84.130 1222.155 84.145 ;
        RECT 1255.190 84.130 1255.490 84.510 ;
        RECT 1297.470 84.500 1297.850 84.510 ;
        RECT 1351.790 84.510 1394.195 84.810 ;
        RECT 1221.825 83.830 1255.490 84.130 ;
        RECT 1345.105 84.130 1345.435 84.145 ;
        RECT 1351.790 84.130 1352.090 84.510 ;
        RECT 1393.865 84.495 1394.195 84.510 ;
        RECT 1617.885 84.810 1618.215 84.825 ;
        RECT 1628.670 84.810 1629.050 84.820 ;
        RECT 1617.885 84.510 1629.050 84.810 ;
        RECT 1617.885 84.495 1618.215 84.510 ;
        RECT 1628.670 84.500 1629.050 84.510 ;
        RECT 1779.805 84.810 1780.135 84.825 ;
        RECT 1786.910 84.810 1787.290 84.820 ;
        RECT 2091.225 84.810 2091.555 84.825 ;
        RECT 2283.965 84.810 2284.295 84.825 ;
        RECT 1779.805 84.510 1787.290 84.810 ;
        RECT 1779.805 84.495 1780.135 84.510 ;
        RECT 1786.910 84.500 1787.290 84.510 ;
        RECT 1876.190 84.510 1907.770 84.810 ;
        RECT 1345.105 83.830 1352.090 84.130 ;
        RECT 1545.205 84.130 1545.535 84.145 ;
        RECT 1617.425 84.130 1617.755 84.145 ;
        RECT 1545.205 83.830 1559.090 84.130 ;
        RECT 1221.825 83.815 1222.155 83.830 ;
        RECT 1345.105 83.815 1345.435 83.830 ;
        RECT 1545.205 83.815 1545.535 83.830 ;
        RECT 1441.705 83.450 1442.035 83.465 ;
        RECT 1496.445 83.450 1496.775 83.465 ;
        RECT 1497.110 83.450 1497.490 83.460 ;
        RECT 1441.705 83.150 1449.610 83.450 ;
        RECT 1441.705 83.135 1442.035 83.150 ;
        RECT 1449.310 82.770 1449.610 83.150 ;
        RECT 1496.445 83.150 1497.490 83.450 ;
        RECT 1558.790 83.450 1559.090 83.830 ;
        RECT 1587.310 83.830 1617.755 84.130 ;
        RECT 1587.310 83.450 1587.610 83.830 ;
        RECT 1617.425 83.815 1617.755 83.830 ;
        RECT 1676.305 84.130 1676.635 84.145 ;
        RECT 1852.485 84.130 1852.815 84.145 ;
        RECT 1876.190 84.130 1876.490 84.510 ;
        RECT 1676.305 83.830 1689.730 84.130 ;
        RECT 1676.305 83.815 1676.635 83.830 ;
        RECT 1558.790 83.150 1587.610 83.450 ;
        RECT 1689.430 83.450 1689.730 83.830 ;
        RECT 1852.485 83.830 1876.490 84.130 ;
        RECT 1907.470 84.130 1907.770 84.510 ;
        RECT 2091.225 84.510 2138.690 84.810 ;
        RECT 2091.225 84.495 2091.555 84.510 ;
        RECT 1932.525 84.130 1932.855 84.145 ;
        RECT 1907.470 83.830 1932.855 84.130 ;
        RECT 1852.485 83.815 1852.815 83.830 ;
        RECT 1932.525 83.815 1932.855 83.830 ;
        RECT 1994.625 84.130 1994.955 84.145 ;
        RECT 2042.005 84.130 2042.335 84.145 ;
        RECT 1994.625 83.830 2042.335 84.130 ;
        RECT 1994.625 83.815 1994.955 83.830 ;
        RECT 2042.005 83.815 2042.335 83.830 ;
        RECT 1731.045 83.450 1731.375 83.465 ;
        RECT 1738.405 83.450 1738.735 83.465 ;
        RECT 1689.430 83.150 1731.375 83.450 ;
        RECT 1496.445 83.135 1496.775 83.150 ;
        RECT 1497.110 83.140 1497.490 83.150 ;
        RECT 1731.045 83.135 1731.375 83.150 ;
        RECT 1731.750 83.150 1738.735 83.450 ;
        RECT 1496.445 82.770 1496.775 82.785 ;
        RECT 1449.310 82.470 1496.775 82.770 ;
        RECT 1496.445 82.455 1496.775 82.470 ;
        RECT 1731.045 82.770 1731.375 82.785 ;
        RECT 1731.750 82.770 1732.050 83.150 ;
        RECT 1738.405 83.135 1738.735 83.150 ;
        RECT 1787.830 83.450 1788.210 83.460 ;
        RECT 1828.310 83.450 1828.690 83.460 ;
        RECT 1787.830 83.150 1828.690 83.450 ;
        RECT 2138.390 83.450 2138.690 84.510 ;
        RECT 2139.310 84.510 2187.450 84.810 ;
        RECT 2139.310 83.450 2139.610 84.510 ;
        RECT 2138.390 83.150 2139.610 83.450 ;
        RECT 2187.150 83.450 2187.450 84.510 ;
        RECT 2283.965 84.510 2284.970 84.810 ;
        RECT 2283.965 84.495 2284.295 84.510 ;
        RECT 2283.505 84.130 2283.835 84.145 ;
        RECT 2235.910 83.830 2283.835 84.130 ;
        RECT 2284.670 84.130 2284.970 84.510 ;
        RECT 2379.645 84.130 2379.975 84.145 ;
        RECT 2284.670 83.830 2331.890 84.130 ;
        RECT 2235.910 83.450 2236.210 83.830 ;
        RECT 2283.505 83.815 2283.835 83.830 ;
        RECT 2187.150 83.150 2236.210 83.450 ;
        RECT 2331.590 83.450 2331.890 83.830 ;
        RECT 2332.510 83.830 2379.975 84.130 ;
        RECT 2332.510 83.450 2332.810 83.830 ;
        RECT 2379.645 83.815 2379.975 83.830 ;
        RECT 2387.465 84.130 2387.795 84.145 ;
        RECT 2476.030 84.130 2476.330 85.190 ;
        RECT 2510.030 85.180 2510.410 85.190 ;
        RECT 2718.910 85.190 2753.290 85.490 ;
        RECT 2622.525 84.810 2622.855 84.825 ;
        RECT 2656.310 84.810 2656.690 84.820 ;
        RECT 2622.525 84.510 2656.690 84.810 ;
        RECT 2622.525 84.495 2622.855 84.510 ;
        RECT 2656.310 84.500 2656.690 84.510 ;
        RECT 2572.845 84.130 2573.175 84.145 ;
        RECT 2387.465 83.830 2414.690 84.130 ;
        RECT 2387.465 83.815 2387.795 83.830 ;
        RECT 2331.590 83.150 2332.810 83.450 ;
        RECT 2414.390 83.450 2414.690 83.830 ;
        RECT 2429.110 83.830 2476.330 84.130 ;
        RECT 2525.710 83.830 2573.175 84.130 ;
        RECT 2429.110 83.450 2429.410 83.830 ;
        RECT 2414.390 83.150 2429.410 83.450 ;
        RECT 2510.950 83.450 2511.330 83.460 ;
        RECT 2525.710 83.450 2526.010 83.830 ;
        RECT 2572.845 83.815 2573.175 83.830 ;
        RECT 2704.405 84.130 2704.735 84.145 ;
        RECT 2718.910 84.130 2719.210 85.190 ;
        RECT 2752.910 85.180 2753.290 85.190 ;
        RECT 2801.005 84.810 2801.335 84.825 ;
        RECT 2801.005 84.510 2815.810 84.810 ;
        RECT 2801.005 84.495 2801.335 84.510 ;
        RECT 2704.405 83.830 2719.210 84.130 ;
        RECT 2704.405 83.815 2704.735 83.830 ;
        RECT 2608.265 83.450 2608.595 83.465 ;
        RECT 2510.950 83.150 2526.010 83.450 ;
        RECT 2607.590 83.150 2608.595 83.450 ;
        RECT 2815.510 83.450 2815.810 84.510 ;
        RECT 2863.105 84.130 2863.435 84.145 ;
        RECT 2916.710 84.130 2917.010 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
        RECT 2849.550 83.830 2863.435 84.130 ;
        RECT 2849.550 83.450 2849.850 83.830 ;
        RECT 2863.105 83.815 2863.435 83.830 ;
        RECT 2884.510 83.830 2917.010 84.130 ;
        RECT 2815.510 83.150 2849.850 83.450 ;
        RECT 2863.565 83.450 2863.895 83.465 ;
        RECT 2884.510 83.450 2884.810 83.830 ;
        RECT 2863.565 83.150 2884.810 83.450 ;
        RECT 1787.830 83.140 1788.210 83.150 ;
        RECT 1828.310 83.140 1828.690 83.150 ;
        RECT 2510.950 83.140 2511.330 83.150 ;
        RECT 1731.045 82.470 1732.050 82.770 ;
        RECT 1932.525 82.770 1932.855 82.785 ;
        RECT 1979.190 82.770 1979.570 82.780 ;
        RECT 1932.525 82.470 1979.570 82.770 ;
        RECT 1731.045 82.455 1731.375 82.470 ;
        RECT 1932.525 82.455 1932.855 82.470 ;
        RECT 1979.190 82.460 1979.570 82.470 ;
        RECT 1980.110 82.770 1980.490 82.780 ;
        RECT 1994.625 82.770 1994.955 82.785 ;
        RECT 1980.110 82.470 1994.955 82.770 ;
        RECT 1980.110 82.460 1980.490 82.470 ;
        RECT 1994.625 82.455 1994.955 82.470 ;
        RECT 1497.110 82.090 1497.490 82.100 ;
        RECT 1545.205 82.090 1545.535 82.105 ;
        RECT 1497.110 81.790 1545.535 82.090 ;
        RECT 1497.110 81.780 1497.490 81.790 ;
        RECT 1545.205 81.775 1545.535 81.790 ;
        RECT 1828.310 82.090 1828.690 82.100 ;
        RECT 1852.485 82.090 1852.815 82.105 ;
        RECT 1828.310 81.790 1852.815 82.090 ;
        RECT 1828.310 81.780 1828.690 81.790 ;
        RECT 1852.485 81.775 1852.815 81.790 ;
        RECT 2572.845 82.090 2573.175 82.105 ;
        RECT 2607.590 82.090 2607.890 83.150 ;
        RECT 2608.265 83.135 2608.595 83.150 ;
        RECT 2863.565 83.135 2863.895 83.150 ;
        RECT 2572.845 81.790 2607.890 82.090 ;
        RECT 2572.845 81.775 2573.175 81.790 ;
      LAYER via3 ;
        RECT 1158.580 3199.580 1158.900 3199.900 ;
        RECT 2752.940 86.540 2753.260 86.860 ;
        RECT 1297.500 85.860 1297.820 86.180 ;
        RECT 1628.700 85.860 1629.020 86.180 ;
        RECT 2656.340 85.860 2656.660 86.180 ;
        RECT 1158.580 83.820 1158.900 84.140 ;
        RECT 1297.500 84.500 1297.820 84.820 ;
        RECT 1628.700 84.500 1629.020 84.820 ;
        RECT 1786.940 84.500 1787.260 84.820 ;
        RECT 1497.140 83.140 1497.460 83.460 ;
        RECT 1787.860 83.140 1788.180 83.460 ;
        RECT 1828.340 83.140 1828.660 83.460 ;
        RECT 2510.060 85.180 2510.380 85.500 ;
        RECT 2656.340 84.500 2656.660 84.820 ;
        RECT 2510.980 83.140 2511.300 83.460 ;
        RECT 2752.940 85.180 2753.260 85.500 ;
        RECT 1979.220 82.460 1979.540 82.780 ;
        RECT 1980.140 82.460 1980.460 82.780 ;
        RECT 1497.140 81.780 1497.460 82.100 ;
        RECT 1828.340 81.780 1828.660 82.100 ;
      LAYER met4 ;
        RECT 1158.575 3199.575 1158.905 3199.905 ;
        RECT 1158.590 84.145 1158.890 3199.575 ;
        RECT 2752.935 86.535 2753.265 86.865 ;
        RECT 1297.495 85.855 1297.825 86.185 ;
        RECT 1628.695 85.855 1629.025 86.185 ;
        RECT 2656.335 85.855 2656.665 86.185 ;
        RECT 1297.510 84.825 1297.810 85.855 ;
        RECT 1628.710 84.825 1629.010 85.855 ;
        RECT 2510.055 85.175 2510.385 85.505 ;
        RECT 1297.495 84.495 1297.825 84.825 ;
        RECT 1628.695 84.495 1629.025 84.825 ;
        RECT 1786.935 84.495 1787.265 84.825 ;
        RECT 1158.575 83.815 1158.905 84.145 ;
        RECT 1497.135 83.135 1497.465 83.465 ;
        RECT 1786.950 83.450 1787.250 84.495 ;
        RECT 1787.855 83.450 1788.185 83.465 ;
        RECT 1786.950 83.150 1788.185 83.450 ;
        RECT 1787.855 83.135 1788.185 83.150 ;
        RECT 1828.335 83.135 1828.665 83.465 ;
        RECT 2510.070 83.450 2510.370 85.175 ;
        RECT 2656.350 84.825 2656.650 85.855 ;
        RECT 2752.950 85.505 2753.250 86.535 ;
        RECT 2752.935 85.175 2753.265 85.505 ;
        RECT 2656.335 84.495 2656.665 84.825 ;
        RECT 2510.975 83.450 2511.305 83.465 ;
        RECT 1979.230 83.150 1980.450 83.450 ;
        RECT 2510.070 83.150 2511.305 83.450 ;
        RECT 1497.150 82.105 1497.450 83.135 ;
        RECT 1828.350 82.105 1828.650 83.135 ;
        RECT 1979.230 82.785 1979.530 83.150 ;
        RECT 1980.150 82.785 1980.450 83.150 ;
        RECT 2510.975 83.135 2511.305 83.150 ;
        RECT 1979.215 82.455 1979.545 82.785 ;
        RECT 1980.135 82.455 1980.465 82.785 ;
        RECT 1497.135 81.775 1497.465 82.105 ;
        RECT 1828.335 81.775 1828.665 82.105 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1549.810 3207.120 1550.130 3207.180 ;
        RECT 2648.750 3207.120 2649.070 3207.180 ;
        RECT 1549.810 3206.980 2649.070 3207.120 ;
        RECT 1549.810 3206.920 1550.130 3206.980 ;
        RECT 2648.750 3206.920 2649.070 3206.980 ;
        RECT 2648.750 2435.660 2649.070 2435.720 ;
        RECT 2898.990 2435.660 2899.310 2435.720 ;
        RECT 2648.750 2435.520 2899.310 2435.660 ;
        RECT 2648.750 2435.460 2649.070 2435.520 ;
        RECT 2898.990 2435.460 2899.310 2435.520 ;
      LAYER via ;
        RECT 1549.840 3206.920 1550.100 3207.180 ;
        RECT 2648.780 3206.920 2649.040 3207.180 ;
        RECT 2648.780 2435.460 2649.040 2435.720 ;
        RECT 2899.020 2435.460 2899.280 2435.720 ;
      LAYER met2 ;
        RECT 1549.840 3206.890 1550.100 3207.210 ;
        RECT 2648.780 3206.890 2649.040 3207.210 ;
        RECT 1549.900 3200.000 1550.040 3206.890 ;
        RECT 1549.760 3197.600 1550.040 3200.000 ;
        RECT 2648.840 2435.750 2648.980 3206.890 ;
        RECT 2648.780 2435.430 2649.040 2435.750 ;
        RECT 2899.020 2435.430 2899.280 2435.750 ;
        RECT 2899.080 2434.245 2899.220 2435.430 ;
        RECT 2899.010 2433.875 2899.290 2434.245 ;
      LAYER via2 ;
        RECT 2899.010 2433.920 2899.290 2434.200 ;
      LAYER met3 ;
        RECT 2898.985 2434.210 2899.315 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2898.985 2433.910 2924.800 2434.210 ;
        RECT 2898.985 2433.895 2899.315 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1588.910 3207.800 1589.230 3207.860 ;
        RECT 2649.210 3207.800 2649.530 3207.860 ;
        RECT 1588.910 3207.660 2649.530 3207.800 ;
        RECT 1588.910 3207.600 1589.230 3207.660 ;
        RECT 2649.210 3207.600 2649.530 3207.660 ;
        RECT 2649.210 2670.260 2649.530 2670.320 ;
        RECT 2898.990 2670.260 2899.310 2670.320 ;
        RECT 2649.210 2670.120 2899.310 2670.260 ;
        RECT 2649.210 2670.060 2649.530 2670.120 ;
        RECT 2898.990 2670.060 2899.310 2670.120 ;
      LAYER via ;
        RECT 1588.940 3207.600 1589.200 3207.860 ;
        RECT 2649.240 3207.600 2649.500 3207.860 ;
        RECT 2649.240 2670.060 2649.500 2670.320 ;
        RECT 2899.020 2670.060 2899.280 2670.320 ;
      LAYER met2 ;
        RECT 1588.940 3207.570 1589.200 3207.890 ;
        RECT 2649.240 3207.570 2649.500 3207.890 ;
        RECT 1589.000 3200.000 1589.140 3207.570 ;
        RECT 1588.860 3197.600 1589.140 3200.000 ;
        RECT 2649.300 2670.350 2649.440 3207.570 ;
        RECT 2649.240 2670.030 2649.500 2670.350 ;
        RECT 2899.020 2670.030 2899.280 2670.350 ;
        RECT 2899.080 2669.525 2899.220 2670.030 ;
        RECT 2899.010 2669.155 2899.290 2669.525 ;
      LAYER via2 ;
        RECT 2899.010 2669.200 2899.290 2669.480 ;
      LAYER met3 ;
        RECT 2898.985 2669.490 2899.315 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2898.985 2669.190 2924.800 2669.490 ;
        RECT 2898.985 2669.175 2899.315 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1628.490 3214.515 1628.770 3214.885 ;
        RECT 1628.560 3200.000 1628.700 3214.515 ;
        RECT 1628.420 3197.600 1628.700 3200.000 ;
      LAYER via2 ;
        RECT 1628.490 3214.560 1628.770 3214.840 ;
      LAYER met3 ;
        RECT 1628.465 3214.850 1628.795 3214.865 ;
        RECT 2630.550 3214.850 2630.930 3214.860 ;
        RECT 1628.465 3214.550 2630.930 3214.850 ;
        RECT 1628.465 3214.535 1628.795 3214.550 ;
        RECT 2630.550 3214.540 2630.930 3214.550 ;
        RECT 2630.550 3189.010 2630.930 3189.020 ;
        RECT 2636.070 3189.010 2636.450 3189.020 ;
        RECT 2630.550 3188.710 2636.450 3189.010 ;
        RECT 2630.550 3188.700 2630.930 3188.710 ;
        RECT 2636.070 3188.700 2636.450 3188.710 ;
        RECT 2636.070 3172.010 2636.450 3172.020 ;
        RECT 2637.910 3172.010 2638.290 3172.020 ;
        RECT 2636.070 3171.710 2638.290 3172.010 ;
        RECT 2636.070 3171.700 2636.450 3171.710 ;
        RECT 2637.910 3171.700 2638.290 3171.710 ;
        RECT 2637.910 3153.650 2638.290 3153.660 ;
        RECT 2637.030 3153.350 2638.290 3153.650 ;
        RECT 2637.030 3152.980 2637.330 3153.350 ;
        RECT 2637.910 3153.340 2638.290 3153.350 ;
        RECT 2636.990 3152.660 2637.370 3152.980 ;
        RECT 2638.830 3139.370 2639.210 3139.380 ;
        RECT 2642.510 3139.370 2642.890 3139.380 ;
        RECT 2638.830 3139.070 2642.890 3139.370 ;
        RECT 2638.830 3139.060 2639.210 3139.070 ;
        RECT 2642.510 3139.060 2642.890 3139.070 ;
        RECT 2637.910 3091.770 2638.290 3091.780 ;
        RECT 2642.510 3091.770 2642.890 3091.780 ;
        RECT 2637.910 3091.470 2642.890 3091.770 ;
        RECT 2637.910 3091.460 2638.290 3091.470 ;
        RECT 2642.510 3091.460 2642.890 3091.470 ;
        RECT 2636.070 3090.410 2636.450 3090.420 ;
        RECT 2637.910 3090.410 2638.290 3090.420 ;
        RECT 2636.070 3090.110 2638.290 3090.410 ;
        RECT 2636.070 3090.100 2636.450 3090.110 ;
        RECT 2637.910 3090.100 2638.290 3090.110 ;
        RECT 2636.070 3043.490 2636.450 3043.500 ;
        RECT 2639.750 3043.490 2640.130 3043.500 ;
        RECT 2636.070 3043.190 2640.130 3043.490 ;
        RECT 2636.070 3043.180 2636.450 3043.190 ;
        RECT 2639.750 3043.180 2640.130 3043.190 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2916.710 2903.790 2924.800 2904.090 ;
        RECT 2691.310 2899.710 2739.450 2900.010 ;
        RECT 2636.990 2899.330 2637.370 2899.340 ;
        RECT 2636.990 2899.030 2690.690 2899.330 ;
        RECT 2636.990 2899.020 2637.370 2899.030 ;
        RECT 2690.390 2898.650 2690.690 2899.030 ;
        RECT 2691.310 2898.650 2691.610 2899.710 ;
        RECT 2739.150 2899.330 2739.450 2899.710 ;
        RECT 2787.910 2899.710 2836.050 2900.010 ;
        RECT 2739.150 2899.030 2787.290 2899.330 ;
        RECT 2690.390 2898.350 2691.610 2898.650 ;
        RECT 2786.990 2898.650 2787.290 2899.030 ;
        RECT 2787.910 2898.650 2788.210 2899.710 ;
        RECT 2835.750 2899.330 2836.050 2899.710 ;
        RECT 2835.750 2899.030 2883.890 2899.330 ;
        RECT 2786.990 2898.350 2788.210 2898.650 ;
        RECT 2883.590 2898.650 2883.890 2899.030 ;
        RECT 2916.710 2898.650 2917.010 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2883.590 2898.350 2917.010 2898.650 ;
      LAYER via3 ;
        RECT 2630.580 3214.540 2630.900 3214.860 ;
        RECT 2630.580 3188.700 2630.900 3189.020 ;
        RECT 2636.100 3188.700 2636.420 3189.020 ;
        RECT 2636.100 3171.700 2636.420 3172.020 ;
        RECT 2637.940 3171.700 2638.260 3172.020 ;
        RECT 2637.940 3153.340 2638.260 3153.660 ;
        RECT 2637.020 3152.660 2637.340 3152.980 ;
        RECT 2638.860 3139.060 2639.180 3139.380 ;
        RECT 2642.540 3139.060 2642.860 3139.380 ;
        RECT 2637.940 3091.460 2638.260 3091.780 ;
        RECT 2642.540 3091.460 2642.860 3091.780 ;
        RECT 2636.100 3090.100 2636.420 3090.420 ;
        RECT 2637.940 3090.100 2638.260 3090.420 ;
        RECT 2636.100 3043.180 2636.420 3043.500 ;
        RECT 2639.780 3043.180 2640.100 3043.500 ;
        RECT 2637.020 2899.020 2637.340 2899.340 ;
      LAYER met4 ;
        RECT 2630.575 3214.535 2630.905 3214.865 ;
        RECT 2630.590 3189.025 2630.890 3214.535 ;
        RECT 2630.575 3188.695 2630.905 3189.025 ;
        RECT 2636.095 3188.695 2636.425 3189.025 ;
        RECT 2636.110 3172.025 2636.410 3188.695 ;
        RECT 2636.095 3171.695 2636.425 3172.025 ;
        RECT 2637.935 3171.695 2638.265 3172.025 ;
        RECT 2637.950 3153.665 2638.250 3171.695 ;
        RECT 2637.935 3153.335 2638.265 3153.665 ;
        RECT 2637.015 3152.655 2637.345 3152.985 ;
        RECT 2637.030 3140.050 2637.330 3152.655 ;
        RECT 2637.030 3139.750 2639.170 3140.050 ;
        RECT 2638.870 3139.385 2639.170 3139.750 ;
        RECT 2638.855 3139.055 2639.185 3139.385 ;
        RECT 2642.535 3139.055 2642.865 3139.385 ;
        RECT 2642.550 3091.785 2642.850 3139.055 ;
        RECT 2637.935 3091.455 2638.265 3091.785 ;
        RECT 2642.535 3091.455 2642.865 3091.785 ;
        RECT 2637.950 3090.425 2638.250 3091.455 ;
        RECT 2636.095 3090.095 2636.425 3090.425 ;
        RECT 2637.935 3090.095 2638.265 3090.425 ;
        RECT 2636.110 3043.505 2636.410 3090.095 ;
        RECT 2636.095 3043.175 2636.425 3043.505 ;
        RECT 2639.775 3043.175 2640.105 3043.505 ;
        RECT 2639.790 2946.250 2640.090 3043.175 ;
        RECT 2637.950 2945.950 2640.090 2946.250 ;
        RECT 2637.950 2912.250 2638.250 2945.950 ;
        RECT 2637.030 2911.950 2638.250 2912.250 ;
        RECT 2637.030 2899.345 2637.330 2911.950 ;
        RECT 2637.015 2899.015 2637.345 2899.345 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1668.030 3208.140 1668.350 3208.200 ;
        RECT 2651.050 3208.140 2651.370 3208.200 ;
        RECT 1668.030 3208.000 2651.370 3208.140 ;
        RECT 1668.030 3207.940 1668.350 3208.000 ;
        RECT 2651.050 3207.940 2651.370 3208.000 ;
        RECT 2651.050 3139.460 2651.370 3139.520 ;
        RECT 2898.990 3139.460 2899.310 3139.520 ;
        RECT 2651.050 3139.320 2899.310 3139.460 ;
        RECT 2651.050 3139.260 2651.370 3139.320 ;
        RECT 2898.990 3139.260 2899.310 3139.320 ;
      LAYER via ;
        RECT 1668.060 3207.940 1668.320 3208.200 ;
        RECT 2651.080 3207.940 2651.340 3208.200 ;
        RECT 2651.080 3139.260 2651.340 3139.520 ;
        RECT 2899.020 3139.260 2899.280 3139.520 ;
      LAYER met2 ;
        RECT 1668.060 3207.910 1668.320 3208.230 ;
        RECT 2651.080 3207.910 2651.340 3208.230 ;
        RECT 1668.120 3200.000 1668.260 3207.910 ;
        RECT 1667.980 3197.600 1668.260 3200.000 ;
        RECT 2651.140 3139.550 2651.280 3207.910 ;
        RECT 2651.080 3139.230 2651.340 3139.550 ;
        RECT 2899.020 3139.230 2899.280 3139.550 ;
        RECT 2899.080 3138.725 2899.220 3139.230 ;
        RECT 2899.010 3138.355 2899.290 3138.725 ;
      LAYER via2 ;
        RECT 2899.010 3138.400 2899.290 3138.680 ;
      LAYER met3 ;
        RECT 2898.985 3138.690 2899.315 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2898.985 3138.390 2924.800 3138.690 ;
        RECT 2898.985 3138.375 2899.315 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 3367.600 1711.130 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1710.810 3367.460 2901.150 3367.600 ;
        RECT 1710.810 3367.400 1711.130 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 1710.840 3367.400 1711.100 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1710.840 3367.370 1711.100 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1707.540 3199.130 1707.820 3200.000 ;
        RECT 1710.900 3199.810 1711.040 3367.370 ;
        RECT 1709.980 3199.670 1711.040 3199.810 ;
        RECT 1709.980 3199.130 1710.120 3199.670 ;
        RECT 1707.540 3198.990 1710.120 3199.130 ;
        RECT 1707.540 3197.600 1707.820 3198.990 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3422.355 ;
        RECT 2796.025 3236.205 2796.195 3284.315 ;
      LAYER mcon ;
        RECT 2796.485 3422.185 2796.655 3422.355 ;
        RECT 2796.025 3284.145 2796.195 3284.315 ;
      LAYER met1 ;
        RECT 2795.490 3443.080 2795.810 3443.140 ;
        RECT 2798.250 3443.080 2798.570 3443.140 ;
        RECT 2795.490 3442.940 2798.570 3443.080 ;
        RECT 2795.490 3442.880 2795.810 3442.940 ;
        RECT 2798.250 3442.880 2798.570 3442.940 ;
        RECT 2795.030 3422.340 2795.350 3422.400 ;
        RECT 2796.425 3422.340 2796.715 3422.385 ;
        RECT 2795.030 3422.200 2796.715 3422.340 ;
        RECT 2795.030 3422.140 2795.350 3422.200 ;
        RECT 2796.425 3422.155 2796.715 3422.200 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.950 3284.300 2796.270 3284.360 ;
        RECT 2795.755 3284.160 2796.270 3284.300 ;
        RECT 2795.950 3284.100 2796.270 3284.160 ;
        RECT 2795.965 3236.360 2796.255 3236.405 ;
        RECT 2796.410 3236.360 2796.730 3236.420 ;
        RECT 2795.965 3236.220 2796.730 3236.360 ;
        RECT 2795.965 3236.175 2796.255 3236.220 ;
        RECT 2796.410 3236.160 2796.730 3236.220 ;
        RECT 1747.150 3218.680 1747.470 3218.740 ;
        RECT 2796.410 3218.680 2796.730 3218.740 ;
        RECT 1747.150 3218.540 2796.730 3218.680 ;
        RECT 1747.150 3218.480 1747.470 3218.540 ;
        RECT 2796.410 3218.480 2796.730 3218.540 ;
      LAYER via ;
        RECT 2795.520 3442.880 2795.780 3443.140 ;
        RECT 2798.280 3442.880 2798.540 3443.140 ;
        RECT 2795.060 3422.140 2795.320 3422.400 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.980 3284.100 2796.240 3284.360 ;
        RECT 2796.440 3236.160 2796.700 3236.420 ;
        RECT 1747.180 3218.480 1747.440 3218.740 ;
        RECT 2796.440 3218.480 2796.700 3218.740 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3443.170 2798.480 3517.600 ;
        RECT 2795.520 3442.850 2795.780 3443.170 ;
        RECT 2798.280 3442.850 2798.540 3443.170 ;
        RECT 2795.580 3429.650 2795.720 3442.850 ;
        RECT 2795.120 3429.510 2795.720 3429.650 ;
        RECT 2795.120 3422.430 2795.260 3429.510 ;
        RECT 2795.060 3422.110 2795.320 3422.430 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3284.390 2796.180 3298.270 ;
        RECT 2795.980 3284.070 2796.240 3284.390 ;
        RECT 2796.440 3236.130 2796.700 3236.450 ;
        RECT 2796.500 3218.770 2796.640 3236.130 ;
        RECT 1747.180 3218.450 1747.440 3218.770 ;
        RECT 2796.440 3218.450 2796.700 3218.770 ;
        RECT 1747.240 3200.000 1747.380 3218.450 ;
        RECT 1747.100 3197.600 1747.380 3200.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 1786.710 3219.360 1787.030 3219.420 ;
        RECT 2470.270 3219.360 2470.590 3219.420 ;
        RECT 1786.710 3219.220 2470.590 3219.360 ;
        RECT 1786.710 3219.160 1787.030 3219.220 ;
        RECT 2470.270 3219.160 2470.590 3219.220 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 1786.740 3219.160 1787.000 3219.420 ;
        RECT 2470.300 3219.160 2470.560 3219.420 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3430.445 2474.640 3517.230 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3219.450 2470.500 3270.470 ;
        RECT 1786.740 3219.130 1787.000 3219.450 ;
        RECT 2470.300 3219.130 2470.560 3219.450 ;
        RECT 1786.800 3200.000 1786.940 3219.130 ;
        RECT 1786.660 3197.600 1786.940 3200.000 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.425 3332.765 2147.595 3422.355 ;
        RECT 2146.045 3236.205 2146.215 3284.315 ;
      LAYER mcon ;
        RECT 2147.425 3422.185 2147.595 3422.355 ;
        RECT 2146.045 3284.145 2146.215 3284.315 ;
      LAYER met1 ;
        RECT 2146.890 3443.080 2147.210 3443.140 ;
        RECT 2149.190 3443.080 2149.510 3443.140 ;
        RECT 2146.890 3442.940 2149.510 3443.080 ;
        RECT 2146.890 3442.880 2147.210 3442.940 ;
        RECT 2149.190 3442.880 2149.510 3442.940 ;
        RECT 2146.430 3422.340 2146.750 3422.400 ;
        RECT 2147.365 3422.340 2147.655 3422.385 ;
        RECT 2146.430 3422.200 2147.655 3422.340 ;
        RECT 2146.430 3422.140 2146.750 3422.200 ;
        RECT 2147.365 3422.155 2147.655 3422.200 ;
        RECT 2147.350 3332.920 2147.670 3332.980 ;
        RECT 2147.155 3332.780 2147.670 3332.920 ;
        RECT 2147.350 3332.720 2147.670 3332.780 ;
        RECT 2145.985 3284.300 2146.275 3284.345 ;
        RECT 2146.430 3284.300 2146.750 3284.360 ;
        RECT 2145.985 3284.160 2146.750 3284.300 ;
        RECT 2145.985 3284.115 2146.275 3284.160 ;
        RECT 2146.430 3284.100 2146.750 3284.160 ;
        RECT 2145.970 3236.360 2146.290 3236.420 ;
        RECT 2145.775 3236.220 2146.290 3236.360 ;
        RECT 2145.970 3236.160 2146.290 3236.220 ;
        RECT 1825.810 3220.040 1826.130 3220.100 ;
        RECT 2145.970 3220.040 2146.290 3220.100 ;
        RECT 1825.810 3219.900 2146.290 3220.040 ;
        RECT 1825.810 3219.840 1826.130 3219.900 ;
        RECT 2145.970 3219.840 2146.290 3219.900 ;
      LAYER via ;
        RECT 2146.920 3442.880 2147.180 3443.140 ;
        RECT 2149.220 3442.880 2149.480 3443.140 ;
        RECT 2146.460 3422.140 2146.720 3422.400 ;
        RECT 2147.380 3332.720 2147.640 3332.980 ;
        RECT 2146.460 3284.100 2146.720 3284.360 ;
        RECT 2146.000 3236.160 2146.260 3236.420 ;
        RECT 1825.840 3219.840 1826.100 3220.100 ;
        RECT 2146.000 3219.840 2146.260 3220.100 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3443.170 2149.420 3517.600 ;
        RECT 2146.920 3442.850 2147.180 3443.170 ;
        RECT 2149.220 3442.850 2149.480 3443.170 ;
        RECT 2146.980 3429.650 2147.120 3442.850 ;
        RECT 2146.520 3429.510 2147.120 3429.650 ;
        RECT 2146.520 3422.430 2146.660 3429.510 ;
        RECT 2146.460 3422.110 2146.720 3422.430 ;
        RECT 2147.380 3332.690 2147.640 3333.010 ;
        RECT 2147.440 3298.410 2147.580 3332.690 ;
        RECT 2146.520 3298.270 2147.580 3298.410 ;
        RECT 2146.520 3284.390 2146.660 3298.270 ;
        RECT 2146.460 3284.070 2146.720 3284.390 ;
        RECT 2146.000 3236.130 2146.260 3236.450 ;
        RECT 2146.060 3220.130 2146.200 3236.130 ;
        RECT 1825.840 3219.810 1826.100 3220.130 ;
        RECT 2146.000 3219.810 2146.260 3220.130 ;
        RECT 1825.900 3200.000 1826.040 3219.810 ;
        RECT 1825.760 3197.600 1826.040 3200.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3498.500 1825.210 3498.560 ;
        RECT 1828.110 3498.500 1828.430 3498.560 ;
        RECT 1824.890 3498.360 1828.430 3498.500 ;
        RECT 1824.890 3498.300 1825.210 3498.360 ;
        RECT 1828.110 3498.300 1828.430 3498.360 ;
        RECT 1828.110 3215.620 1828.430 3215.680 ;
        RECT 1865.370 3215.620 1865.690 3215.680 ;
        RECT 1828.110 3215.480 1865.690 3215.620 ;
        RECT 1828.110 3215.420 1828.430 3215.480 ;
        RECT 1865.370 3215.420 1865.690 3215.480 ;
      LAYER via ;
        RECT 1824.920 3498.300 1825.180 3498.560 ;
        RECT 1828.140 3498.300 1828.400 3498.560 ;
        RECT 1828.140 3215.420 1828.400 3215.680 ;
        RECT 1865.400 3215.420 1865.660 3215.680 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3498.590 1825.120 3517.600 ;
        RECT 1824.920 3498.270 1825.180 3498.590 ;
        RECT 1828.140 3498.270 1828.400 3498.590 ;
        RECT 1828.200 3215.710 1828.340 3498.270 ;
        RECT 1828.140 3215.390 1828.400 3215.710 ;
        RECT 1865.400 3215.390 1865.660 3215.710 ;
        RECT 1865.460 3200.000 1865.600 3215.390 ;
        RECT 1865.320 3197.600 1865.600 3200.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 3219.700 1504.130 3219.760 ;
        RECT 1904.930 3219.700 1905.250 3219.760 ;
        RECT 1503.810 3219.560 1905.250 3219.700 ;
        RECT 1503.810 3219.500 1504.130 3219.560 ;
        RECT 1904.930 3219.500 1905.250 3219.560 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 3219.500 1504.100 3219.760 ;
        RECT 1904.960 3219.500 1905.220 3219.760 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 3219.790 1504.040 3498.270 ;
        RECT 1503.840 3219.470 1504.100 3219.790 ;
        RECT 1904.960 3219.470 1905.220 3219.790 ;
        RECT 1905.020 3200.000 1905.160 3219.470 ;
        RECT 1904.880 3197.600 1905.160 3200.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1194.230 3204.740 1194.550 3204.800 ;
        RECT 2647.370 3204.740 2647.690 3204.800 ;
        RECT 1194.230 3204.600 2647.690 3204.740 ;
        RECT 1194.230 3204.540 1194.550 3204.600 ;
        RECT 2647.370 3204.540 2647.690 3204.600 ;
        RECT 2647.370 324.260 2647.690 324.320 ;
        RECT 2900.830 324.260 2901.150 324.320 ;
        RECT 2647.370 324.120 2901.150 324.260 ;
        RECT 2647.370 324.060 2647.690 324.120 ;
        RECT 2900.830 324.060 2901.150 324.120 ;
      LAYER via ;
        RECT 1194.260 3204.540 1194.520 3204.800 ;
        RECT 2647.400 3204.540 2647.660 3204.800 ;
        RECT 2647.400 324.060 2647.660 324.320 ;
        RECT 2900.860 324.060 2901.120 324.320 ;
      LAYER met2 ;
        RECT 1194.260 3204.510 1194.520 3204.830 ;
        RECT 2647.400 3204.510 2647.660 3204.830 ;
        RECT 1194.320 3200.000 1194.460 3204.510 ;
        RECT 1194.180 3197.600 1194.460 3200.000 ;
        RECT 2647.460 324.350 2647.600 3204.510 ;
        RECT 2647.400 324.030 2647.660 324.350 ;
        RECT 2900.860 324.030 2901.120 324.350 ;
        RECT 2900.920 322.845 2901.060 324.030 ;
        RECT 2900.850 322.475 2901.130 322.845 ;
      LAYER via2 ;
        RECT 2900.850 322.520 2901.130 322.800 ;
      LAYER met3 ;
        RECT 2900.825 322.810 2901.155 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2900.825 322.510 2924.800 322.810 ;
        RECT 2900.825 322.495 2901.155 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 3219.020 1179.830 3219.080 ;
        RECT 1944.490 3219.020 1944.810 3219.080 ;
        RECT 1179.510 3218.880 1944.810 3219.020 ;
        RECT 1179.510 3218.820 1179.830 3218.880 ;
        RECT 1944.490 3218.820 1944.810 3218.880 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 3218.820 1179.800 3219.080 ;
        RECT 1944.520 3218.820 1944.780 3219.080 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 3219.110 1179.740 3498.270 ;
        RECT 1179.540 3218.790 1179.800 3219.110 ;
        RECT 1944.520 3218.790 1944.780 3219.110 ;
        RECT 1944.580 3200.000 1944.720 3218.790 ;
        RECT 1944.440 3197.600 1944.720 3200.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3503.940 851.850 3504.000 ;
        RECT 1980.370 3503.940 1980.690 3504.000 ;
        RECT 851.530 3503.800 1980.690 3503.940 ;
        RECT 851.530 3503.740 851.850 3503.800 ;
        RECT 1980.370 3503.740 1980.690 3503.800 ;
      LAYER via ;
        RECT 851.560 3503.740 851.820 3504.000 ;
        RECT 1980.400 3503.740 1980.660 3504.000 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3504.030 851.760 3517.600 ;
        RECT 851.560 3503.710 851.820 3504.030 ;
        RECT 1980.400 3503.710 1980.660 3504.030 ;
        RECT 1980.460 3199.130 1980.600 3503.710 ;
        RECT 1984.000 3199.130 1984.280 3200.000 ;
        RECT 1980.460 3198.990 1984.280 3199.130 ;
        RECT 1984.000 3197.600 1984.280 3198.990 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3502.920 527.550 3502.980 ;
        RECT 2021.770 3502.920 2022.090 3502.980 ;
        RECT 527.230 3502.780 2022.090 3502.920 ;
        RECT 527.230 3502.720 527.550 3502.780 ;
        RECT 2021.770 3502.720 2022.090 3502.780 ;
      LAYER via ;
        RECT 527.260 3502.720 527.520 3502.980 ;
        RECT 2021.800 3502.720 2022.060 3502.980 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.010 527.460 3517.600 ;
        RECT 527.260 3502.690 527.520 3503.010 ;
        RECT 2021.800 3502.690 2022.060 3503.010 ;
        RECT 2021.860 3199.810 2022.000 3502.690 ;
        RECT 2023.100 3199.810 2023.380 3200.000 ;
        RECT 2021.860 3199.670 2023.380 3199.810 ;
        RECT 2023.100 3197.600 2023.380 3199.670 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 2056.270 3501.900 2056.590 3501.960 ;
        RECT 202.470 3501.760 2056.590 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 2056.270 3501.700 2056.590 3501.760 ;
        RECT 2056.270 3225.820 2056.590 3225.880 ;
        RECT 2062.710 3225.820 2063.030 3225.880 ;
        RECT 2056.270 3225.680 2063.030 3225.820 ;
        RECT 2056.270 3225.620 2056.590 3225.680 ;
        RECT 2062.710 3225.620 2063.030 3225.680 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 2056.300 3501.700 2056.560 3501.960 ;
        RECT 2056.300 3225.620 2056.560 3225.880 ;
        RECT 2062.740 3225.620 2063.000 3225.880 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 2056.300 3501.670 2056.560 3501.990 ;
        RECT 2056.360 3225.910 2056.500 3501.670 ;
        RECT 2056.300 3225.590 2056.560 3225.910 ;
        RECT 2062.740 3225.590 2063.000 3225.910 ;
        RECT 2062.800 3200.000 2062.940 3225.590 ;
        RECT 2062.660 3197.600 2062.940 3200.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 2097.670 3408.740 2097.990 3408.800 ;
        RECT 17.550 3408.600 2097.990 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 2097.670 3408.540 2097.990 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 2097.700 3408.540 2097.960 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 2097.700 3408.510 2097.960 3408.830 ;
        RECT 2097.760 3200.490 2097.900 3408.510 ;
        RECT 2097.760 3200.350 2100.660 3200.490 ;
        RECT 2100.520 3199.810 2100.660 3200.350 ;
        RECT 2102.220 3199.810 2102.500 3200.000 ;
        RECT 2100.520 3199.670 2102.500 3199.810 ;
        RECT 2102.220 3197.600 2102.500 3199.670 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 41.010 3204.400 41.330 3204.460 ;
        RECT 2141.830 3204.400 2142.150 3204.460 ;
        RECT 41.010 3204.260 2142.150 3204.400 ;
        RECT 41.010 3204.200 41.330 3204.260 ;
        RECT 2141.830 3204.200 2142.150 3204.260 ;
        RECT 16.170 3124.500 16.490 3124.560 ;
        RECT 41.010 3124.500 41.330 3124.560 ;
        RECT 16.170 3124.360 41.330 3124.500 ;
        RECT 16.170 3124.300 16.490 3124.360 ;
        RECT 41.010 3124.300 41.330 3124.360 ;
      LAYER via ;
        RECT 41.040 3204.200 41.300 3204.460 ;
        RECT 2141.860 3204.200 2142.120 3204.460 ;
        RECT 16.200 3124.300 16.460 3124.560 ;
        RECT 41.040 3124.300 41.300 3124.560 ;
      LAYER met2 ;
        RECT 41.040 3204.170 41.300 3204.490 ;
        RECT 2141.860 3204.170 2142.120 3204.490 ;
        RECT 41.100 3124.590 41.240 3204.170 ;
        RECT 2141.920 3200.000 2142.060 3204.170 ;
        RECT 2141.780 3197.600 2142.060 3200.000 ;
        RECT 16.200 3124.445 16.460 3124.590 ;
        RECT 16.190 3124.075 16.470 3124.445 ;
        RECT 41.040 3124.270 41.300 3124.590 ;
      LAYER via2 ;
        RECT 16.190 3124.120 16.470 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 16.165 3124.410 16.495 3124.425 ;
        RECT -4.800 3124.110 16.495 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 16.165 3124.095 16.495 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 40.090 3203.720 40.410 3203.780 ;
        RECT 2181.390 3203.720 2181.710 3203.780 ;
        RECT 40.090 3203.580 2181.710 3203.720 ;
        RECT 40.090 3203.520 40.410 3203.580 ;
        RECT 2181.390 3203.520 2181.710 3203.580 ;
        RECT 16.170 2838.900 16.490 2838.960 ;
        RECT 40.090 2838.900 40.410 2838.960 ;
        RECT 16.170 2838.760 40.410 2838.900 ;
        RECT 16.170 2838.700 16.490 2838.760 ;
        RECT 40.090 2838.700 40.410 2838.760 ;
      LAYER via ;
        RECT 40.120 3203.520 40.380 3203.780 ;
        RECT 2181.420 3203.520 2181.680 3203.780 ;
        RECT 16.200 2838.700 16.460 2838.960 ;
        RECT 40.120 2838.700 40.380 2838.960 ;
      LAYER met2 ;
        RECT 40.120 3203.490 40.380 3203.810 ;
        RECT 2181.420 3203.490 2181.680 3203.810 ;
        RECT 40.180 2838.990 40.320 3203.490 ;
        RECT 2181.480 3200.000 2181.620 3203.490 ;
        RECT 2181.340 3197.600 2181.620 3200.000 ;
        RECT 16.200 2838.670 16.460 2838.990 ;
        RECT 40.120 2838.670 40.380 2838.990 ;
        RECT 16.260 2836.805 16.400 2838.670 ;
        RECT 16.190 2836.435 16.470 2836.805 ;
      LAYER via2 ;
        RECT 16.190 2836.480 16.470 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 16.165 2836.770 16.495 2836.785 ;
        RECT -4.800 2836.470 16.495 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 16.165 2836.455 16.495 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2220.950 3204.060 2221.270 3204.120 ;
        RECT 2204.020 3203.920 2221.270 3204.060 ;
        RECT 32.730 3203.380 33.050 3203.440 ;
        RECT 2204.020 3203.380 2204.160 3203.920 ;
        RECT 2220.950 3203.860 2221.270 3203.920 ;
        RECT 32.730 3203.240 2204.160 3203.380 ;
        RECT 32.730 3203.180 33.050 3203.240 ;
        RECT 16.170 2551.940 16.490 2552.000 ;
        RECT 32.730 2551.940 33.050 2552.000 ;
        RECT 16.170 2551.800 33.050 2551.940 ;
        RECT 16.170 2551.740 16.490 2551.800 ;
        RECT 32.730 2551.740 33.050 2551.800 ;
      LAYER via ;
        RECT 32.760 3203.180 33.020 3203.440 ;
        RECT 2220.980 3203.860 2221.240 3204.120 ;
        RECT 16.200 2551.740 16.460 2552.000 ;
        RECT 32.760 2551.740 33.020 2552.000 ;
      LAYER met2 ;
        RECT 2220.980 3203.830 2221.240 3204.150 ;
        RECT 32.760 3203.150 33.020 3203.470 ;
        RECT 32.820 2552.030 32.960 3203.150 ;
        RECT 2221.040 3200.000 2221.180 3203.830 ;
        RECT 2220.900 3197.600 2221.180 3200.000 ;
        RECT 16.200 2551.710 16.460 2552.030 ;
        RECT 32.760 2551.710 33.020 2552.030 ;
        RECT 16.260 2549.845 16.400 2551.710 ;
        RECT 16.190 2549.475 16.470 2549.845 ;
      LAYER via2 ;
        RECT 16.190 2549.520 16.470 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 16.165 2549.810 16.495 2549.825 ;
        RECT -4.800 2549.510 16.495 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 16.165 2549.495 16.495 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 3203.040 32.590 3203.100 ;
        RECT 2260.050 3203.040 2260.370 3203.100 ;
        RECT 32.270 3202.900 2260.370 3203.040 ;
        RECT 32.270 3202.840 32.590 3202.900 ;
        RECT 2260.050 3202.840 2260.370 3202.900 ;
        RECT 15.710 2262.260 16.030 2262.320 ;
        RECT 32.270 2262.260 32.590 2262.320 ;
        RECT 15.710 2262.120 32.590 2262.260 ;
        RECT 15.710 2262.060 16.030 2262.120 ;
        RECT 32.270 2262.060 32.590 2262.120 ;
      LAYER via ;
        RECT 32.300 3202.840 32.560 3203.100 ;
        RECT 2260.080 3202.840 2260.340 3203.100 ;
        RECT 15.740 2262.060 16.000 2262.320 ;
        RECT 32.300 2262.060 32.560 2262.320 ;
      LAYER met2 ;
        RECT 32.300 3202.810 32.560 3203.130 ;
        RECT 2260.080 3202.810 2260.340 3203.130 ;
        RECT 32.360 2262.350 32.500 3202.810 ;
        RECT 2260.140 3200.000 2260.280 3202.810 ;
        RECT 2260.000 3197.600 2260.280 3200.000 ;
        RECT 15.740 2262.205 16.000 2262.350 ;
        RECT 15.730 2261.835 16.010 2262.205 ;
        RECT 32.300 2262.030 32.560 2262.350 ;
      LAYER via2 ;
        RECT 15.730 2261.880 16.010 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 15.705 2262.170 16.035 2262.185 ;
        RECT -4.800 2261.870 16.035 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 15.705 2261.855 16.035 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.710 3202.700 39.030 3202.760 ;
        RECT 2299.610 3202.700 2299.930 3202.760 ;
        RECT 38.710 3202.560 2299.930 3202.700 ;
        RECT 38.710 3202.500 39.030 3202.560 ;
        RECT 2299.610 3202.500 2299.930 3202.560 ;
        RECT 15.710 1977.340 16.030 1977.400 ;
        RECT 38.710 1977.340 39.030 1977.400 ;
        RECT 15.710 1977.200 39.030 1977.340 ;
        RECT 15.710 1977.140 16.030 1977.200 ;
        RECT 38.710 1977.140 39.030 1977.200 ;
      LAYER via ;
        RECT 38.740 3202.500 39.000 3202.760 ;
        RECT 2299.640 3202.500 2299.900 3202.760 ;
        RECT 15.740 1977.140 16.000 1977.400 ;
        RECT 38.740 1977.140 39.000 1977.400 ;
      LAYER met2 ;
        RECT 38.740 3202.470 39.000 3202.790 ;
        RECT 2299.640 3202.470 2299.900 3202.790 ;
        RECT 38.800 1977.430 38.940 3202.470 ;
        RECT 2299.700 3200.000 2299.840 3202.470 ;
        RECT 2299.560 3197.600 2299.840 3200.000 ;
        RECT 15.740 1977.110 16.000 1977.430 ;
        RECT 38.740 1977.110 39.000 1977.430 ;
        RECT 15.800 1975.245 15.940 1977.110 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 3205.420 1234.110 3205.480 ;
        RECT 2647.830 3205.420 2648.150 3205.480 ;
        RECT 1233.790 3205.280 2648.150 3205.420 ;
        RECT 1233.790 3205.220 1234.110 3205.280 ;
        RECT 2647.830 3205.220 2648.150 3205.280 ;
        RECT 2647.830 558.860 2648.150 558.920 ;
        RECT 2900.830 558.860 2901.150 558.920 ;
        RECT 2647.830 558.720 2901.150 558.860 ;
        RECT 2647.830 558.660 2648.150 558.720 ;
        RECT 2900.830 558.660 2901.150 558.720 ;
      LAYER via ;
        RECT 1233.820 3205.220 1234.080 3205.480 ;
        RECT 2647.860 3205.220 2648.120 3205.480 ;
        RECT 2647.860 558.660 2648.120 558.920 ;
        RECT 2900.860 558.660 2901.120 558.920 ;
      LAYER met2 ;
        RECT 1233.820 3205.190 1234.080 3205.510 ;
        RECT 2647.860 3205.190 2648.120 3205.510 ;
        RECT 1233.880 3200.000 1234.020 3205.190 ;
        RECT 1233.740 3197.600 1234.020 3200.000 ;
        RECT 2647.920 558.950 2648.060 3205.190 ;
        RECT 2647.860 558.630 2648.120 558.950 ;
        RECT 2900.860 558.630 2901.120 558.950 ;
        RECT 2900.920 557.445 2901.060 558.630 ;
        RECT 2900.850 557.075 2901.130 557.445 ;
      LAYER via2 ;
        RECT 2900.850 557.120 2901.130 557.400 ;
      LAYER met3 ;
        RECT 2900.825 557.410 2901.155 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2900.825 557.110 2924.800 557.410 ;
        RECT 2900.825 557.095 2901.155 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 31.810 3202.360 32.130 3202.420 ;
        RECT 2339.170 3202.360 2339.490 3202.420 ;
        RECT 31.810 3202.220 2339.490 3202.360 ;
        RECT 31.810 3202.160 32.130 3202.220 ;
        RECT 2339.170 3202.160 2339.490 3202.220 ;
        RECT 16.170 1689.700 16.490 1689.760 ;
        RECT 31.810 1689.700 32.130 1689.760 ;
        RECT 16.170 1689.560 32.130 1689.700 ;
        RECT 16.170 1689.500 16.490 1689.560 ;
        RECT 31.810 1689.500 32.130 1689.560 ;
      LAYER via ;
        RECT 31.840 3202.160 32.100 3202.420 ;
        RECT 2339.200 3202.160 2339.460 3202.420 ;
        RECT 16.200 1689.500 16.460 1689.760 ;
        RECT 31.840 1689.500 32.100 1689.760 ;
      LAYER met2 ;
        RECT 31.840 3202.130 32.100 3202.450 ;
        RECT 2339.200 3202.130 2339.460 3202.450 ;
        RECT 31.900 1689.790 32.040 3202.130 ;
        RECT 2339.260 3200.000 2339.400 3202.130 ;
        RECT 2339.120 3197.600 2339.400 3200.000 ;
        RECT 16.200 1689.470 16.460 1689.790 ;
        RECT 31.840 1689.470 32.100 1689.790 ;
        RECT 16.260 1687.605 16.400 1689.470 ;
        RECT 16.190 1687.235 16.470 1687.605 ;
      LAYER via2 ;
        RECT 16.190 1687.280 16.470 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 16.165 1687.570 16.495 1687.585 ;
        RECT -4.800 1687.270 16.495 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 16.165 1687.255 16.495 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 37.790 3202.020 38.110 3202.080 ;
        RECT 2378.730 3202.020 2379.050 3202.080 ;
        RECT 37.790 3201.880 2379.050 3202.020 ;
        RECT 37.790 3201.820 38.110 3201.880 ;
        RECT 2378.730 3201.820 2379.050 3201.880 ;
        RECT 16.630 1472.100 16.950 1472.160 ;
        RECT 37.790 1472.100 38.110 1472.160 ;
        RECT 16.630 1471.960 38.110 1472.100 ;
        RECT 16.630 1471.900 16.950 1471.960 ;
        RECT 37.790 1471.900 38.110 1471.960 ;
      LAYER via ;
        RECT 37.820 3201.820 38.080 3202.080 ;
        RECT 2378.760 3201.820 2379.020 3202.080 ;
        RECT 16.660 1471.900 16.920 1472.160 ;
        RECT 37.820 1471.900 38.080 1472.160 ;
      LAYER met2 ;
        RECT 37.820 3201.790 38.080 3202.110 ;
        RECT 2378.760 3201.790 2379.020 3202.110 ;
        RECT 37.880 1472.190 38.020 3201.790 ;
        RECT 2378.820 3200.000 2378.960 3201.790 ;
        RECT 2378.680 3197.600 2378.960 3200.000 ;
        RECT 16.660 1472.045 16.920 1472.190 ;
        RECT 16.650 1471.675 16.930 1472.045 ;
        RECT 37.820 1471.870 38.080 1472.190 ;
      LAYER via2 ;
        RECT 16.650 1471.720 16.930 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 16.625 1472.010 16.955 1472.025 ;
        RECT -4.800 1471.710 16.955 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 16.625 1471.695 16.955 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2418.310 3213.155 2418.590 3213.525 ;
        RECT 2418.380 3200.000 2418.520 3213.155 ;
        RECT 2418.240 3197.600 2418.520 3200.000 ;
        RECT 15.730 1262.235 16.010 1262.605 ;
        RECT 15.800 1256.485 15.940 1262.235 ;
        RECT 15.730 1256.115 16.010 1256.485 ;
      LAYER via2 ;
        RECT 2418.310 3213.200 2418.590 3213.480 ;
        RECT 15.730 1262.280 16.010 1262.560 ;
        RECT 15.730 1256.160 16.010 1256.440 ;
      LAYER met3 ;
        RECT 1164.070 3213.490 1164.450 3213.500 ;
        RECT 2418.285 3213.490 2418.615 3213.505 ;
        RECT 1164.070 3213.190 2418.615 3213.490 ;
        RECT 1164.070 3213.180 1164.450 3213.190 ;
        RECT 2418.285 3213.175 2418.615 3213.190 ;
        RECT 15.705 1262.570 16.035 1262.585 ;
        RECT 1164.070 1262.570 1164.450 1262.580 ;
        RECT 15.705 1262.270 1164.450 1262.570 ;
        RECT 15.705 1262.255 16.035 1262.270 ;
        RECT 1164.070 1262.260 1164.450 1262.270 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 15.705 1256.450 16.035 1256.465 ;
        RECT -4.800 1256.150 16.035 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 15.705 1256.135 16.035 1256.150 ;
      LAYER via3 ;
        RECT 1164.100 3213.180 1164.420 3213.500 ;
        RECT 1164.100 1262.260 1164.420 1262.580 ;
      LAYER met4 ;
        RECT 1164.095 3213.175 1164.425 3213.505 ;
        RECT 1164.110 1262.585 1164.410 3213.175 ;
        RECT 1164.095 1262.255 1164.425 1262.585 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2457.410 3212.475 2457.690 3212.845 ;
        RECT 2457.480 3200.000 2457.620 3212.475 ;
        RECT 2457.340 3197.600 2457.620 3200.000 ;
      LAYER via2 ;
        RECT 2457.410 3212.520 2457.690 3212.800 ;
      LAYER met3 ;
        RECT 1163.150 3212.810 1163.530 3212.820 ;
        RECT 2457.385 3212.810 2457.715 3212.825 ;
        RECT 1163.150 3212.510 2457.715 3212.810 ;
        RECT 1163.150 3212.500 1163.530 3212.510 ;
        RECT 2457.385 3212.495 2457.715 3212.510 ;
        RECT 1163.150 1041.570 1163.530 1041.580 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 3.070 1041.270 1163.530 1041.570 ;
        RECT 3.070 1040.890 3.370 1041.270 ;
        RECT 1163.150 1041.260 1163.530 1041.270 ;
        RECT -4.800 1040.590 3.370 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
      LAYER via3 ;
        RECT 1163.180 3212.500 1163.500 3212.820 ;
        RECT 1163.180 1041.260 1163.500 1041.580 ;
      LAYER met4 ;
        RECT 1163.175 3212.495 1163.505 3212.825 ;
        RECT 1163.190 1041.585 1163.490 3212.495 ;
        RECT 1163.175 1041.255 1163.505 1041.585 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2496.970 3211.795 2497.250 3212.165 ;
        RECT 2497.040 3200.000 2497.180 3211.795 ;
        RECT 2496.900 3197.600 2497.180 3200.000 ;
      LAYER via2 ;
        RECT 2496.970 3211.840 2497.250 3212.120 ;
      LAYER met3 ;
        RECT 1162.230 3212.130 1162.610 3212.140 ;
        RECT 2496.945 3212.130 2497.275 3212.145 ;
        RECT 1162.230 3211.830 2497.275 3212.130 ;
        RECT 1162.230 3211.820 1162.610 3211.830 ;
        RECT 2496.945 3211.815 2497.275 3211.830 ;
        RECT 1162.230 828.050 1162.610 828.060 ;
        RECT 3.070 827.750 1162.610 828.050 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 3.070 825.330 3.370 827.750 ;
        RECT 1162.230 827.740 1162.610 827.750 ;
        RECT -4.800 825.030 3.370 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
      LAYER via3 ;
        RECT 1162.260 3211.820 1162.580 3212.140 ;
        RECT 1162.260 827.740 1162.580 828.060 ;
      LAYER met4 ;
        RECT 1162.255 3211.815 1162.585 3212.145 ;
        RECT 1162.270 828.065 1162.570 3211.815 ;
        RECT 1162.255 827.735 1162.585 828.065 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2536.530 3210.435 2536.810 3210.805 ;
        RECT 2536.600 3200.000 2536.740 3210.435 ;
        RECT 2536.460 3197.600 2536.740 3200.000 ;
        RECT 18.950 3190.715 19.230 3191.085 ;
        RECT 19.020 610.485 19.160 3190.715 ;
        RECT 18.950 610.115 19.230 610.485 ;
      LAYER via2 ;
        RECT 2536.530 3210.480 2536.810 3210.760 ;
        RECT 18.950 3190.760 19.230 3191.040 ;
        RECT 18.950 610.160 19.230 610.440 ;
      LAYER met3 ;
        RECT 2172.390 3210.770 2172.770 3210.780 ;
        RECT 2536.505 3210.770 2536.835 3210.785 ;
        RECT 2172.390 3210.470 2536.835 3210.770 ;
        RECT 2172.390 3210.460 2172.770 3210.470 ;
        RECT 2536.505 3210.455 2536.835 3210.470 ;
        RECT 18.925 3191.050 19.255 3191.065 ;
        RECT 2172.390 3191.050 2172.770 3191.060 ;
        RECT 18.925 3190.750 2172.770 3191.050 ;
        RECT 18.925 3190.735 19.255 3190.750 ;
        RECT 2172.390 3190.740 2172.770 3190.750 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 18.925 610.450 19.255 610.465 ;
        RECT -4.800 610.150 19.255 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 18.925 610.135 19.255 610.150 ;
      LAYER via3 ;
        RECT 2172.420 3210.460 2172.740 3210.780 ;
        RECT 2172.420 3190.740 2172.740 3191.060 ;
      LAYER met4 ;
        RECT 2172.415 3210.455 2172.745 3210.785 ;
        RECT 2172.430 3191.065 2172.730 3210.455 ;
        RECT 2172.415 3190.735 2172.745 3191.065 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 3201.680 24.310 3201.740 ;
        RECT 2576.070 3201.680 2576.390 3201.740 ;
        RECT 23.990 3201.540 2576.390 3201.680 ;
        RECT 23.990 3201.480 24.310 3201.540 ;
        RECT 2576.070 3201.480 2576.390 3201.540 ;
        RECT 13.870 399.400 14.190 399.460 ;
        RECT 23.990 399.400 24.310 399.460 ;
        RECT 13.870 399.260 24.310 399.400 ;
        RECT 13.870 399.200 14.190 399.260 ;
        RECT 23.990 399.200 24.310 399.260 ;
      LAYER via ;
        RECT 24.020 3201.480 24.280 3201.740 ;
        RECT 2576.100 3201.480 2576.360 3201.740 ;
        RECT 13.900 399.200 14.160 399.460 ;
        RECT 24.020 399.200 24.280 399.460 ;
      LAYER met2 ;
        RECT 24.020 3201.450 24.280 3201.770 ;
        RECT 2576.100 3201.450 2576.360 3201.770 ;
        RECT 24.080 399.490 24.220 3201.450 ;
        RECT 2576.160 3200.000 2576.300 3201.450 ;
        RECT 2576.020 3197.600 2576.300 3200.000 ;
        RECT 13.900 399.170 14.160 399.490 ;
        RECT 24.020 399.170 24.280 399.490 ;
        RECT 13.960 394.925 14.100 399.170 ;
        RECT 13.890 394.555 14.170 394.925 ;
      LAYER via2 ;
        RECT 13.890 394.600 14.170 394.880 ;
      LAYER met3 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 13.865 394.890 14.195 394.905 ;
        RECT -4.800 394.590 14.195 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 13.865 394.575 14.195 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.050 3215.280 2145.370 3215.340 ;
        RECT 2615.630 3215.280 2615.950 3215.340 ;
        RECT 2145.050 3215.140 2615.950 3215.280 ;
        RECT 2145.050 3215.080 2145.370 3215.140 ;
        RECT 2615.630 3215.080 2615.950 3215.140 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 362.090 179.420 362.410 179.480 ;
        RECT 17.090 179.280 362.410 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 362.090 179.220 362.410 179.280 ;
      LAYER via ;
        RECT 2145.080 3215.080 2145.340 3215.340 ;
        RECT 2615.660 3215.080 2615.920 3215.340 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 362.120 179.220 362.380 179.480 ;
      LAYER met2 ;
        RECT 2145.080 3215.050 2145.340 3215.370 ;
        RECT 2615.660 3215.050 2615.920 3215.370 ;
        RECT 2145.140 3210.805 2145.280 3215.050 ;
        RECT 362.110 3210.435 362.390 3210.805 ;
        RECT 2145.070 3210.435 2145.350 3210.805 ;
        RECT 362.180 179.510 362.320 3210.435 ;
        RECT 2615.720 3200.000 2615.860 3215.050 ;
        RECT 2615.580 3197.600 2615.860 3200.000 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 362.120 179.190 362.380 179.510 ;
      LAYER via2 ;
        RECT 362.110 3210.480 362.390 3210.760 ;
        RECT 2145.070 3210.480 2145.350 3210.760 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 362.085 3210.770 362.415 3210.785 ;
        RECT 2145.045 3210.770 2145.375 3210.785 ;
        RECT 362.085 3210.470 2145.375 3210.770 ;
        RECT 362.085 3210.455 362.415 3210.470 ;
        RECT 2145.045 3210.455 2145.375 3210.470 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2648.290 793.460 2648.610 793.520 ;
        RECT 2898.530 793.460 2898.850 793.520 ;
        RECT 2648.290 793.320 2898.850 793.460 ;
        RECT 2648.290 793.260 2648.610 793.320 ;
        RECT 2898.530 793.260 2898.850 793.320 ;
      LAYER via ;
        RECT 2648.320 793.260 2648.580 793.520 ;
        RECT 2898.560 793.260 2898.820 793.520 ;
      LAYER met2 ;
        RECT 1273.300 3199.130 1273.580 3200.000 ;
        RECT 1274.750 3199.130 1275.030 3199.245 ;
        RECT 1273.300 3198.990 1275.030 3199.130 ;
        RECT 1273.300 3197.600 1273.580 3198.990 ;
        RECT 1274.750 3198.875 1275.030 3198.990 ;
        RECT 2648.310 3191.395 2648.590 3191.765 ;
        RECT 2648.380 793.550 2648.520 3191.395 ;
        RECT 2648.320 793.230 2648.580 793.550 ;
        RECT 2898.560 793.230 2898.820 793.550 ;
        RECT 2898.620 792.045 2898.760 793.230 ;
        RECT 2898.550 791.675 2898.830 792.045 ;
      LAYER via2 ;
        RECT 1274.750 3198.920 1275.030 3199.200 ;
        RECT 2648.310 3191.440 2648.590 3191.720 ;
        RECT 2898.550 791.720 2898.830 792.000 ;
      LAYER met3 ;
        RECT 1274.725 3199.210 1275.055 3199.225 ;
        RECT 1278.150 3199.210 1278.530 3199.220 ;
        RECT 1274.725 3198.910 1278.530 3199.210 ;
        RECT 1274.725 3198.895 1275.055 3198.910 ;
        RECT 1278.150 3198.900 1278.530 3198.910 ;
        RECT 1278.150 3191.730 1278.530 3191.740 ;
        RECT 2648.285 3191.730 2648.615 3191.745 ;
        RECT 1278.150 3191.430 2648.615 3191.730 ;
        RECT 1278.150 3191.420 1278.530 3191.430 ;
        RECT 2648.285 3191.415 2648.615 3191.430 ;
        RECT 2898.525 792.010 2898.855 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.525 791.710 2924.800 792.010 ;
        RECT 2898.525 791.695 2898.855 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
      LAYER via3 ;
        RECT 1278.180 3198.900 1278.500 3199.220 ;
        RECT 1278.180 3191.420 1278.500 3191.740 ;
      LAYER met4 ;
        RECT 1278.175 3198.895 1278.505 3199.225 ;
        RECT 1278.190 3191.745 1278.490 3198.895 ;
        RECT 1278.175 3191.415 1278.505 3191.745 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1312.910 3205.760 1313.230 3205.820 ;
        RECT 2652.890 3205.760 2653.210 3205.820 ;
        RECT 1312.910 3205.620 2653.210 3205.760 ;
        RECT 1312.910 3205.560 1313.230 3205.620 ;
        RECT 2652.890 3205.560 2653.210 3205.620 ;
        RECT 2652.890 1028.060 2653.210 1028.120 ;
        RECT 2900.830 1028.060 2901.150 1028.120 ;
        RECT 2652.890 1027.920 2901.150 1028.060 ;
        RECT 2652.890 1027.860 2653.210 1027.920 ;
        RECT 2900.830 1027.860 2901.150 1027.920 ;
      LAYER via ;
        RECT 1312.940 3205.560 1313.200 3205.820 ;
        RECT 2652.920 3205.560 2653.180 3205.820 ;
        RECT 2652.920 1027.860 2653.180 1028.120 ;
        RECT 2900.860 1027.860 2901.120 1028.120 ;
      LAYER met2 ;
        RECT 1312.940 3205.530 1313.200 3205.850 ;
        RECT 2652.920 3205.530 2653.180 3205.850 ;
        RECT 1313.000 3200.000 1313.140 3205.530 ;
        RECT 1312.860 3197.600 1313.140 3200.000 ;
        RECT 2652.980 1028.150 2653.120 3205.530 ;
        RECT 2652.920 1027.830 2653.180 1028.150 ;
        RECT 2900.860 1027.830 2901.120 1028.150 ;
        RECT 2900.920 1026.645 2901.060 1027.830 ;
        RECT 2900.850 1026.275 2901.130 1026.645 ;
      LAYER via2 ;
        RECT 2900.850 1026.320 2901.130 1026.600 ;
      LAYER met3 ;
        RECT 2900.825 1026.610 2901.155 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2900.825 1026.310 2924.800 1026.610 ;
        RECT 2900.825 1026.295 2901.155 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.470 3212.560 1352.790 3212.620 ;
        RECT 2653.350 3212.560 2653.670 3212.620 ;
        RECT 1352.470 3212.420 2653.670 3212.560 ;
        RECT 1352.470 3212.360 1352.790 3212.420 ;
        RECT 2653.350 3212.360 2653.670 3212.420 ;
        RECT 2653.350 1262.660 2653.670 1262.720 ;
        RECT 2898.070 1262.660 2898.390 1262.720 ;
        RECT 2653.350 1262.520 2898.390 1262.660 ;
        RECT 2653.350 1262.460 2653.670 1262.520 ;
        RECT 2898.070 1262.460 2898.390 1262.520 ;
      LAYER via ;
        RECT 1352.500 3212.360 1352.760 3212.620 ;
        RECT 2653.380 3212.360 2653.640 3212.620 ;
        RECT 2653.380 1262.460 2653.640 1262.720 ;
        RECT 2898.100 1262.460 2898.360 1262.720 ;
      LAYER met2 ;
        RECT 1352.500 3212.330 1352.760 3212.650 ;
        RECT 2653.380 3212.330 2653.640 3212.650 ;
        RECT 1352.560 3200.000 1352.700 3212.330 ;
        RECT 1352.420 3197.600 1352.700 3200.000 ;
        RECT 2653.440 1262.750 2653.580 3212.330 ;
        RECT 2653.380 1262.430 2653.640 1262.750 ;
        RECT 2898.100 1262.430 2898.360 1262.750 ;
        RECT 2898.160 1261.245 2898.300 1262.430 ;
        RECT 2898.090 1260.875 2898.370 1261.245 ;
      LAYER via2 ;
        RECT 2898.090 1260.920 2898.370 1261.200 ;
      LAYER met3 ;
        RECT 2898.065 1261.210 2898.395 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.065 1260.910 2924.800 1261.210 ;
        RECT 2898.065 1260.895 2898.395 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1391.570 3212.220 1391.890 3212.280 ;
        RECT 2904.510 3212.220 2904.830 3212.280 ;
        RECT 1391.570 3212.080 2904.830 3212.220 ;
        RECT 1391.570 3212.020 1391.890 3212.080 ;
        RECT 2904.510 3212.020 2904.830 3212.080 ;
      LAYER via ;
        RECT 1391.600 3212.020 1391.860 3212.280 ;
        RECT 2904.540 3212.020 2904.800 3212.280 ;
      LAYER met2 ;
        RECT 1391.600 3211.990 1391.860 3212.310 ;
        RECT 2904.540 3211.990 2904.800 3212.310 ;
        RECT 1391.660 3200.000 1391.800 3211.990 ;
        RECT 1391.520 3197.600 1391.800 3200.000 ;
        RECT 2904.600 1495.845 2904.740 3211.990 ;
        RECT 2904.530 1495.475 2904.810 1495.845 ;
      LAYER via2 ;
        RECT 2904.530 1495.520 2904.810 1495.800 ;
      LAYER met3 ;
        RECT 2904.505 1495.810 2904.835 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2904.505 1495.510 2924.800 1495.810 ;
        RECT 2904.505 1495.495 2904.835 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1431.130 3206.440 1431.450 3206.500 ;
        RECT 2654.730 3206.440 2655.050 3206.500 ;
        RECT 1431.130 3206.300 2655.050 3206.440 ;
        RECT 1431.130 3206.240 1431.450 3206.300 ;
        RECT 2654.730 3206.240 2655.050 3206.300 ;
        RECT 2654.730 1731.860 2655.050 1731.920 ;
        RECT 2898.990 1731.860 2899.310 1731.920 ;
        RECT 2654.730 1731.720 2899.310 1731.860 ;
        RECT 2654.730 1731.660 2655.050 1731.720 ;
        RECT 2898.990 1731.660 2899.310 1731.720 ;
      LAYER via ;
        RECT 1431.160 3206.240 1431.420 3206.500 ;
        RECT 2654.760 3206.240 2655.020 3206.500 ;
        RECT 2654.760 1731.660 2655.020 1731.920 ;
        RECT 2899.020 1731.660 2899.280 1731.920 ;
      LAYER met2 ;
        RECT 1431.160 3206.210 1431.420 3206.530 ;
        RECT 2654.760 3206.210 2655.020 3206.530 ;
        RECT 1431.220 3200.000 1431.360 3206.210 ;
        RECT 1431.080 3197.600 1431.360 3200.000 ;
        RECT 2654.820 1731.950 2654.960 3206.210 ;
        RECT 2654.760 1731.630 2655.020 1731.950 ;
        RECT 2899.020 1731.630 2899.280 1731.950 ;
        RECT 2899.080 1730.445 2899.220 1731.630 ;
        RECT 2899.010 1730.075 2899.290 1730.445 ;
      LAYER via2 ;
        RECT 2899.010 1730.120 2899.290 1730.400 ;
      LAYER met3 ;
        RECT 2898.985 1730.410 2899.315 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2898.985 1730.110 2924.800 1730.410 ;
        RECT 2898.985 1730.095 2899.315 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1470.690 3212.900 1471.010 3212.960 ;
        RECT 2655.190 3212.900 2655.510 3212.960 ;
        RECT 1470.690 3212.760 2655.510 3212.900 ;
        RECT 1470.690 3212.700 1471.010 3212.760 ;
        RECT 2655.190 3212.700 2655.510 3212.760 ;
        RECT 2655.190 1966.460 2655.510 1966.520 ;
        RECT 2899.450 1966.460 2899.770 1966.520 ;
        RECT 2655.190 1966.320 2899.770 1966.460 ;
        RECT 2655.190 1966.260 2655.510 1966.320 ;
        RECT 2899.450 1966.260 2899.770 1966.320 ;
      LAYER via ;
        RECT 1470.720 3212.700 1470.980 3212.960 ;
        RECT 2655.220 3212.700 2655.480 3212.960 ;
        RECT 2655.220 1966.260 2655.480 1966.520 ;
        RECT 2899.480 1966.260 2899.740 1966.520 ;
      LAYER met2 ;
        RECT 1470.720 3212.670 1470.980 3212.990 ;
        RECT 2655.220 3212.670 2655.480 3212.990 ;
        RECT 1470.780 3200.000 1470.920 3212.670 ;
        RECT 1470.640 3197.600 1470.920 3200.000 ;
        RECT 2655.280 1966.550 2655.420 3212.670 ;
        RECT 2655.220 1966.230 2655.480 1966.550 ;
        RECT 2899.480 1966.230 2899.740 1966.550 ;
        RECT 2899.540 1965.045 2899.680 1966.230 ;
        RECT 2899.470 1964.675 2899.750 1965.045 ;
      LAYER via2 ;
        RECT 2899.470 1964.720 2899.750 1965.000 ;
      LAYER met3 ;
        RECT 2899.445 1965.010 2899.775 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2899.445 1964.710 2924.800 1965.010 ;
        RECT 2899.445 1964.695 2899.775 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2656.110 2201.060 2656.430 2201.120 ;
        RECT 2899.450 2201.060 2899.770 2201.120 ;
        RECT 2656.110 2200.920 2899.770 2201.060 ;
        RECT 2656.110 2200.860 2656.430 2200.920 ;
        RECT 2899.450 2200.860 2899.770 2200.920 ;
      LAYER via ;
        RECT 2656.140 2200.860 2656.400 2201.120 ;
        RECT 2899.480 2200.860 2899.740 2201.120 ;
      LAYER met2 ;
        RECT 1510.270 3200.235 1510.550 3200.605 ;
        RECT 1510.340 3200.000 1510.480 3200.235 ;
        RECT 1510.200 3197.600 1510.480 3200.000 ;
        RECT 2656.130 3192.075 2656.410 3192.445 ;
        RECT 2656.200 2201.150 2656.340 3192.075 ;
        RECT 2656.140 2200.830 2656.400 2201.150 ;
        RECT 2899.480 2200.830 2899.740 2201.150 ;
        RECT 2899.540 2199.645 2899.680 2200.830 ;
        RECT 2899.470 2199.275 2899.750 2199.645 ;
      LAYER via2 ;
        RECT 1510.270 3200.280 1510.550 3200.560 ;
        RECT 2656.130 3192.120 2656.410 3192.400 ;
        RECT 2899.470 2199.320 2899.750 2199.600 ;
      LAYER met3 ;
        RECT 1510.245 3200.580 1510.575 3200.585 ;
        RECT 1509.990 3200.570 1510.575 3200.580 ;
        RECT 1509.790 3200.270 1510.575 3200.570 ;
        RECT 1509.990 3200.260 1510.575 3200.270 ;
        RECT 1510.245 3200.255 1510.575 3200.260 ;
        RECT 1509.990 3192.410 1510.370 3192.420 ;
        RECT 2656.105 3192.410 2656.435 3192.425 ;
        RECT 1509.990 3192.110 2656.435 3192.410 ;
        RECT 1509.990 3192.100 1510.370 3192.110 ;
        RECT 2656.105 3192.095 2656.435 3192.110 ;
        RECT 2899.445 2199.610 2899.775 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2899.445 2199.310 2924.800 2199.610 ;
        RECT 2899.445 2199.295 2899.775 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
      LAYER via3 ;
        RECT 1510.020 3200.260 1510.340 3200.580 ;
        RECT 1510.020 3192.100 1510.340 3192.420 ;
      LAYER met4 ;
        RECT 1510.015 3200.255 1510.345 3200.585 ;
        RECT 1510.030 3192.425 1510.330 3200.255 ;
        RECT 1510.015 3192.095 1510.345 3192.425 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1988.190 201.860 1988.510 201.920 ;
        RECT 2028.210 201.860 2028.530 201.920 ;
        RECT 1988.190 201.720 2028.530 201.860 ;
        RECT 1988.190 201.660 1988.510 201.720 ;
        RECT 2028.210 201.660 2028.530 201.720 ;
        RECT 2379.650 201.180 2379.970 201.240 ;
        RECT 2391.150 201.180 2391.470 201.240 ;
        RECT 2379.650 201.040 2391.470 201.180 ;
        RECT 2379.650 200.980 2379.970 201.040 ;
        RECT 2391.150 200.980 2391.470 201.040 ;
        RECT 2572.850 201.180 2573.170 201.240 ;
        RECT 2574.230 201.180 2574.550 201.240 ;
        RECT 2572.850 201.040 2574.550 201.180 ;
        RECT 2572.850 200.980 2573.170 201.040 ;
        RECT 2574.230 200.980 2574.550 201.040 ;
        RECT 2704.870 200.500 2705.190 200.560 ;
        RECT 2729.250 200.500 2729.570 200.560 ;
        RECT 2704.870 200.360 2729.570 200.500 ;
        RECT 2704.870 200.300 2705.190 200.360 ;
        RECT 2729.250 200.300 2729.570 200.360 ;
        RECT 1510.710 200.160 1511.030 200.220 ;
        RECT 1536.470 200.160 1536.790 200.220 ;
        RECT 1510.710 200.020 1536.790 200.160 ;
        RECT 1510.710 199.960 1511.030 200.020 ;
        RECT 1536.470 199.960 1536.790 200.020 ;
      LAYER via ;
        RECT 1988.220 201.660 1988.480 201.920 ;
        RECT 2028.240 201.660 2028.500 201.920 ;
        RECT 2379.680 200.980 2379.940 201.240 ;
        RECT 2391.180 200.980 2391.440 201.240 ;
        RECT 2572.880 200.980 2573.140 201.240 ;
        RECT 2574.260 200.980 2574.520 201.240 ;
        RECT 2704.900 200.300 2705.160 200.560 ;
        RECT 2729.280 200.300 2729.540 200.560 ;
        RECT 1510.740 199.960 1511.000 200.220 ;
        RECT 1536.500 199.960 1536.760 200.220 ;
      LAYER met2 ;
        RECT 1167.960 3199.130 1168.240 3200.000 ;
        RECT 1169.870 3199.130 1170.150 3199.245 ;
        RECT 1167.960 3198.990 1170.150 3199.130 ;
        RECT 1167.960 3197.600 1168.240 3198.990 ;
        RECT 1169.870 3198.875 1170.150 3198.990 ;
        RECT 1869.530 202.795 1869.810 203.165 ;
        RECT 1821.230 202.115 1821.510 202.485 ;
        RECT 1365.370 201.690 1365.650 201.805 ;
        RECT 1366.290 201.690 1366.570 201.805 ;
        RECT 1365.370 201.550 1366.570 201.690 ;
        RECT 1365.370 201.435 1365.650 201.550 ;
        RECT 1366.290 201.435 1366.570 201.550 ;
        RECT 1724.630 201.435 1724.910 201.805 ;
        RECT 1449.090 200.755 1449.370 201.125 ;
        RECT 1536.490 200.755 1536.770 201.125 ;
        RECT 1676.330 200.755 1676.610 201.125 ;
        RECT 1449.160 200.445 1449.300 200.755 ;
        RECT 1449.090 200.075 1449.370 200.445 ;
        RECT 1510.730 200.075 1511.010 200.445 ;
        RECT 1536.560 200.250 1536.700 200.755 ;
        RECT 1676.400 200.445 1676.540 200.755 ;
        RECT 1724.700 200.445 1724.840 201.435 ;
        RECT 1821.300 201.125 1821.440 202.115 ;
        RECT 1869.600 201.125 1869.740 202.795 ;
        RECT 1988.220 201.805 1988.480 201.950 ;
        RECT 2028.240 201.805 2028.500 201.950 ;
        RECT 1988.210 201.435 1988.490 201.805 ;
        RECT 2028.230 201.435 2028.510 201.805 ;
        RECT 2090.330 201.435 2090.610 201.805 ;
        RECT 2283.990 201.435 2284.270 201.805 ;
        RECT 2772.510 201.435 2772.790 201.805 ;
        RECT 1821.230 200.755 1821.510 201.125 ;
        RECT 1869.530 200.755 1869.810 201.125 ;
        RECT 2090.400 201.010 2090.540 201.435 ;
        RECT 2090.790 201.010 2091.070 201.125 ;
        RECT 2090.400 200.870 2091.070 201.010 ;
        RECT 2090.790 200.755 2091.070 200.870 ;
        RECT 2283.530 201.010 2283.810 201.125 ;
        RECT 2284.060 201.010 2284.200 201.435 ;
        RECT 2379.680 201.125 2379.940 201.270 ;
        RECT 2391.180 201.125 2391.440 201.270 ;
        RECT 2572.880 201.125 2573.140 201.270 ;
        RECT 2574.260 201.125 2574.520 201.270 ;
        RECT 2283.530 200.870 2284.200 201.010 ;
        RECT 2283.530 200.755 2283.810 200.870 ;
        RECT 2379.670 200.755 2379.950 201.125 ;
        RECT 2391.170 200.755 2391.450 201.125 ;
        RECT 2572.870 200.755 2573.150 201.125 ;
        RECT 2574.250 200.755 2574.530 201.125 ;
        RECT 2729.270 200.755 2729.550 201.125 ;
        RECT 2729.340 200.590 2729.480 200.755 ;
        RECT 2704.900 200.445 2705.160 200.590 ;
        RECT 1510.740 199.930 1511.000 200.075 ;
        RECT 1536.500 199.930 1536.760 200.250 ;
        RECT 1676.330 200.075 1676.610 200.445 ;
        RECT 1724.630 200.075 1724.910 200.445 ;
        RECT 2704.890 200.075 2705.170 200.445 ;
        RECT 2729.280 200.270 2729.540 200.590 ;
        RECT 2772.580 199.765 2772.720 201.435 ;
        RECT 2863.130 200.755 2863.410 201.125 ;
        RECT 2863.200 200.330 2863.340 200.755 ;
        RECT 2863.590 200.330 2863.870 200.445 ;
        RECT 2863.200 200.190 2863.870 200.330 ;
        RECT 2863.590 200.075 2863.870 200.190 ;
        RECT 2772.510 199.395 2772.790 199.765 ;
      LAYER via2 ;
        RECT 1169.870 3198.920 1170.150 3199.200 ;
        RECT 1869.530 202.840 1869.810 203.120 ;
        RECT 1821.230 202.160 1821.510 202.440 ;
        RECT 1365.370 201.480 1365.650 201.760 ;
        RECT 1366.290 201.480 1366.570 201.760 ;
        RECT 1724.630 201.480 1724.910 201.760 ;
        RECT 1449.090 200.800 1449.370 201.080 ;
        RECT 1536.490 200.800 1536.770 201.080 ;
        RECT 1676.330 200.800 1676.610 201.080 ;
        RECT 1449.090 200.120 1449.370 200.400 ;
        RECT 1510.730 200.120 1511.010 200.400 ;
        RECT 1988.210 201.480 1988.490 201.760 ;
        RECT 2028.230 201.480 2028.510 201.760 ;
        RECT 2090.330 201.480 2090.610 201.760 ;
        RECT 2283.990 201.480 2284.270 201.760 ;
        RECT 2772.510 201.480 2772.790 201.760 ;
        RECT 1821.230 200.800 1821.510 201.080 ;
        RECT 1869.530 200.800 1869.810 201.080 ;
        RECT 2090.790 200.800 2091.070 201.080 ;
        RECT 2283.530 200.800 2283.810 201.080 ;
        RECT 2379.670 200.800 2379.950 201.080 ;
        RECT 2391.170 200.800 2391.450 201.080 ;
        RECT 2572.870 200.800 2573.150 201.080 ;
        RECT 2574.250 200.800 2574.530 201.080 ;
        RECT 2729.270 200.800 2729.550 201.080 ;
        RECT 1676.330 200.120 1676.610 200.400 ;
        RECT 1724.630 200.120 1724.910 200.400 ;
        RECT 2704.890 200.120 2705.170 200.400 ;
        RECT 2863.130 200.800 2863.410 201.080 ;
        RECT 2863.590 200.120 2863.870 200.400 ;
        RECT 2772.510 199.440 2772.790 199.720 ;
      LAYER met3 ;
        RECT 1169.845 3199.210 1170.175 3199.225 ;
        RECT 1172.350 3199.210 1172.730 3199.220 ;
        RECT 1169.845 3198.910 1172.730 3199.210 ;
        RECT 1169.845 3198.895 1170.175 3198.910 ;
        RECT 1172.350 3198.900 1172.730 3198.910 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 1869.505 203.140 1869.835 203.145 ;
        RECT 1869.505 203.130 1870.090 203.140 ;
        RECT 1869.505 202.830 1870.470 203.130 ;
        RECT 1869.505 202.820 1870.090 202.830 ;
        RECT 1869.505 202.815 1869.835 202.820 ;
        RECT 1773.110 202.450 1773.490 202.460 ;
        RECT 1821.205 202.450 1821.535 202.465 ;
        RECT 1268.990 202.150 1270.210 202.450 ;
        RECT 1268.990 201.090 1269.290 202.150 ;
        RECT 1269.910 201.770 1270.210 202.150 ;
        RECT 1773.110 202.150 1821.535 202.450 ;
        RECT 1773.110 202.140 1773.490 202.150 ;
        RECT 1821.205 202.135 1821.535 202.150 ;
        RECT 2463.150 202.150 2511.290 202.450 ;
        RECT 1365.345 201.770 1365.675 201.785 ;
        RECT 1269.910 201.470 1365.675 201.770 ;
        RECT 1365.345 201.455 1365.675 201.470 ;
        RECT 1366.265 201.770 1366.595 201.785 ;
        RECT 1676.510 201.770 1676.890 201.780 ;
        RECT 1724.605 201.770 1724.935 201.785 ;
        RECT 1366.265 201.470 1424.770 201.770 ;
        RECT 1366.265 201.455 1366.595 201.470 ;
        RECT 1173.310 200.790 1269.290 201.090 ;
        RECT 1424.470 201.090 1424.770 201.470 ;
        RECT 1676.510 201.470 1724.935 201.770 ;
        RECT 1676.510 201.460 1676.890 201.470 ;
        RECT 1724.605 201.455 1724.935 201.470 ;
        RECT 1869.710 201.770 1870.090 201.780 ;
        RECT 1988.185 201.770 1988.515 201.785 ;
        RECT 1869.710 201.470 1870.970 201.770 ;
        RECT 1869.710 201.460 1870.090 201.470 ;
        RECT 1449.065 201.090 1449.395 201.105 ;
        RECT 1424.470 200.790 1449.395 201.090 ;
        RECT 1172.350 200.410 1172.730 200.420 ;
        RECT 1173.310 200.410 1173.610 200.790 ;
        RECT 1449.065 200.775 1449.395 200.790 ;
        RECT 1536.465 201.090 1536.795 201.105 ;
        RECT 1676.305 201.090 1676.635 201.105 ;
        RECT 1773.110 201.090 1773.490 201.100 ;
        RECT 1536.465 200.790 1676.635 201.090 ;
        RECT 1536.465 200.775 1536.795 200.790 ;
        RECT 1676.305 200.775 1676.635 200.790 ;
        RECT 1725.310 200.790 1773.490 201.090 ;
        RECT 1172.350 200.110 1173.610 200.410 ;
        RECT 1449.065 200.410 1449.395 200.425 ;
        RECT 1510.705 200.410 1511.035 200.425 ;
        RECT 1449.065 200.110 1511.035 200.410 ;
        RECT 1172.350 200.100 1172.730 200.110 ;
        RECT 1449.065 200.095 1449.395 200.110 ;
        RECT 1510.705 200.095 1511.035 200.110 ;
        RECT 1676.305 200.420 1676.635 200.425 ;
        RECT 1676.305 200.410 1676.890 200.420 ;
        RECT 1724.605 200.410 1724.935 200.425 ;
        RECT 1725.310 200.410 1725.610 200.790 ;
        RECT 1773.110 200.780 1773.490 200.790 ;
        RECT 1821.205 201.090 1821.535 201.105 ;
        RECT 1869.505 201.090 1869.835 201.105 ;
        RECT 1821.205 200.790 1869.835 201.090 ;
        RECT 1870.670 201.090 1870.970 201.470 ;
        RECT 1946.110 201.470 1988.515 201.770 ;
        RECT 1946.110 201.090 1946.410 201.470 ;
        RECT 1988.185 201.455 1988.515 201.470 ;
        RECT 2028.205 201.770 2028.535 201.785 ;
        RECT 2090.305 201.770 2090.635 201.785 ;
        RECT 2283.965 201.770 2284.295 201.785 ;
        RECT 2028.205 201.470 2042.090 201.770 ;
        RECT 2028.205 201.455 2028.535 201.470 ;
        RECT 1870.670 200.790 1946.410 201.090 ;
        RECT 1821.205 200.775 1821.535 200.790 ;
        RECT 1869.505 200.775 1869.835 200.790 ;
        RECT 1676.305 200.110 1677.270 200.410 ;
        RECT 1724.605 200.110 1725.610 200.410 ;
        RECT 2041.790 200.410 2042.090 201.470 ;
        RECT 2076.750 201.470 2090.635 201.770 ;
        RECT 2076.750 201.090 2077.050 201.470 ;
        RECT 2090.305 201.455 2090.635 201.470 ;
        RECT 2124.590 201.470 2138.690 201.770 ;
        RECT 2042.710 200.790 2077.050 201.090 ;
        RECT 2090.765 201.090 2091.095 201.105 ;
        RECT 2124.590 201.090 2124.890 201.470 ;
        RECT 2090.765 200.790 2124.890 201.090 ;
        RECT 2042.710 200.410 2043.010 200.790 ;
        RECT 2090.765 200.775 2091.095 200.790 ;
        RECT 2041.790 200.110 2043.010 200.410 ;
        RECT 2138.390 200.410 2138.690 201.470 ;
        RECT 2139.310 201.470 2187.450 201.770 ;
        RECT 2139.310 200.410 2139.610 201.470 ;
        RECT 2138.390 200.110 2139.610 200.410 ;
        RECT 2187.150 200.410 2187.450 201.470 ;
        RECT 2283.965 201.470 2284.970 201.770 ;
        RECT 2283.965 201.455 2284.295 201.470 ;
        RECT 2283.505 201.090 2283.835 201.105 ;
        RECT 2235.910 200.790 2283.835 201.090 ;
        RECT 2284.670 201.090 2284.970 201.470 ;
        RECT 2379.645 201.090 2379.975 201.105 ;
        RECT 2284.670 200.790 2331.890 201.090 ;
        RECT 2235.910 200.410 2236.210 200.790 ;
        RECT 2283.505 200.775 2283.835 200.790 ;
        RECT 2187.150 200.110 2236.210 200.410 ;
        RECT 2331.590 200.410 2331.890 200.790 ;
        RECT 2332.510 200.790 2379.975 201.090 ;
        RECT 2332.510 200.410 2332.810 200.790 ;
        RECT 2379.645 200.775 2379.975 200.790 ;
        RECT 2391.145 201.090 2391.475 201.105 ;
        RECT 2463.150 201.090 2463.450 202.150 ;
        RECT 2510.990 201.780 2511.290 202.150 ;
        RECT 2510.950 201.460 2511.330 201.780 ;
        RECT 2772.485 201.770 2772.815 201.785 ;
        RECT 2772.485 201.470 2815.810 201.770 ;
        RECT 2772.485 201.455 2772.815 201.470 ;
        RECT 2572.845 201.090 2573.175 201.105 ;
        RECT 2391.145 200.790 2414.690 201.090 ;
        RECT 2391.145 200.775 2391.475 200.790 ;
        RECT 2331.590 200.110 2332.810 200.410 ;
        RECT 2414.390 200.410 2414.690 200.790 ;
        RECT 2429.110 200.790 2463.450 201.090 ;
        RECT 2525.710 200.790 2573.175 201.090 ;
        RECT 2429.110 200.410 2429.410 200.790 ;
        RECT 2414.390 200.110 2429.410 200.410 ;
        RECT 2510.950 200.410 2511.330 200.420 ;
        RECT 2525.710 200.410 2526.010 200.790 ;
        RECT 2572.845 200.775 2573.175 200.790 ;
        RECT 2574.225 201.090 2574.555 201.105 ;
        RECT 2656.310 201.090 2656.690 201.100 ;
        RECT 2574.225 200.790 2621.690 201.090 ;
        RECT 2574.225 200.775 2574.555 200.790 ;
        RECT 2510.950 200.110 2526.010 200.410 ;
        RECT 2621.390 200.410 2621.690 200.790 ;
        RECT 2622.310 200.790 2656.690 201.090 ;
        RECT 2622.310 200.410 2622.610 200.790 ;
        RECT 2656.310 200.780 2656.690 200.790 ;
        RECT 2729.245 201.090 2729.575 201.105 ;
        RECT 2752.910 201.090 2753.290 201.100 ;
        RECT 2729.245 200.790 2753.290 201.090 ;
        RECT 2729.245 200.775 2729.575 200.790 ;
        RECT 2752.910 200.780 2753.290 200.790 ;
        RECT 2704.865 200.410 2705.195 200.425 ;
        RECT 2621.390 200.110 2622.610 200.410 ;
        RECT 2704.190 200.110 2705.195 200.410 ;
        RECT 2815.510 200.410 2815.810 201.470 ;
        RECT 2863.105 201.090 2863.435 201.105 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2849.550 200.790 2863.435 201.090 ;
        RECT 2849.550 200.410 2849.850 200.790 ;
        RECT 2863.105 200.775 2863.435 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2815.510 200.110 2849.850 200.410 ;
        RECT 2863.565 200.410 2863.895 200.425 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2863.565 200.110 2884.810 200.410 ;
        RECT 1676.305 200.100 1676.890 200.110 ;
        RECT 1676.305 200.095 1676.635 200.100 ;
        RECT 1724.605 200.095 1724.935 200.110 ;
        RECT 2510.950 200.100 2511.330 200.110 ;
        RECT 2656.310 199.050 2656.690 199.060 ;
        RECT 2704.190 199.050 2704.490 200.110 ;
        RECT 2704.865 200.095 2705.195 200.110 ;
        RECT 2863.565 200.095 2863.895 200.110 ;
        RECT 2752.910 199.730 2753.290 199.740 ;
        RECT 2772.485 199.730 2772.815 199.745 ;
        RECT 2752.910 199.430 2772.815 199.730 ;
        RECT 2752.910 199.420 2753.290 199.430 ;
        RECT 2772.485 199.415 2772.815 199.430 ;
        RECT 2656.310 198.750 2704.490 199.050 ;
        RECT 2656.310 198.740 2656.690 198.750 ;
      LAYER via3 ;
        RECT 1172.380 3198.900 1172.700 3199.220 ;
        RECT 1869.740 202.820 1870.060 203.140 ;
        RECT 1773.140 202.140 1773.460 202.460 ;
        RECT 1676.540 201.460 1676.860 201.780 ;
        RECT 1869.740 201.460 1870.060 201.780 ;
        RECT 1172.380 200.100 1172.700 200.420 ;
        RECT 1676.540 200.100 1676.860 200.420 ;
        RECT 1773.140 200.780 1773.460 201.100 ;
        RECT 2510.980 201.460 2511.300 201.780 ;
        RECT 2510.980 200.100 2511.300 200.420 ;
        RECT 2656.340 200.780 2656.660 201.100 ;
        RECT 2752.940 200.780 2753.260 201.100 ;
        RECT 2656.340 198.740 2656.660 199.060 ;
        RECT 2752.940 199.420 2753.260 199.740 ;
      LAYER met4 ;
        RECT 1172.375 3198.895 1172.705 3199.225 ;
        RECT 1172.390 200.425 1172.690 3198.895 ;
        RECT 1869.735 202.815 1870.065 203.145 ;
        RECT 1773.135 202.135 1773.465 202.465 ;
        RECT 1676.535 201.455 1676.865 201.785 ;
        RECT 1676.550 200.425 1676.850 201.455 ;
        RECT 1773.150 201.105 1773.450 202.135 ;
        RECT 1869.750 201.785 1870.050 202.815 ;
        RECT 1869.735 201.455 1870.065 201.785 ;
        RECT 2510.975 201.455 2511.305 201.785 ;
        RECT 1773.135 200.775 1773.465 201.105 ;
        RECT 2510.990 200.425 2511.290 201.455 ;
        RECT 2656.335 200.775 2656.665 201.105 ;
        RECT 2752.935 200.775 2753.265 201.105 ;
        RECT 1172.375 200.095 1172.705 200.425 ;
        RECT 1676.535 200.095 1676.865 200.425 ;
        RECT 2510.975 200.095 2511.305 200.425 ;
        RECT 2656.350 199.065 2656.650 200.775 ;
        RECT 2752.950 199.745 2753.250 200.775 ;
        RECT 2752.935 199.415 2753.265 199.745 ;
        RECT 2656.335 198.735 2656.665 199.065 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1562.690 3207.460 1563.010 3207.520 ;
        RECT 2652.430 3207.460 2652.750 3207.520 ;
        RECT 1562.690 3207.320 2652.750 3207.460 ;
        RECT 1562.690 3207.260 1563.010 3207.320 ;
        RECT 2652.430 3207.260 2652.750 3207.320 ;
        RECT 2652.430 2552.960 2652.750 2553.020 ;
        RECT 2898.990 2552.960 2899.310 2553.020 ;
        RECT 2652.430 2552.820 2899.310 2552.960 ;
        RECT 2652.430 2552.760 2652.750 2552.820 ;
        RECT 2898.990 2552.760 2899.310 2552.820 ;
      LAYER via ;
        RECT 1562.720 3207.260 1562.980 3207.520 ;
        RECT 2652.460 3207.260 2652.720 3207.520 ;
        RECT 2652.460 2552.760 2652.720 2553.020 ;
        RECT 2899.020 2552.760 2899.280 2553.020 ;
      LAYER met2 ;
        RECT 1562.720 3207.230 1562.980 3207.550 ;
        RECT 2652.460 3207.230 2652.720 3207.550 ;
        RECT 1562.780 3200.000 1562.920 3207.230 ;
        RECT 1562.640 3197.600 1562.920 3200.000 ;
        RECT 2652.520 2553.050 2652.660 3207.230 ;
        RECT 2652.460 2552.730 2652.720 2553.050 ;
        RECT 2899.020 2552.730 2899.280 2553.050 ;
        RECT 2899.080 2551.885 2899.220 2552.730 ;
        RECT 2899.010 2551.515 2899.290 2551.885 ;
      LAYER via2 ;
        RECT 2899.010 2551.560 2899.290 2551.840 ;
      LAYER met3 ;
        RECT 2898.985 2551.850 2899.315 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2898.985 2551.550 2924.800 2551.850 ;
        RECT 2898.985 2551.535 2899.315 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1602.250 3213.920 1602.570 3213.980 ;
        RECT 2651.970 3213.920 2652.290 3213.980 ;
        RECT 1602.250 3213.780 2652.290 3213.920 ;
        RECT 1602.250 3213.720 1602.570 3213.780 ;
        RECT 2651.970 3213.720 2652.290 3213.780 ;
        RECT 2651.970 2787.560 2652.290 2787.620 ;
        RECT 2898.990 2787.560 2899.310 2787.620 ;
        RECT 2651.970 2787.420 2899.310 2787.560 ;
        RECT 2651.970 2787.360 2652.290 2787.420 ;
        RECT 2898.990 2787.360 2899.310 2787.420 ;
      LAYER via ;
        RECT 1602.280 3213.720 1602.540 3213.980 ;
        RECT 2652.000 3213.720 2652.260 3213.980 ;
        RECT 2652.000 2787.360 2652.260 2787.620 ;
        RECT 2899.020 2787.360 2899.280 2787.620 ;
      LAYER met2 ;
        RECT 1602.280 3213.690 1602.540 3214.010 ;
        RECT 2652.000 3213.690 2652.260 3214.010 ;
        RECT 1602.340 3200.000 1602.480 3213.690 ;
        RECT 1602.200 3197.600 1602.480 3200.000 ;
        RECT 2652.060 2787.650 2652.200 3213.690 ;
        RECT 2652.000 2787.330 2652.260 2787.650 ;
        RECT 2899.020 2787.330 2899.280 2787.650 ;
        RECT 2899.080 2786.485 2899.220 2787.330 ;
        RECT 2899.010 2786.115 2899.290 2786.485 ;
      LAYER via2 ;
        RECT 2899.010 2786.160 2899.290 2786.440 ;
      LAYER met3 ;
        RECT 2898.985 2786.450 2899.315 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2898.985 2786.150 2924.800 2786.450 ;
        RECT 2898.985 2786.135 2899.315 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2651.510 3022.160 2651.830 3022.220 ;
        RECT 2898.990 3022.160 2899.310 3022.220 ;
        RECT 2651.510 3022.020 2899.310 3022.160 ;
        RECT 2651.510 3021.960 2651.830 3022.020 ;
        RECT 2898.990 3021.960 2899.310 3022.020 ;
      LAYER via ;
        RECT 2651.540 3021.960 2651.800 3022.220 ;
        RECT 2899.020 3021.960 2899.280 3022.220 ;
      LAYER met2 ;
        RECT 1640.910 3199.810 1641.190 3199.925 ;
        RECT 1641.760 3199.810 1642.040 3200.000 ;
        RECT 1640.910 3199.670 1642.040 3199.810 ;
        RECT 1640.910 3199.555 1641.190 3199.670 ;
        RECT 1641.760 3197.600 1642.040 3199.670 ;
        RECT 2651.530 3192.755 2651.810 3193.125 ;
        RECT 2651.600 3022.250 2651.740 3192.755 ;
        RECT 2651.540 3021.930 2651.800 3022.250 ;
        RECT 2899.020 3021.930 2899.280 3022.250 ;
        RECT 2899.080 3021.085 2899.220 3021.930 ;
        RECT 2899.010 3020.715 2899.290 3021.085 ;
      LAYER via2 ;
        RECT 1640.910 3199.600 1641.190 3199.880 ;
        RECT 2651.530 3192.800 2651.810 3193.080 ;
        RECT 2899.010 3020.760 2899.290 3021.040 ;
      LAYER met3 ;
        RECT 1640.885 3199.900 1641.215 3199.905 ;
        RECT 1640.630 3199.890 1641.215 3199.900 ;
        RECT 1640.430 3199.590 1641.215 3199.890 ;
        RECT 1640.630 3199.580 1641.215 3199.590 ;
        RECT 1640.885 3199.575 1641.215 3199.580 ;
        RECT 1640.630 3193.090 1641.010 3193.100 ;
        RECT 2651.505 3193.090 2651.835 3193.105 ;
        RECT 1640.630 3192.790 2651.835 3193.090 ;
        RECT 1640.630 3192.780 1641.010 3192.790 ;
        RECT 2651.505 3192.775 2651.835 3192.790 ;
        RECT 2898.985 3021.050 2899.315 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2898.985 3020.750 2924.800 3021.050 ;
        RECT 2898.985 3020.735 2899.315 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
      LAYER via3 ;
        RECT 1640.660 3199.580 1640.980 3199.900 ;
        RECT 1640.660 3192.780 1640.980 3193.100 ;
      LAYER met4 ;
        RECT 1640.655 3199.575 1640.985 3199.905 ;
        RECT 1640.670 3193.105 1640.970 3199.575 ;
        RECT 1640.655 3192.775 1640.985 3193.105 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1683.210 3250.300 1683.530 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1683.210 3250.160 2901.150 3250.300 ;
        RECT 1683.210 3250.100 1683.530 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 1683.240 3250.100 1683.500 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1683.240 3250.070 1683.500 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1681.320 3199.810 1681.600 3200.000 ;
        RECT 1683.300 3199.810 1683.440 3250.070 ;
        RECT 1681.320 3199.670 1683.440 3199.810 ;
        RECT 1681.320 3197.600 1681.600 3199.670 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1724.610 3484.900 1724.930 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1724.610 3484.760 2901.150 3484.900 ;
        RECT 1724.610 3484.700 1724.930 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 1724.640 3484.700 1724.900 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1724.640 3484.670 1724.900 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1720.880 3199.130 1721.160 3200.000 ;
        RECT 1724.700 3199.810 1724.840 3484.670 ;
        RECT 1723.780 3199.670 1724.840 3199.810 ;
        RECT 1723.780 3199.130 1723.920 3199.670 ;
        RECT 1720.880 3198.990 1723.920 3199.130 ;
        RECT 1720.880 3197.600 1721.160 3198.990 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1766.010 3501.220 1766.330 3501.280 ;
        RECT 2635.870 3501.220 2636.190 3501.280 ;
        RECT 1766.010 3501.080 2636.190 3501.220 ;
        RECT 1766.010 3501.020 1766.330 3501.080 ;
        RECT 2635.870 3501.020 2636.190 3501.080 ;
      LAYER via ;
        RECT 1766.040 3501.020 1766.300 3501.280 ;
        RECT 2635.900 3501.020 2636.160 3501.280 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.310 2636.100 3517.600 ;
        RECT 1766.040 3500.990 1766.300 3501.310 ;
        RECT 2635.900 3500.990 2636.160 3501.310 ;
        RECT 1766.100 3200.490 1766.240 3500.990 ;
        RECT 1762.880 3200.350 1766.240 3200.490 ;
        RECT 1759.980 3199.810 1760.260 3200.000 ;
        RECT 1762.880 3199.810 1763.020 3200.350 ;
        RECT 1759.980 3199.670 1763.020 3199.810 ;
        RECT 1759.980 3197.600 1760.260 3199.670 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.510 3500.200 1800.830 3500.260 ;
        RECT 2311.570 3500.200 2311.890 3500.260 ;
        RECT 1800.510 3500.060 2311.890 3500.200 ;
        RECT 1800.510 3500.000 1800.830 3500.060 ;
        RECT 2311.570 3500.000 2311.890 3500.060 ;
      LAYER via ;
        RECT 1800.540 3500.000 1800.800 3500.260 ;
        RECT 2311.600 3500.000 2311.860 3500.260 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3500.290 2311.800 3517.600 ;
        RECT 1800.540 3499.970 1800.800 3500.290 ;
        RECT 2311.600 3499.970 2311.860 3500.290 ;
        RECT 1799.540 3199.810 1799.820 3200.000 ;
        RECT 1800.600 3199.810 1800.740 3499.970 ;
        RECT 1799.540 3199.670 1800.740 3199.810 ;
        RECT 1799.540 3197.600 1799.820 3199.670 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1841.910 3498.500 1842.230 3498.560 ;
        RECT 1987.270 3498.500 1987.590 3498.560 ;
        RECT 1841.910 3498.360 1987.590 3498.500 ;
        RECT 1841.910 3498.300 1842.230 3498.360 ;
        RECT 1987.270 3498.300 1987.590 3498.360 ;
      LAYER via ;
        RECT 1841.940 3498.300 1842.200 3498.560 ;
        RECT 1987.300 3498.300 1987.560 3498.560 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3498.590 1987.500 3517.600 ;
        RECT 1841.940 3498.270 1842.200 3498.590 ;
        RECT 1987.300 3498.270 1987.560 3498.590 ;
        RECT 1839.100 3199.130 1839.380 3200.000 ;
        RECT 1842.000 3199.130 1842.140 3498.270 ;
        RECT 1839.100 3198.990 1842.140 3199.130 ;
        RECT 1839.100 3197.600 1839.380 3198.990 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 3499.520 1662.830 3499.580 ;
        RECT 1876.870 3499.520 1877.190 3499.580 ;
        RECT 1662.510 3499.380 1877.190 3499.520 ;
        RECT 1662.510 3499.320 1662.830 3499.380 ;
        RECT 1876.870 3499.320 1877.190 3499.380 ;
      LAYER via ;
        RECT 1662.540 3499.320 1662.800 3499.580 ;
        RECT 1876.900 3499.320 1877.160 3499.580 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3499.610 1662.740 3517.600 ;
        RECT 1662.540 3499.290 1662.800 3499.610 ;
        RECT 1876.900 3499.290 1877.160 3499.610 ;
        RECT 1876.960 3199.810 1877.100 3499.290 ;
        RECT 1878.660 3199.810 1878.940 3200.000 ;
        RECT 1876.960 3199.670 1878.940 3199.810 ;
        RECT 1878.660 3197.600 1878.940 3199.670 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3500.880 1338.530 3500.940 ;
        RECT 1918.270 3500.880 1918.590 3500.940 ;
        RECT 1338.210 3500.740 1918.590 3500.880 ;
        RECT 1338.210 3500.680 1338.530 3500.740 ;
        RECT 1918.270 3500.680 1918.590 3500.740 ;
      LAYER via ;
        RECT 1338.240 3500.680 1338.500 3500.940 ;
        RECT 1918.300 3500.680 1918.560 3500.940 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3500.970 1338.440 3517.600 ;
        RECT 1338.240 3500.650 1338.500 3500.970 ;
        RECT 1918.300 3500.650 1918.560 3500.970 ;
        RECT 1918.360 3200.000 1918.500 3500.650 ;
        RECT 1918.220 3197.600 1918.500 3200.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2898.990 3195.900 2899.310 3195.960 ;
        RECT 2901.750 3195.900 2902.070 3195.960 ;
        RECT 2898.990 3195.760 2902.070 3195.900 ;
        RECT 2898.990 3195.700 2899.310 3195.760 ;
        RECT 2901.750 3195.700 2902.070 3195.760 ;
      LAYER via ;
        RECT 2899.020 3195.700 2899.280 3195.960 ;
        RECT 2901.780 3195.700 2902.040 3195.960 ;
      LAYER met2 ;
        RECT 1207.590 3211.115 1207.870 3211.485 ;
        RECT 2899.010 3211.115 2899.290 3211.485 ;
        RECT 1207.660 3200.000 1207.800 3211.115 ;
        RECT 1207.520 3197.600 1207.800 3200.000 ;
        RECT 2899.080 3195.990 2899.220 3211.115 ;
        RECT 2899.020 3195.670 2899.280 3195.990 ;
        RECT 2901.780 3195.670 2902.040 3195.990 ;
        RECT 2901.840 439.805 2901.980 3195.670 ;
        RECT 2901.770 439.435 2902.050 439.805 ;
      LAYER via2 ;
        RECT 1207.590 3211.160 1207.870 3211.440 ;
        RECT 2899.010 3211.160 2899.290 3211.440 ;
        RECT 2901.770 439.480 2902.050 439.760 ;
      LAYER met3 ;
        RECT 1207.565 3211.450 1207.895 3211.465 ;
        RECT 2898.985 3211.450 2899.315 3211.465 ;
        RECT 1207.565 3211.150 2899.315 3211.450 ;
        RECT 1207.565 3211.135 1207.895 3211.150 ;
        RECT 2898.985 3211.135 2899.315 3211.150 ;
        RECT 2901.745 439.770 2902.075 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2901.745 439.470 2924.800 439.770 ;
        RECT 2901.745 439.455 2902.075 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3504.280 1014.230 3504.340 ;
        RECT 1952.770 3504.280 1953.090 3504.340 ;
        RECT 1013.910 3504.140 1953.090 3504.280 ;
        RECT 1013.910 3504.080 1014.230 3504.140 ;
        RECT 1952.770 3504.080 1953.090 3504.140 ;
      LAYER via ;
        RECT 1013.940 3504.080 1014.200 3504.340 ;
        RECT 1952.800 3504.080 1953.060 3504.340 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3504.370 1014.140 3517.600 ;
        RECT 1013.940 3504.050 1014.200 3504.370 ;
        RECT 1952.800 3504.050 1953.060 3504.370 ;
        RECT 1952.860 3200.490 1953.000 3504.050 ;
        RECT 1952.860 3200.350 1956.220 3200.490 ;
        RECT 1956.080 3199.810 1956.220 3200.350 ;
        RECT 1957.320 3199.810 1957.600 3200.000 ;
        RECT 1956.080 3199.670 1957.600 3199.810 ;
        RECT 1957.320 3197.600 1957.600 3199.670 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3503.260 689.470 3503.320 ;
        RECT 1994.170 3503.260 1994.490 3503.320 ;
        RECT 689.150 3503.120 1994.490 3503.260 ;
        RECT 689.150 3503.060 689.470 3503.120 ;
        RECT 1994.170 3503.060 1994.490 3503.120 ;
      LAYER via ;
        RECT 689.180 3503.060 689.440 3503.320 ;
        RECT 1994.200 3503.060 1994.460 3503.320 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.350 689.380 3517.600 ;
        RECT 689.180 3503.030 689.440 3503.350 ;
        RECT 1994.200 3503.030 1994.460 3503.350 ;
        RECT 1994.260 3199.130 1994.400 3503.030 ;
        RECT 1996.880 3199.130 1997.160 3200.000 ;
        RECT 1994.260 3198.990 1997.160 3199.130 ;
        RECT 1996.880 3197.600 1997.160 3198.990 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.240 365.170 3502.300 ;
        RECT 2035.570 3502.240 2035.890 3502.300 ;
        RECT 364.850 3502.100 2035.890 3502.240 ;
        RECT 364.850 3502.040 365.170 3502.100 ;
        RECT 2035.570 3502.040 2035.890 3502.100 ;
      LAYER via ;
        RECT 364.880 3502.040 365.140 3502.300 ;
        RECT 2035.600 3502.040 2035.860 3502.300 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3502.330 365.080 3517.600 ;
        RECT 364.880 3502.010 365.140 3502.330 ;
        RECT 2035.600 3502.010 2035.860 3502.330 ;
        RECT 2035.660 3199.810 2035.800 3502.010 ;
        RECT 2036.440 3199.810 2036.720 3200.000 ;
        RECT 2035.660 3199.670 2036.720 3199.810 ;
        RECT 2036.440 3197.600 2036.720 3199.670 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
        RECT 2070.090 3501.475 2070.370 3501.845 ;
        RECT 2070.160 3199.130 2070.300 3501.475 ;
        RECT 2076.000 3199.130 2076.280 3200.000 ;
        RECT 2070.160 3198.990 2076.280 3199.130 ;
        RECT 2076.000 3197.600 2076.280 3198.990 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
        RECT 2070.090 3501.520 2070.370 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 2070.065 3501.810 2070.395 3501.825 ;
        RECT 40.545 3501.510 2070.395 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 2070.065 3501.495 2070.395 3501.510 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 2111.470 3263.900 2111.790 3263.960 ;
        RECT 15.250 3263.760 2111.790 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 2111.470 3263.700 2111.790 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 2111.500 3263.700 2111.760 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 2111.500 3263.670 2111.760 3263.990 ;
        RECT 2111.560 3201.170 2111.700 3263.670 ;
        RECT 2111.560 3201.030 2114.000 3201.170 ;
        RECT 2113.860 3199.810 2114.000 3201.030 ;
        RECT 2115.560 3199.810 2115.840 3200.000 ;
        RECT 2113.860 3199.670 2115.840 3199.810 ;
        RECT 2115.560 3197.600 2115.840 3199.670 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3204.060 40.870 3204.120 ;
        RECT 2155.170 3204.060 2155.490 3204.120 ;
        RECT 40.550 3203.920 2155.490 3204.060 ;
        RECT 40.550 3203.860 40.870 3203.920 ;
        RECT 2155.170 3203.860 2155.490 3203.920 ;
        RECT 16.170 2980.340 16.490 2980.400 ;
        RECT 40.550 2980.340 40.870 2980.400 ;
        RECT 16.170 2980.200 40.870 2980.340 ;
        RECT 16.170 2980.140 16.490 2980.200 ;
        RECT 40.550 2980.140 40.870 2980.200 ;
      LAYER via ;
        RECT 40.580 3203.860 40.840 3204.120 ;
        RECT 2155.200 3203.860 2155.460 3204.120 ;
        RECT 16.200 2980.140 16.460 2980.400 ;
        RECT 40.580 2980.140 40.840 2980.400 ;
      LAYER met2 ;
        RECT 40.580 3203.830 40.840 3204.150 ;
        RECT 2155.200 3203.830 2155.460 3204.150 ;
        RECT 40.640 2980.430 40.780 3203.830 ;
        RECT 2155.260 3200.000 2155.400 3203.830 ;
        RECT 2155.120 3197.600 2155.400 3200.000 ;
        RECT 16.200 2980.285 16.460 2980.430 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 40.580 2980.110 40.840 2980.430 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 431.090 3211.540 431.410 3211.600 ;
        RECT 2194.270 3211.540 2194.590 3211.600 ;
        RECT 431.090 3211.400 2194.590 3211.540 ;
        RECT 431.090 3211.340 431.410 3211.400 ;
        RECT 2194.270 3211.340 2194.590 3211.400 ;
        RECT 16.170 2697.800 16.490 2697.860 ;
        RECT 431.090 2697.800 431.410 2697.860 ;
        RECT 16.170 2697.660 431.410 2697.800 ;
        RECT 16.170 2697.600 16.490 2697.660 ;
        RECT 431.090 2697.600 431.410 2697.660 ;
      LAYER via ;
        RECT 431.120 3211.340 431.380 3211.600 ;
        RECT 2194.300 3211.340 2194.560 3211.600 ;
        RECT 16.200 2697.600 16.460 2697.860 ;
        RECT 431.120 2697.600 431.380 2697.860 ;
      LAYER met2 ;
        RECT 431.120 3211.310 431.380 3211.630 ;
        RECT 2194.300 3211.310 2194.560 3211.630 ;
        RECT 431.180 2697.890 431.320 3211.310 ;
        RECT 2194.360 3200.000 2194.500 3211.310 ;
        RECT 2194.220 3197.600 2194.500 3200.000 ;
        RECT 16.200 2697.570 16.460 2697.890 ;
        RECT 431.120 2697.570 431.380 2697.890 ;
        RECT 16.260 2693.325 16.400 2697.570 ;
        RECT 16.190 2692.955 16.470 2693.325 ;
      LAYER via2 ;
        RECT 16.190 2693.000 16.470 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 16.165 2693.290 16.495 2693.305 ;
        RECT -4.800 2692.990 16.495 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 16.165 2692.975 16.495 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 39.630 3210.520 39.950 3210.580 ;
        RECT 2233.830 3210.520 2234.150 3210.580 ;
        RECT 39.630 3210.380 2234.150 3210.520 ;
        RECT 39.630 3210.320 39.950 3210.380 ;
        RECT 2233.830 3210.320 2234.150 3210.380 ;
        RECT 16.170 2405.740 16.490 2405.800 ;
        RECT 39.630 2405.740 39.950 2405.800 ;
        RECT 16.170 2405.600 39.950 2405.740 ;
        RECT 16.170 2405.540 16.490 2405.600 ;
        RECT 39.630 2405.540 39.950 2405.600 ;
      LAYER via ;
        RECT 39.660 3210.320 39.920 3210.580 ;
        RECT 2233.860 3210.320 2234.120 3210.580 ;
        RECT 16.200 2405.540 16.460 2405.800 ;
        RECT 39.660 2405.540 39.920 2405.800 ;
      LAYER met2 ;
        RECT 39.660 3210.290 39.920 3210.610 ;
        RECT 2233.860 3210.290 2234.120 3210.610 ;
        RECT 39.720 2405.830 39.860 3210.290 ;
        RECT 2233.920 3200.000 2234.060 3210.290 ;
        RECT 2233.780 3197.600 2234.060 3200.000 ;
        RECT 16.200 2405.685 16.460 2405.830 ;
        RECT 16.190 2405.315 16.470 2405.685 ;
        RECT 39.660 2405.510 39.920 2405.830 ;
      LAYER via2 ;
        RECT 16.190 2405.360 16.470 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 16.165 2405.650 16.495 2405.665 ;
        RECT -4.800 2405.350 16.495 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 16.165 2405.335 16.495 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2194.730 3211.540 2195.050 3211.600 ;
        RECT 2273.390 3211.540 2273.710 3211.600 ;
        RECT 2194.730 3211.400 2273.710 3211.540 ;
        RECT 2194.730 3211.340 2195.050 3211.400 ;
        RECT 2273.390 3211.340 2273.710 3211.400 ;
        RECT 16.630 3198.620 16.950 3198.680 ;
        RECT 2194.730 3198.620 2195.050 3198.680 ;
        RECT 16.630 3198.480 2195.050 3198.620 ;
        RECT 16.630 3198.420 16.950 3198.480 ;
        RECT 2194.730 3198.420 2195.050 3198.480 ;
      LAYER via ;
        RECT 2194.760 3211.340 2195.020 3211.600 ;
        RECT 2273.420 3211.340 2273.680 3211.600 ;
        RECT 16.660 3198.420 16.920 3198.680 ;
        RECT 2194.760 3198.420 2195.020 3198.680 ;
      LAYER met2 ;
        RECT 2194.760 3211.310 2195.020 3211.630 ;
        RECT 2273.420 3211.310 2273.680 3211.630 ;
        RECT 2194.820 3198.710 2194.960 3211.310 ;
        RECT 2273.480 3200.000 2273.620 3211.310 ;
        RECT 16.660 3198.390 16.920 3198.710 ;
        RECT 2194.760 3198.390 2195.020 3198.710 ;
        RECT 16.720 2118.725 16.860 3198.390 ;
        RECT 2273.340 3197.600 2273.620 3200.000 ;
        RECT 16.650 2118.355 16.930 2118.725 ;
      LAYER via2 ;
        RECT 16.650 2118.400 16.930 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.625 2118.690 16.955 2118.705 ;
        RECT -4.800 2118.390 16.955 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.625 2118.375 16.955 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 38.250 3209.840 38.570 3209.900 ;
        RECT 2312.950 3209.840 2313.270 3209.900 ;
        RECT 38.250 3209.700 2313.270 3209.840 ;
        RECT 38.250 3209.640 38.570 3209.700 ;
        RECT 2312.950 3209.640 2313.270 3209.700 ;
        RECT 16.630 1832.500 16.950 1832.560 ;
        RECT 38.250 1832.500 38.570 1832.560 ;
        RECT 16.630 1832.360 38.570 1832.500 ;
        RECT 16.630 1832.300 16.950 1832.360 ;
        RECT 38.250 1832.300 38.570 1832.360 ;
      LAYER via ;
        RECT 38.280 3209.640 38.540 3209.900 ;
        RECT 2312.980 3209.640 2313.240 3209.900 ;
        RECT 16.660 1832.300 16.920 1832.560 ;
        RECT 38.280 1832.300 38.540 1832.560 ;
      LAYER met2 ;
        RECT 38.280 3209.610 38.540 3209.930 ;
        RECT 2312.980 3209.610 2313.240 3209.930 ;
        RECT 38.340 1832.590 38.480 3209.610 ;
        RECT 2313.040 3200.000 2313.180 3209.610 ;
        RECT 2312.900 3197.600 2313.180 3200.000 ;
        RECT 16.660 1832.270 16.920 1832.590 ;
        RECT 38.280 1832.270 38.540 1832.590 ;
        RECT 16.720 1831.085 16.860 1832.270 ;
        RECT 16.650 1830.715 16.930 1831.085 ;
      LAYER via2 ;
        RECT 16.650 1830.760 16.930 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 16.625 1831.050 16.955 1831.065 ;
        RECT -4.800 1830.750 16.955 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 16.625 1830.735 16.955 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1421.470 670.380 1421.790 670.440 ;
        RECT 1468.850 670.380 1469.170 670.440 ;
        RECT 1421.470 670.240 1469.170 670.380 ;
        RECT 1421.470 670.180 1421.790 670.240 ;
        RECT 1468.850 670.180 1469.170 670.240 ;
        RECT 2572.850 670.380 2573.170 670.440 ;
        RECT 2574.230 670.380 2574.550 670.440 ;
        RECT 2572.850 670.240 2574.550 670.380 ;
        RECT 2572.850 670.180 2573.170 670.240 ;
        RECT 2574.230 670.180 2574.550 670.240 ;
        RECT 2704.870 669.700 2705.190 669.760 ;
        RECT 2729.250 669.700 2729.570 669.760 ;
        RECT 2704.870 669.560 2729.570 669.700 ;
        RECT 2704.870 669.500 2705.190 669.560 ;
        RECT 2729.250 669.500 2729.570 669.560 ;
        RECT 1628.010 669.360 1628.330 669.420 ;
        RECT 1669.410 669.360 1669.730 669.420 ;
        RECT 1628.010 669.220 1669.730 669.360 ;
        RECT 1628.010 669.160 1628.330 669.220 ;
        RECT 1669.410 669.160 1669.730 669.220 ;
        RECT 1742.090 668.680 1742.410 668.740 ;
        RECT 1772.910 668.680 1773.230 668.740 ;
        RECT 1742.090 668.540 1773.230 668.680 ;
        RECT 1742.090 668.480 1742.410 668.540 ;
        RECT 1772.910 668.480 1773.230 668.540 ;
      LAYER via ;
        RECT 1421.500 670.180 1421.760 670.440 ;
        RECT 1468.880 670.180 1469.140 670.440 ;
        RECT 2572.880 670.180 2573.140 670.440 ;
        RECT 2574.260 670.180 2574.520 670.440 ;
        RECT 2704.900 669.500 2705.160 669.760 ;
        RECT 2729.280 669.500 2729.540 669.760 ;
        RECT 1628.040 669.160 1628.300 669.420 ;
        RECT 1669.440 669.160 1669.700 669.420 ;
        RECT 1742.120 668.480 1742.380 668.740 ;
        RECT 1772.940 668.480 1773.200 668.740 ;
      LAYER met2 ;
        RECT 1247.080 3199.130 1247.360 3200.000 ;
        RECT 1247.610 3199.130 1247.890 3199.245 ;
        RECT 1247.080 3198.990 1247.890 3199.130 ;
        RECT 1247.080 3197.600 1247.360 3198.990 ;
        RECT 1247.610 3198.875 1247.890 3198.990 ;
        RECT 1246.230 1538.315 1246.510 1538.685 ;
        RECT 1246.300 1491.765 1246.440 1538.315 ;
        RECT 1246.230 1491.395 1246.510 1491.765 ;
        RECT 1246.230 1398.915 1246.510 1399.285 ;
        RECT 1246.300 1353.045 1246.440 1398.915 ;
        RECT 1246.230 1352.675 1246.510 1353.045 ;
        RECT 1246.230 1351.995 1246.510 1352.365 ;
        RECT 1246.300 1304.765 1246.440 1351.995 ;
        RECT 1246.230 1304.395 1246.510 1304.765 ;
        RECT 1246.230 1255.435 1246.510 1255.805 ;
        RECT 1246.300 1208.885 1246.440 1255.435 ;
        RECT 1246.230 1208.515 1246.510 1208.885 ;
        RECT 1247.150 1110.595 1247.430 1110.965 ;
        RECT 1247.220 1072.885 1247.360 1110.595 ;
        RECT 1247.150 1072.515 1247.430 1072.885 ;
        RECT 1247.610 999.075 1247.890 999.445 ;
        RECT 1247.680 928.045 1247.820 999.075 ;
        RECT 1247.610 927.675 1247.890 928.045 ;
        RECT 1248.070 896.395 1248.350 896.765 ;
        RECT 1248.140 849.845 1248.280 896.395 ;
        RECT 1248.070 849.475 1248.350 849.845 ;
        RECT 1907.250 672.675 1907.530 673.045 ;
        RECT 1572.830 671.995 1573.110 672.365 ;
        RECT 1468.870 671.315 1469.150 671.685 ;
        RECT 1476.230 671.315 1476.510 671.685 ;
        RECT 1468.940 670.470 1469.080 671.315 ;
        RECT 1421.500 670.325 1421.760 670.470 ;
        RECT 1421.490 669.955 1421.770 670.325 ;
        RECT 1468.880 670.150 1469.140 670.470 ;
        RECT 1476.300 669.645 1476.440 671.315 ;
        RECT 1572.900 671.005 1573.040 671.995 ;
        RECT 1572.830 670.635 1573.110 671.005 ;
        RECT 1907.320 670.325 1907.460 672.675 ;
        RECT 2076.530 671.315 2076.810 671.685 ;
        RECT 2076.600 671.005 2076.740 671.315 ;
        RECT 1979.930 670.635 1980.210 671.005 ;
        RECT 2076.530 670.635 2076.810 671.005 ;
        RECT 2137.710 670.890 2137.990 671.005 ;
        RECT 2138.630 670.890 2138.910 671.005 ;
        RECT 2137.710 670.750 2138.910 670.890 ;
        RECT 2137.710 670.635 2137.990 670.750 ;
        RECT 2138.630 670.635 2138.910 670.750 ;
        RECT 2772.510 670.635 2772.790 671.005 ;
        RECT 1907.250 669.955 1907.530 670.325 ;
        RECT 1476.230 669.275 1476.510 669.645 ;
        RECT 1628.030 669.275 1628.310 669.645 ;
        RECT 1669.430 669.275 1669.710 669.645 ;
        RECT 1628.040 669.130 1628.300 669.275 ;
        RECT 1669.440 669.130 1669.700 669.275 ;
        RECT 1980.000 668.965 1980.140 670.635 ;
        RECT 2572.880 670.325 2573.140 670.470 ;
        RECT 2574.260 670.325 2574.520 670.470 ;
        RECT 2294.110 669.955 2294.390 670.325 ;
        RECT 2572.870 669.955 2573.150 670.325 ;
        RECT 2574.250 669.955 2574.530 670.325 ;
        RECT 2729.270 669.955 2729.550 670.325 ;
        RECT 2294.180 668.965 2294.320 669.955 ;
        RECT 2729.340 669.790 2729.480 669.955 ;
        RECT 2704.900 669.645 2705.160 669.790 ;
        RECT 2704.890 669.275 2705.170 669.645 ;
        RECT 2729.280 669.470 2729.540 669.790 ;
        RECT 2772.580 668.965 2772.720 670.635 ;
        RECT 2863.130 669.955 2863.410 670.325 ;
        RECT 2863.200 669.530 2863.340 669.955 ;
        RECT 2863.590 669.530 2863.870 669.645 ;
        RECT 2863.200 669.390 2863.870 669.530 ;
        RECT 2863.590 669.275 2863.870 669.390 ;
        RECT 1742.120 668.450 1742.380 668.770 ;
        RECT 1772.940 668.450 1773.200 668.770 ;
        RECT 1979.930 668.595 1980.210 668.965 ;
        RECT 2294.110 668.595 2294.390 668.965 ;
        RECT 2772.510 668.595 2772.790 668.965 ;
        RECT 1742.180 668.285 1742.320 668.450 ;
        RECT 1773.000 668.285 1773.140 668.450 ;
        RECT 1742.110 667.915 1742.390 668.285 ;
        RECT 1772.930 667.915 1773.210 668.285 ;
      LAYER via2 ;
        RECT 1247.610 3198.920 1247.890 3199.200 ;
        RECT 1246.230 1538.360 1246.510 1538.640 ;
        RECT 1246.230 1491.440 1246.510 1491.720 ;
        RECT 1246.230 1398.960 1246.510 1399.240 ;
        RECT 1246.230 1352.720 1246.510 1353.000 ;
        RECT 1246.230 1352.040 1246.510 1352.320 ;
        RECT 1246.230 1304.440 1246.510 1304.720 ;
        RECT 1246.230 1255.480 1246.510 1255.760 ;
        RECT 1246.230 1208.560 1246.510 1208.840 ;
        RECT 1247.150 1110.640 1247.430 1110.920 ;
        RECT 1247.150 1072.560 1247.430 1072.840 ;
        RECT 1247.610 999.120 1247.890 999.400 ;
        RECT 1247.610 927.720 1247.890 928.000 ;
        RECT 1248.070 896.440 1248.350 896.720 ;
        RECT 1248.070 849.520 1248.350 849.800 ;
        RECT 1907.250 672.720 1907.530 673.000 ;
        RECT 1572.830 672.040 1573.110 672.320 ;
        RECT 1468.870 671.360 1469.150 671.640 ;
        RECT 1476.230 671.360 1476.510 671.640 ;
        RECT 1421.490 670.000 1421.770 670.280 ;
        RECT 1572.830 670.680 1573.110 670.960 ;
        RECT 2076.530 671.360 2076.810 671.640 ;
        RECT 1979.930 670.680 1980.210 670.960 ;
        RECT 2076.530 670.680 2076.810 670.960 ;
        RECT 2137.710 670.680 2137.990 670.960 ;
        RECT 2138.630 670.680 2138.910 670.960 ;
        RECT 2772.510 670.680 2772.790 670.960 ;
        RECT 1907.250 670.000 1907.530 670.280 ;
        RECT 1476.230 669.320 1476.510 669.600 ;
        RECT 1628.030 669.320 1628.310 669.600 ;
        RECT 1669.430 669.320 1669.710 669.600 ;
        RECT 2294.110 670.000 2294.390 670.280 ;
        RECT 2572.870 670.000 2573.150 670.280 ;
        RECT 2574.250 670.000 2574.530 670.280 ;
        RECT 2729.270 670.000 2729.550 670.280 ;
        RECT 2704.890 669.320 2705.170 669.600 ;
        RECT 2863.130 670.000 2863.410 670.280 ;
        RECT 2863.590 669.320 2863.870 669.600 ;
        RECT 1979.930 668.640 1980.210 668.920 ;
        RECT 2294.110 668.640 2294.390 668.920 ;
        RECT 2772.510 668.640 2772.790 668.920 ;
        RECT 1742.110 667.960 1742.390 668.240 ;
        RECT 1772.930 667.960 1773.210 668.240 ;
      LAYER met3 ;
        RECT 1246.870 3199.210 1247.250 3199.220 ;
        RECT 1247.585 3199.210 1247.915 3199.225 ;
        RECT 1246.870 3198.910 1247.915 3199.210 ;
        RECT 1246.870 3198.900 1247.250 3198.910 ;
        RECT 1247.585 3198.895 1247.915 3198.910 ;
        RECT 1246.205 1538.650 1246.535 1538.665 ;
        RECT 1246.870 1538.650 1247.250 1538.660 ;
        RECT 1246.205 1538.350 1247.250 1538.650 ;
        RECT 1246.205 1538.335 1246.535 1538.350 ;
        RECT 1246.870 1538.340 1247.250 1538.350 ;
        RECT 1246.205 1491.730 1246.535 1491.745 ;
        RECT 1245.990 1491.415 1246.535 1491.730 ;
        RECT 1245.990 1491.060 1246.290 1491.415 ;
        RECT 1245.950 1490.740 1246.330 1491.060 ;
        RECT 1245.950 1449.260 1246.330 1449.580 ;
        RECT 1245.990 1448.210 1246.290 1449.260 ;
        RECT 1247.790 1448.210 1248.170 1448.220 ;
        RECT 1245.990 1447.910 1248.170 1448.210 ;
        RECT 1247.790 1447.900 1248.170 1447.910 ;
        RECT 1246.205 1399.260 1246.535 1399.265 ;
        RECT 1245.950 1399.250 1246.535 1399.260 ;
        RECT 1245.750 1398.950 1246.535 1399.250 ;
        RECT 1245.950 1398.940 1246.535 1398.950 ;
        RECT 1246.205 1398.935 1246.535 1398.940 ;
        RECT 1246.205 1353.010 1246.535 1353.025 ;
        RECT 1246.870 1353.010 1247.250 1353.020 ;
        RECT 1246.205 1352.710 1247.250 1353.010 ;
        RECT 1246.205 1352.695 1246.535 1352.710 ;
        RECT 1246.870 1352.700 1247.250 1352.710 ;
        RECT 1246.205 1352.330 1246.535 1352.345 ;
        RECT 1246.870 1352.330 1247.250 1352.340 ;
        RECT 1246.205 1352.030 1247.250 1352.330 ;
        RECT 1246.205 1352.015 1246.535 1352.030 ;
        RECT 1246.870 1352.020 1247.250 1352.030 ;
        RECT 1246.205 1304.730 1246.535 1304.745 ;
        RECT 1245.990 1304.415 1246.535 1304.730 ;
        RECT 1245.990 1303.370 1246.290 1304.415 ;
        RECT 1247.790 1303.370 1248.170 1303.380 ;
        RECT 1245.990 1303.070 1248.170 1303.370 ;
        RECT 1247.790 1303.060 1248.170 1303.070 ;
        RECT 1246.205 1255.770 1246.535 1255.785 ;
        RECT 1246.870 1255.770 1247.250 1255.780 ;
        RECT 1246.205 1255.470 1247.250 1255.770 ;
        RECT 1246.205 1255.455 1246.535 1255.470 ;
        RECT 1246.870 1255.460 1247.250 1255.470 ;
        RECT 1246.205 1208.850 1246.535 1208.865 ;
        RECT 1245.990 1208.535 1246.535 1208.850 ;
        RECT 1245.990 1208.180 1246.290 1208.535 ;
        RECT 1245.950 1207.860 1246.330 1208.180 ;
        RECT 1245.950 1159.890 1246.330 1159.900 ;
        RECT 1246.870 1159.890 1247.250 1159.900 ;
        RECT 1245.950 1159.590 1247.250 1159.890 ;
        RECT 1245.950 1159.580 1246.330 1159.590 ;
        RECT 1246.870 1159.580 1247.250 1159.590 ;
        RECT 1246.870 1111.610 1247.250 1111.620 ;
        RECT 1246.870 1111.310 1248.130 1111.610 ;
        RECT 1246.870 1111.300 1247.250 1111.310 ;
        RECT 1247.125 1110.930 1247.455 1110.945 ;
        RECT 1247.830 1110.930 1248.130 1111.310 ;
        RECT 1247.125 1110.630 1248.130 1110.930 ;
        RECT 1247.125 1110.615 1247.455 1110.630 ;
        RECT 1247.125 1072.860 1247.455 1072.865 ;
        RECT 1246.870 1072.850 1247.455 1072.860 ;
        RECT 1246.670 1072.550 1247.455 1072.850 ;
        RECT 1246.870 1072.540 1247.455 1072.550 ;
        RECT 1247.125 1072.535 1247.455 1072.540 ;
        RECT 1247.790 999.780 1248.170 1000.100 ;
        RECT 1247.830 999.425 1248.130 999.780 ;
        RECT 1247.585 999.110 1248.130 999.425 ;
        RECT 1247.585 999.095 1247.915 999.110 ;
        RECT 1247.585 928.020 1247.915 928.025 ;
        RECT 1247.585 928.010 1248.170 928.020 ;
        RECT 1247.360 927.710 1248.170 928.010 ;
        RECT 1247.585 927.700 1248.170 927.710 ;
        RECT 1247.585 927.695 1247.915 927.700 ;
        RECT 1248.045 896.740 1248.375 896.745 ;
        RECT 1247.790 896.730 1248.375 896.740 ;
        RECT 1247.790 896.430 1248.600 896.730 ;
        RECT 1247.790 896.420 1248.375 896.430 ;
        RECT 1248.045 896.415 1248.375 896.420 ;
        RECT 1248.045 849.810 1248.375 849.825 ;
        RECT 1247.830 849.495 1248.375 849.810 ;
        RECT 1247.830 849.140 1248.130 849.495 ;
        RECT 1247.790 848.820 1248.170 849.140 ;
        RECT 1247.790 835.220 1248.170 835.540 ;
        RECT 1247.830 834.860 1248.130 835.220 ;
        RECT 1247.790 834.540 1248.170 834.860 ;
        RECT 1248.710 772.660 1249.090 772.980 ;
        RECT 1248.750 772.300 1249.050 772.660 ;
        RECT 1248.710 771.980 1249.090 772.300 ;
        RECT 1246.870 724.690 1247.250 724.700 ;
        RECT 1248.710 724.690 1249.090 724.700 ;
        RECT 1246.870 724.390 1249.090 724.690 ;
        RECT 1246.870 724.380 1247.250 724.390 ;
        RECT 1248.710 724.380 1249.090 724.390 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2916.710 674.070 2924.800 674.370 ;
        RECT 1883.510 673.010 1883.890 673.020 ;
        RECT 1907.225 673.010 1907.555 673.025 ;
        RECT 1883.510 672.710 1907.555 673.010 ;
        RECT 1883.510 672.700 1883.890 672.710 ;
        RECT 1907.225 672.695 1907.555 672.710 ;
        RECT 1524.710 672.330 1525.090 672.340 ;
        RECT 1572.805 672.330 1573.135 672.345 ;
        RECT 1524.710 672.030 1573.135 672.330 ;
        RECT 1524.710 672.020 1525.090 672.030 ;
        RECT 1572.805 672.015 1573.135 672.030 ;
        RECT 2088.710 672.030 2124.890 672.330 ;
        RECT 1468.845 671.650 1469.175 671.665 ;
        RECT 1476.205 671.650 1476.535 671.665 ;
        RECT 1468.845 671.350 1476.535 671.650 ;
        RECT 1468.845 671.335 1469.175 671.350 ;
        RECT 1476.205 671.335 1476.535 671.350 ;
        RECT 1835.670 671.650 1836.050 671.660 ;
        RECT 1883.510 671.650 1883.890 671.660 ;
        RECT 2076.505 671.650 2076.835 671.665 ;
        RECT 1835.670 671.350 1883.890 671.650 ;
        RECT 1835.670 671.340 1836.050 671.350 ;
        RECT 1883.510 671.340 1883.890 671.350 ;
        RECT 2041.790 671.350 2076.835 671.650 ;
        RECT 1572.805 670.970 1573.135 670.985 ;
        RECT 1579.910 670.970 1580.290 670.980 ;
        RECT 1572.805 670.670 1580.290 670.970 ;
        RECT 1572.805 670.655 1573.135 670.670 ;
        RECT 1579.910 670.660 1580.290 670.670 ;
        RECT 1979.905 670.970 1980.235 670.985 ;
        RECT 2041.790 670.970 2042.090 671.350 ;
        RECT 2076.505 671.335 2076.835 671.350 ;
        RECT 1979.905 670.670 2042.090 670.970 ;
        RECT 2076.505 670.970 2076.835 670.985 ;
        RECT 2088.710 670.970 2089.010 672.030 ;
        RECT 2076.505 670.670 2089.010 670.970 ;
        RECT 2124.590 670.970 2124.890 672.030 ;
        RECT 2463.150 671.350 2511.290 671.650 ;
        RECT 2137.685 670.970 2138.015 670.985 ;
        RECT 2124.590 670.670 2138.015 670.970 ;
        RECT 1979.905 670.655 1980.235 670.670 ;
        RECT 2076.505 670.655 2076.835 670.670 ;
        RECT 2137.685 670.655 2138.015 670.670 ;
        RECT 2138.605 670.970 2138.935 670.985 ;
        RECT 2138.605 670.670 2187.450 670.970 ;
        RECT 2138.605 670.655 2138.935 670.670 ;
        RECT 1421.465 670.290 1421.795 670.305 ;
        RECT 1297.510 669.990 1421.795 670.290 ;
        RECT 1246.870 669.610 1247.250 669.620 ;
        RECT 1297.510 669.610 1297.810 669.990 ;
        RECT 1421.465 669.975 1421.795 669.990 ;
        RECT 1786.910 670.290 1787.290 670.300 ;
        RECT 1835.670 670.290 1836.050 670.300 ;
        RECT 1786.910 669.990 1836.050 670.290 ;
        RECT 1786.910 669.980 1787.290 669.990 ;
        RECT 1835.670 669.980 1836.050 669.990 ;
        RECT 1907.225 670.290 1907.555 670.305 ;
        RECT 1907.225 669.990 1932.610 670.290 ;
        RECT 1907.225 669.975 1907.555 669.990 ;
        RECT 1246.870 669.310 1297.810 669.610 ;
        RECT 1476.205 669.610 1476.535 669.625 ;
        RECT 1579.910 669.610 1580.290 669.620 ;
        RECT 1628.005 669.610 1628.335 669.625 ;
        RECT 1476.205 669.310 1477.210 669.610 ;
        RECT 1246.870 669.300 1247.250 669.310 ;
        RECT 1476.205 669.295 1476.535 669.310 ;
        RECT 1476.910 668.930 1477.210 669.310 ;
        RECT 1498.070 669.310 1525.050 669.610 ;
        RECT 1498.070 668.930 1498.370 669.310 ;
        RECT 1524.750 668.940 1525.050 669.310 ;
        RECT 1579.910 669.310 1628.335 669.610 ;
        RECT 1579.910 669.300 1580.290 669.310 ;
        RECT 1628.005 669.295 1628.335 669.310 ;
        RECT 1669.405 669.610 1669.735 669.625 ;
        RECT 1717.910 669.610 1718.290 669.620 ;
        RECT 1669.405 669.310 1718.290 669.610 ;
        RECT 1669.405 669.295 1669.735 669.310 ;
        RECT 1717.910 669.300 1718.290 669.310 ;
        RECT 1476.910 668.630 1498.370 668.930 ;
        RECT 1524.710 668.620 1525.090 668.940 ;
        RECT 1932.310 668.930 1932.610 669.990 ;
        RECT 2187.150 669.610 2187.450 670.670 ;
        RECT 2269.910 670.290 2270.290 670.300 ;
        RECT 2235.910 669.990 2270.290 670.290 ;
        RECT 2235.910 669.610 2236.210 669.990 ;
        RECT 2269.910 669.980 2270.290 669.990 ;
        RECT 2294.085 670.290 2294.415 670.305 ;
        RECT 2366.510 670.290 2366.890 670.300 ;
        RECT 2463.150 670.290 2463.450 671.350 ;
        RECT 2510.990 670.980 2511.290 671.350 ;
        RECT 2510.950 670.660 2511.330 670.980 ;
        RECT 2772.485 670.970 2772.815 670.985 ;
        RECT 2772.485 670.670 2815.810 670.970 ;
        RECT 2772.485 670.655 2772.815 670.670 ;
        RECT 2572.845 670.290 2573.175 670.305 ;
        RECT 2294.085 669.990 2331.890 670.290 ;
        RECT 2294.085 669.975 2294.415 669.990 ;
        RECT 2187.150 669.310 2236.210 669.610 ;
        RECT 2331.590 669.610 2331.890 669.990 ;
        RECT 2332.510 669.990 2366.890 670.290 ;
        RECT 2332.510 669.610 2332.810 669.990 ;
        RECT 2366.510 669.980 2366.890 669.990 ;
        RECT 2429.110 669.990 2463.450 670.290 ;
        RECT 2525.710 669.990 2573.175 670.290 ;
        RECT 2429.110 669.610 2429.410 669.990 ;
        RECT 2331.590 669.310 2332.810 669.610 ;
        RECT 2414.390 669.310 2429.410 669.610 ;
        RECT 2510.950 669.610 2511.330 669.620 ;
        RECT 2525.710 669.610 2526.010 669.990 ;
        RECT 2572.845 669.975 2573.175 669.990 ;
        RECT 2574.225 670.290 2574.555 670.305 ;
        RECT 2656.310 670.290 2656.690 670.300 ;
        RECT 2574.225 669.990 2621.690 670.290 ;
        RECT 2574.225 669.975 2574.555 669.990 ;
        RECT 2510.950 669.310 2526.010 669.610 ;
        RECT 2621.390 669.610 2621.690 669.990 ;
        RECT 2622.310 669.990 2656.690 670.290 ;
        RECT 2622.310 669.610 2622.610 669.990 ;
        RECT 2656.310 669.980 2656.690 669.990 ;
        RECT 2729.245 670.290 2729.575 670.305 ;
        RECT 2752.910 670.290 2753.290 670.300 ;
        RECT 2729.245 669.990 2753.290 670.290 ;
        RECT 2729.245 669.975 2729.575 669.990 ;
        RECT 2752.910 669.980 2753.290 669.990 ;
        RECT 2704.865 669.610 2705.195 669.625 ;
        RECT 2621.390 669.310 2622.610 669.610 ;
        RECT 2704.190 669.310 2705.195 669.610 ;
        RECT 2815.510 669.610 2815.810 670.670 ;
        RECT 2863.105 670.290 2863.435 670.305 ;
        RECT 2916.710 670.290 2917.010 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
        RECT 2849.550 669.990 2863.435 670.290 ;
        RECT 2849.550 669.610 2849.850 669.990 ;
        RECT 2863.105 669.975 2863.435 669.990 ;
        RECT 2884.510 669.990 2917.010 670.290 ;
        RECT 2815.510 669.310 2849.850 669.610 ;
        RECT 2863.565 669.610 2863.895 669.625 ;
        RECT 2884.510 669.610 2884.810 669.990 ;
        RECT 2863.565 669.310 2884.810 669.610 ;
        RECT 1979.905 668.930 1980.235 668.945 ;
        RECT 1932.310 668.630 1980.235 668.930 ;
        RECT 1979.905 668.615 1980.235 668.630 ;
        RECT 2269.910 668.930 2270.290 668.940 ;
        RECT 2294.085 668.930 2294.415 668.945 ;
        RECT 2269.910 668.630 2294.415 668.930 ;
        RECT 2269.910 668.620 2270.290 668.630 ;
        RECT 2294.085 668.615 2294.415 668.630 ;
        RECT 1717.910 668.250 1718.290 668.260 ;
        RECT 1742.085 668.250 1742.415 668.265 ;
        RECT 1717.910 667.950 1742.415 668.250 ;
        RECT 1717.910 667.940 1718.290 667.950 ;
        RECT 1742.085 667.935 1742.415 667.950 ;
        RECT 1772.905 668.250 1773.235 668.265 ;
        RECT 1785.990 668.250 1786.370 668.260 ;
        RECT 1772.905 667.950 1786.370 668.250 ;
        RECT 1772.905 667.935 1773.235 667.950 ;
        RECT 1785.990 667.940 1786.370 667.950 ;
        RECT 2366.510 668.250 2366.890 668.260 ;
        RECT 2414.390 668.250 2414.690 669.310 ;
        RECT 2510.950 669.300 2511.330 669.310 ;
        RECT 2366.510 667.950 2414.690 668.250 ;
        RECT 2656.310 668.250 2656.690 668.260 ;
        RECT 2704.190 668.250 2704.490 669.310 ;
        RECT 2704.865 669.295 2705.195 669.310 ;
        RECT 2863.565 669.295 2863.895 669.310 ;
        RECT 2752.910 668.930 2753.290 668.940 ;
        RECT 2772.485 668.930 2772.815 668.945 ;
        RECT 2752.910 668.630 2772.815 668.930 ;
        RECT 2752.910 668.620 2753.290 668.630 ;
        RECT 2772.485 668.615 2772.815 668.630 ;
        RECT 2656.310 667.950 2704.490 668.250 ;
        RECT 2366.510 667.940 2366.890 667.950 ;
        RECT 2656.310 667.940 2656.690 667.950 ;
      LAYER via3 ;
        RECT 1246.900 3198.900 1247.220 3199.220 ;
        RECT 1246.900 1538.340 1247.220 1538.660 ;
        RECT 1245.980 1490.740 1246.300 1491.060 ;
        RECT 1245.980 1449.260 1246.300 1449.580 ;
        RECT 1247.820 1447.900 1248.140 1448.220 ;
        RECT 1245.980 1398.940 1246.300 1399.260 ;
        RECT 1246.900 1352.700 1247.220 1353.020 ;
        RECT 1246.900 1352.020 1247.220 1352.340 ;
        RECT 1247.820 1303.060 1248.140 1303.380 ;
        RECT 1246.900 1255.460 1247.220 1255.780 ;
        RECT 1245.980 1207.860 1246.300 1208.180 ;
        RECT 1245.980 1159.580 1246.300 1159.900 ;
        RECT 1246.900 1159.580 1247.220 1159.900 ;
        RECT 1246.900 1111.300 1247.220 1111.620 ;
        RECT 1246.900 1072.540 1247.220 1072.860 ;
        RECT 1247.820 999.780 1248.140 1000.100 ;
        RECT 1247.820 927.700 1248.140 928.020 ;
        RECT 1247.820 896.420 1248.140 896.740 ;
        RECT 1247.820 848.820 1248.140 849.140 ;
        RECT 1247.820 835.220 1248.140 835.540 ;
        RECT 1247.820 834.540 1248.140 834.860 ;
        RECT 1248.740 772.660 1249.060 772.980 ;
        RECT 1248.740 771.980 1249.060 772.300 ;
        RECT 1246.900 724.380 1247.220 724.700 ;
        RECT 1248.740 724.380 1249.060 724.700 ;
        RECT 1883.540 672.700 1883.860 673.020 ;
        RECT 1524.740 672.020 1525.060 672.340 ;
        RECT 1835.700 671.340 1836.020 671.660 ;
        RECT 1883.540 671.340 1883.860 671.660 ;
        RECT 1579.940 670.660 1580.260 670.980 ;
        RECT 1246.900 669.300 1247.220 669.620 ;
        RECT 1786.940 669.980 1787.260 670.300 ;
        RECT 1835.700 669.980 1836.020 670.300 ;
        RECT 1579.940 669.300 1580.260 669.620 ;
        RECT 1717.940 669.300 1718.260 669.620 ;
        RECT 1524.740 668.620 1525.060 668.940 ;
        RECT 2269.940 669.980 2270.260 670.300 ;
        RECT 2366.540 669.980 2366.860 670.300 ;
        RECT 2510.980 670.660 2511.300 670.980 ;
        RECT 2269.940 668.620 2270.260 668.940 ;
        RECT 1717.940 667.940 1718.260 668.260 ;
        RECT 1786.020 667.940 1786.340 668.260 ;
        RECT 2366.540 667.940 2366.860 668.260 ;
        RECT 2510.980 669.300 2511.300 669.620 ;
        RECT 2656.340 669.980 2656.660 670.300 ;
        RECT 2752.940 669.980 2753.260 670.300 ;
        RECT 2656.340 667.940 2656.660 668.260 ;
        RECT 2752.940 668.620 2753.260 668.940 ;
      LAYER met4 ;
        RECT 1246.895 3198.895 1247.225 3199.225 ;
        RECT 1246.910 3188.080 1247.210 3198.895 ;
        RECT 1246.390 3153.650 1247.990 3188.080 ;
        RECT 1246.390 3150.690 1248.130 3153.650 ;
        RECT 1246.390 3149.510 1248.570 3150.690 ;
        RECT 1246.390 3126.450 1247.990 3149.510 ;
        RECT 1246.390 3088.750 1248.130 3126.450 ;
        RECT 1246.390 3075.890 1247.990 3088.750 ;
        RECT 1246.390 3074.710 1248.570 3075.890 ;
        RECT 1246.390 3064.950 1248.130 3074.710 ;
        RECT 1246.390 3045.290 1247.990 3064.950 ;
        RECT 1245.550 3044.110 1247.990 3045.290 ;
        RECT 1245.990 3041.450 1246.290 3044.110 ;
        RECT 1246.390 3041.450 1247.990 3044.110 ;
        RECT 1245.990 3041.150 1247.990 3041.450 ;
        RECT 1246.390 1848.050 1247.990 3041.150 ;
        RECT 1246.390 1738.950 1248.130 1848.050 ;
        RECT 1246.390 1715.450 1247.990 1738.950 ;
        RECT 1246.390 1712.490 1248.130 1715.450 ;
        RECT 1246.390 1711.310 1248.570 1712.490 ;
        RECT 1246.390 1710.640 1247.990 1711.310 ;
        RECT 1245.550 1707.910 1246.730 1709.090 ;
        RECT 1245.990 1661.050 1246.290 1707.910 ;
        RECT 1245.990 1660.750 1247.210 1661.050 ;
        RECT 1246.910 1538.665 1247.210 1660.750 ;
        RECT 1246.895 1538.335 1247.225 1538.665 ;
        RECT 1245.975 1490.735 1246.305 1491.065 ;
        RECT 1245.990 1449.585 1246.290 1490.735 ;
        RECT 1245.975 1449.255 1246.305 1449.585 ;
        RECT 1247.815 1447.895 1248.145 1448.225 ;
        RECT 1247.830 1409.450 1248.130 1447.895 ;
        RECT 1245.990 1409.150 1248.130 1409.450 ;
        RECT 1245.990 1399.265 1246.290 1409.150 ;
        RECT 1245.975 1398.935 1246.305 1399.265 ;
        RECT 1246.895 1352.695 1247.225 1353.025 ;
        RECT 1246.910 1352.345 1247.210 1352.695 ;
        RECT 1246.895 1352.015 1247.225 1352.345 ;
        RECT 1247.815 1303.055 1248.145 1303.385 ;
        RECT 1247.830 1256.450 1248.130 1303.055 ;
        RECT 1246.910 1256.150 1248.130 1256.450 ;
        RECT 1246.910 1255.785 1247.210 1256.150 ;
        RECT 1246.895 1255.455 1247.225 1255.785 ;
        RECT 1245.975 1207.855 1246.305 1208.185 ;
        RECT 1245.990 1159.905 1246.290 1207.855 ;
        RECT 1245.975 1159.575 1246.305 1159.905 ;
        RECT 1246.895 1159.575 1247.225 1159.905 ;
        RECT 1246.910 1111.625 1247.210 1159.575 ;
        RECT 1246.895 1111.295 1247.225 1111.625 ;
        RECT 1246.895 1072.535 1247.225 1072.865 ;
        RECT 1246.910 1032.050 1247.210 1072.535 ;
        RECT 1246.910 1031.750 1248.130 1032.050 ;
        RECT 1247.830 1000.105 1248.130 1031.750 ;
        RECT 1247.815 999.775 1248.145 1000.105 ;
        RECT 1247.815 927.695 1248.145 928.025 ;
        RECT 1247.830 896.745 1248.130 927.695 ;
        RECT 1247.815 896.415 1248.145 896.745 ;
        RECT 1247.815 848.815 1248.145 849.145 ;
        RECT 1247.830 835.545 1248.130 848.815 ;
        RECT 1247.815 835.215 1248.145 835.545 ;
        RECT 1247.815 834.535 1248.145 834.865 ;
        RECT 1247.830 804.250 1248.130 834.535 ;
        RECT 1247.830 803.950 1249.050 804.250 ;
        RECT 1248.750 772.985 1249.050 803.950 ;
        RECT 1248.735 772.655 1249.065 772.985 ;
        RECT 1248.735 771.975 1249.065 772.305 ;
        RECT 1248.750 724.705 1249.050 771.975 ;
        RECT 1246.895 724.375 1247.225 724.705 ;
        RECT 1248.735 724.375 1249.065 724.705 ;
        RECT 1246.910 669.625 1247.210 724.375 ;
        RECT 1883.535 672.695 1883.865 673.025 ;
        RECT 1524.735 672.015 1525.065 672.345 ;
        RECT 1246.895 669.295 1247.225 669.625 ;
        RECT 1524.750 668.945 1525.050 672.015 ;
        RECT 1883.550 671.665 1883.850 672.695 ;
        RECT 1835.695 671.335 1836.025 671.665 ;
        RECT 1883.535 671.335 1883.865 671.665 ;
        RECT 1579.935 670.655 1580.265 670.985 ;
        RECT 1579.950 669.625 1580.250 670.655 ;
        RECT 1835.710 670.305 1836.010 671.335 ;
        RECT 2510.975 670.655 2511.305 670.985 ;
        RECT 1786.935 669.975 1787.265 670.305 ;
        RECT 1835.695 669.975 1836.025 670.305 ;
        RECT 2269.935 669.975 2270.265 670.305 ;
        RECT 2366.535 669.975 2366.865 670.305 ;
        RECT 1579.935 669.295 1580.265 669.625 ;
        RECT 1717.935 669.295 1718.265 669.625 ;
        RECT 1524.735 668.615 1525.065 668.945 ;
        RECT 1717.950 668.265 1718.250 669.295 ;
        RECT 1717.935 667.935 1718.265 668.265 ;
        RECT 1786.015 668.250 1786.345 668.265 ;
        RECT 1786.950 668.250 1787.250 669.975 ;
        RECT 2269.950 668.945 2270.250 669.975 ;
        RECT 2269.935 668.615 2270.265 668.945 ;
        RECT 2366.550 668.265 2366.850 669.975 ;
        RECT 2510.990 669.625 2511.290 670.655 ;
        RECT 2656.335 669.975 2656.665 670.305 ;
        RECT 2752.935 669.975 2753.265 670.305 ;
        RECT 2510.975 669.295 2511.305 669.625 ;
        RECT 2656.350 668.265 2656.650 669.975 ;
        RECT 2752.950 668.945 2753.250 669.975 ;
        RECT 2752.935 668.615 2753.265 668.945 ;
        RECT 1786.015 667.950 1787.250 668.250 ;
        RECT 1786.015 667.935 1786.345 667.950 ;
        RECT 2366.535 667.935 2366.865 668.265 ;
        RECT 2656.335 667.935 2656.665 668.265 ;
      LAYER via4 ;
        RECT 1247.390 3149.510 1248.570 3150.690 ;
        RECT 1246.470 3135.910 1247.650 3137.090 ;
        RECT 1246.470 3078.110 1247.650 3079.290 ;
        RECT 1247.390 3074.710 1248.570 3075.890 ;
        RECT 1246.470 3064.510 1247.650 3065.690 ;
        RECT 1247.390 1711.310 1248.570 1712.490 ;
      LAYER met5 ;
        RECT 1247.180 3149.300 1249.700 3150.900 ;
        RECT 1248.100 3137.300 1249.700 3149.300 ;
        RECT 1246.260 3135.700 1249.700 3137.300 ;
        RECT 1246.260 3077.900 1249.700 3079.500 ;
        RECT 1248.100 3076.100 1249.700 3077.900 ;
        RECT 1247.180 3074.500 1249.700 3076.100 ;
        RECT 1243.500 3064.300 1247.860 3065.900 ;
        RECT 1243.500 3045.500 1245.100 3064.300 ;
        RECT 1243.500 3043.900 1246.940 3045.500 ;
        RECT 1246.260 1711.100 1248.780 1712.700 ;
        RECT 1246.260 1709.300 1247.860 1711.100 ;
        RECT 1245.340 1707.700 1247.860 1709.300 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2317.110 3200.235 2317.390 3200.605 ;
        RECT 2317.180 3198.565 2317.320 3200.235 ;
        RECT 2317.110 3198.195 2317.390 3198.565 ;
        RECT 2350.690 3198.450 2350.970 3198.565 ;
        RECT 2352.460 3198.450 2352.740 3200.000 ;
        RECT 2350.690 3198.310 2352.740 3198.450 ;
        RECT 2350.690 3198.195 2350.970 3198.310 ;
        RECT 2352.460 3197.600 2352.740 3198.310 ;
      LAYER via2 ;
        RECT 2317.110 3200.280 2317.390 3200.560 ;
        RECT 2317.110 3198.240 2317.390 3198.520 ;
        RECT 2350.690 3198.240 2350.970 3198.520 ;
      LAYER met3 ;
        RECT 1631.430 3200.570 1631.810 3200.580 ;
        RECT 1682.030 3200.570 1682.410 3200.580 ;
        RECT 1631.430 3200.270 1682.410 3200.570 ;
        RECT 1631.430 3200.260 1631.810 3200.270 ;
        RECT 1682.030 3200.260 1682.410 3200.270 ;
        RECT 2017.830 3200.570 2018.210 3200.580 ;
        RECT 2066.590 3200.570 2066.970 3200.580 ;
        RECT 2017.830 3200.270 2066.970 3200.570 ;
        RECT 2017.830 3200.260 2018.210 3200.270 ;
        RECT 2066.590 3200.260 2066.970 3200.270 ;
        RECT 2283.710 3200.570 2284.090 3200.580 ;
        RECT 2317.085 3200.570 2317.415 3200.585 ;
        RECT 2283.710 3200.270 2317.415 3200.570 ;
        RECT 2283.710 3200.260 2284.090 3200.270 ;
        RECT 2317.085 3200.255 2317.415 3200.270 ;
        RECT 1164.990 3199.890 1165.370 3199.900 ;
        RECT 1197.190 3199.890 1197.570 3199.900 ;
        RECT 1164.990 3199.590 1197.570 3199.890 ;
        RECT 1164.990 3199.580 1165.370 3199.590 ;
        RECT 1197.190 3199.580 1197.570 3199.590 ;
        RECT 1258.830 3199.890 1259.210 3199.900 ;
        RECT 1289.190 3199.890 1289.570 3199.900 ;
        RECT 1258.830 3199.590 1289.570 3199.890 ;
        RECT 1258.830 3199.580 1259.210 3199.590 ;
        RECT 1289.190 3199.580 1289.570 3199.590 ;
        RECT 1435.470 3199.890 1435.850 3199.900 ;
        RECT 1486.990 3199.890 1487.370 3199.900 ;
        RECT 1435.470 3199.590 1487.370 3199.890 ;
        RECT 1435.470 3199.580 1435.850 3199.590 ;
        RECT 1486.990 3199.580 1487.370 3199.590 ;
        RECT 1532.990 3199.890 1533.370 3199.900 ;
        RECT 1583.590 3199.890 1583.970 3199.900 ;
        RECT 1532.990 3199.590 1583.970 3199.890 ;
        RECT 1532.990 3199.580 1533.370 3199.590 ;
        RECT 1583.590 3199.580 1583.970 3199.590 ;
        RECT 1728.030 3199.890 1728.410 3199.900 ;
        RECT 1861.430 3199.890 1861.810 3199.900 ;
        RECT 1728.030 3199.590 1861.810 3199.890 ;
        RECT 1728.030 3199.580 1728.410 3199.590 ;
        RECT 1861.430 3199.580 1861.810 3199.590 ;
        RECT 1921.230 3199.890 1921.610 3199.900 ;
        RECT 1965.390 3199.890 1965.770 3199.900 ;
        RECT 1921.230 3199.590 1965.770 3199.890 ;
        RECT 1921.230 3199.580 1921.610 3199.590 ;
        RECT 1965.390 3199.580 1965.770 3199.590 ;
        RECT 2208.270 3199.890 2208.650 3199.900 ;
        RECT 2259.790 3199.890 2260.170 3199.900 ;
        RECT 2208.270 3199.590 2260.170 3199.890 ;
        RECT 2208.270 3199.580 2208.650 3199.590 ;
        RECT 2259.790 3199.580 2260.170 3199.590 ;
        RECT 1338.870 3199.210 1339.250 3199.220 ;
        RECT 1411.550 3199.210 1411.930 3199.220 ;
        RECT 1338.870 3198.910 1411.930 3199.210 ;
        RECT 1338.870 3198.900 1339.250 3198.910 ;
        RECT 1411.550 3198.900 1411.930 3198.910 ;
        RECT 2317.085 3198.530 2317.415 3198.545 ;
        RECT 2350.665 3198.530 2350.995 3198.545 ;
        RECT 2317.085 3198.230 2350.995 3198.530 ;
        RECT 2317.085 3198.215 2317.415 3198.230 ;
        RECT 2350.665 3198.215 2350.995 3198.230 ;
        RECT 1197.190 3197.170 1197.570 3197.180 ;
        RECT 1258.830 3197.170 1259.210 3197.180 ;
        RECT 1197.190 3196.870 1259.210 3197.170 ;
        RECT 1197.190 3196.860 1197.570 3196.870 ;
        RECT 1258.830 3196.860 1259.210 3196.870 ;
        RECT 1289.190 3197.170 1289.570 3197.180 ;
        RECT 1338.870 3197.170 1339.250 3197.180 ;
        RECT 1289.190 3196.870 1339.250 3197.170 ;
        RECT 1289.190 3196.860 1289.570 3196.870 ;
        RECT 1338.870 3196.860 1339.250 3196.870 ;
        RECT 1411.550 3197.170 1411.930 3197.180 ;
        RECT 1435.470 3197.170 1435.850 3197.180 ;
        RECT 1411.550 3196.870 1435.850 3197.170 ;
        RECT 1411.550 3196.860 1411.930 3196.870 ;
        RECT 1435.470 3196.860 1435.850 3196.870 ;
        RECT 1486.990 3197.170 1487.370 3197.180 ;
        RECT 1532.990 3197.170 1533.370 3197.180 ;
        RECT 1486.990 3196.870 1533.370 3197.170 ;
        RECT 1486.990 3196.860 1487.370 3196.870 ;
        RECT 1532.990 3196.860 1533.370 3196.870 ;
        RECT 1583.590 3197.170 1583.970 3197.180 ;
        RECT 1631.430 3197.170 1631.810 3197.180 ;
        RECT 1583.590 3196.870 1631.810 3197.170 ;
        RECT 1583.590 3196.860 1583.970 3196.870 ;
        RECT 1631.430 3196.860 1631.810 3196.870 ;
        RECT 1682.030 3197.170 1682.410 3197.180 ;
        RECT 1728.030 3197.170 1728.410 3197.180 ;
        RECT 1682.030 3196.870 1728.410 3197.170 ;
        RECT 1682.030 3196.860 1682.410 3196.870 ;
        RECT 1728.030 3196.860 1728.410 3196.870 ;
        RECT 1861.430 3197.170 1861.810 3197.180 ;
        RECT 1921.230 3197.170 1921.610 3197.180 ;
        RECT 1861.430 3196.870 1921.610 3197.170 ;
        RECT 1861.430 3196.860 1861.810 3196.870 ;
        RECT 1921.230 3196.860 1921.610 3196.870 ;
        RECT 1965.390 3197.170 1965.770 3197.180 ;
        RECT 2017.830 3197.170 2018.210 3197.180 ;
        RECT 1965.390 3196.870 2018.210 3197.170 ;
        RECT 1965.390 3196.860 1965.770 3196.870 ;
        RECT 2017.830 3196.860 2018.210 3196.870 ;
        RECT 2066.590 3197.170 2066.970 3197.180 ;
        RECT 2208.270 3197.170 2208.650 3197.180 ;
        RECT 2066.590 3196.870 2208.650 3197.170 ;
        RECT 2066.590 3196.860 2066.970 3196.870 ;
        RECT 2208.270 3196.860 2208.650 3196.870 ;
        RECT 2259.790 3197.170 2260.170 3197.180 ;
        RECT 2283.710 3197.170 2284.090 3197.180 ;
        RECT 2259.790 3196.870 2284.090 3197.170 ;
        RECT 2259.790 3196.860 2260.170 3196.870 ;
        RECT 2283.710 3196.860 2284.090 3196.870 ;
        RECT 1164.990 1545.450 1165.370 1545.460 ;
        RECT 3.070 1545.150 1165.370 1545.450 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 3.070 1544.090 3.370 1545.150 ;
        RECT 1164.990 1545.140 1165.370 1545.150 ;
        RECT -4.800 1543.790 3.370 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
      LAYER via3 ;
        RECT 1631.460 3200.260 1631.780 3200.580 ;
        RECT 1682.060 3200.260 1682.380 3200.580 ;
        RECT 2017.860 3200.260 2018.180 3200.580 ;
        RECT 2066.620 3200.260 2066.940 3200.580 ;
        RECT 2283.740 3200.260 2284.060 3200.580 ;
        RECT 1165.020 3199.580 1165.340 3199.900 ;
        RECT 1197.220 3199.580 1197.540 3199.900 ;
        RECT 1258.860 3199.580 1259.180 3199.900 ;
        RECT 1289.220 3199.580 1289.540 3199.900 ;
        RECT 1435.500 3199.580 1435.820 3199.900 ;
        RECT 1487.020 3199.580 1487.340 3199.900 ;
        RECT 1533.020 3199.580 1533.340 3199.900 ;
        RECT 1583.620 3199.580 1583.940 3199.900 ;
        RECT 1728.060 3199.580 1728.380 3199.900 ;
        RECT 1861.460 3199.580 1861.780 3199.900 ;
        RECT 1921.260 3199.580 1921.580 3199.900 ;
        RECT 1965.420 3199.580 1965.740 3199.900 ;
        RECT 2208.300 3199.580 2208.620 3199.900 ;
        RECT 2259.820 3199.580 2260.140 3199.900 ;
        RECT 1338.900 3198.900 1339.220 3199.220 ;
        RECT 1411.580 3198.900 1411.900 3199.220 ;
        RECT 1197.220 3196.860 1197.540 3197.180 ;
        RECT 1258.860 3196.860 1259.180 3197.180 ;
        RECT 1289.220 3196.860 1289.540 3197.180 ;
        RECT 1338.900 3196.860 1339.220 3197.180 ;
        RECT 1411.580 3196.860 1411.900 3197.180 ;
        RECT 1435.500 3196.860 1435.820 3197.180 ;
        RECT 1487.020 3196.860 1487.340 3197.180 ;
        RECT 1533.020 3196.860 1533.340 3197.180 ;
        RECT 1583.620 3196.860 1583.940 3197.180 ;
        RECT 1631.460 3196.860 1631.780 3197.180 ;
        RECT 1682.060 3196.860 1682.380 3197.180 ;
        RECT 1728.060 3196.860 1728.380 3197.180 ;
        RECT 1861.460 3196.860 1861.780 3197.180 ;
        RECT 1921.260 3196.860 1921.580 3197.180 ;
        RECT 1965.420 3196.860 1965.740 3197.180 ;
        RECT 2017.860 3196.860 2018.180 3197.180 ;
        RECT 2066.620 3196.860 2066.940 3197.180 ;
        RECT 2208.300 3196.860 2208.620 3197.180 ;
        RECT 2259.820 3196.860 2260.140 3197.180 ;
        RECT 2283.740 3196.860 2284.060 3197.180 ;
        RECT 1165.020 1545.140 1165.340 1545.460 ;
      LAYER met4 ;
        RECT 1631.455 3200.255 1631.785 3200.585 ;
        RECT 1682.055 3200.255 1682.385 3200.585 ;
        RECT 2017.855 3200.255 2018.185 3200.585 ;
        RECT 2066.615 3200.255 2066.945 3200.585 ;
        RECT 2283.735 3200.255 2284.065 3200.585 ;
        RECT 1165.015 3199.575 1165.345 3199.905 ;
        RECT 1197.215 3199.575 1197.545 3199.905 ;
        RECT 1258.855 3199.575 1259.185 3199.905 ;
        RECT 1289.215 3199.575 1289.545 3199.905 ;
        RECT 1435.495 3199.575 1435.825 3199.905 ;
        RECT 1487.015 3199.575 1487.345 3199.905 ;
        RECT 1533.015 3199.575 1533.345 3199.905 ;
        RECT 1583.615 3199.575 1583.945 3199.905 ;
        RECT 1165.030 1545.465 1165.330 3199.575 ;
        RECT 1197.230 3197.185 1197.530 3199.575 ;
        RECT 1258.870 3197.185 1259.170 3199.575 ;
        RECT 1289.230 3197.185 1289.530 3199.575 ;
        RECT 1338.895 3198.895 1339.225 3199.225 ;
        RECT 1411.575 3198.895 1411.905 3199.225 ;
        RECT 1338.910 3197.185 1339.210 3198.895 ;
        RECT 1411.590 3197.185 1411.890 3198.895 ;
        RECT 1435.510 3197.185 1435.810 3199.575 ;
        RECT 1487.030 3197.185 1487.330 3199.575 ;
        RECT 1533.030 3197.185 1533.330 3199.575 ;
        RECT 1583.630 3197.185 1583.930 3199.575 ;
        RECT 1631.470 3197.185 1631.770 3200.255 ;
        RECT 1682.070 3197.185 1682.370 3200.255 ;
        RECT 1728.055 3199.575 1728.385 3199.905 ;
        RECT 1861.455 3199.575 1861.785 3199.905 ;
        RECT 1921.255 3199.575 1921.585 3199.905 ;
        RECT 1965.415 3199.575 1965.745 3199.905 ;
        RECT 1728.070 3197.185 1728.370 3199.575 ;
        RECT 1861.470 3197.185 1861.770 3199.575 ;
        RECT 1921.270 3197.185 1921.570 3199.575 ;
        RECT 1965.430 3197.185 1965.730 3199.575 ;
        RECT 2017.870 3197.185 2018.170 3200.255 ;
        RECT 2066.630 3197.185 2066.930 3200.255 ;
        RECT 2208.295 3199.575 2208.625 3199.905 ;
        RECT 2259.815 3199.575 2260.145 3199.905 ;
        RECT 2208.310 3197.185 2208.610 3199.575 ;
        RECT 2259.830 3197.185 2260.130 3199.575 ;
        RECT 2283.750 3197.185 2284.050 3200.255 ;
        RECT 1197.215 3196.855 1197.545 3197.185 ;
        RECT 1258.855 3196.855 1259.185 3197.185 ;
        RECT 1289.215 3196.855 1289.545 3197.185 ;
        RECT 1338.895 3196.855 1339.225 3197.185 ;
        RECT 1411.575 3196.855 1411.905 3197.185 ;
        RECT 1435.495 3196.855 1435.825 3197.185 ;
        RECT 1487.015 3196.855 1487.345 3197.185 ;
        RECT 1533.015 3196.855 1533.345 3197.185 ;
        RECT 1583.615 3196.855 1583.945 3197.185 ;
        RECT 1631.455 3196.855 1631.785 3197.185 ;
        RECT 1682.055 3196.855 1682.385 3197.185 ;
        RECT 1728.055 3196.855 1728.385 3197.185 ;
        RECT 1861.455 3196.855 1861.785 3197.185 ;
        RECT 1921.255 3196.855 1921.585 3197.185 ;
        RECT 1965.415 3196.855 1965.745 3197.185 ;
        RECT 2017.855 3196.855 2018.185 3197.185 ;
        RECT 2066.615 3196.855 2066.945 3197.185 ;
        RECT 2208.295 3196.855 2208.625 3197.185 ;
        RECT 2259.815 3196.855 2260.145 3197.185 ;
        RECT 2283.735 3196.855 2284.065 3197.185 ;
        RECT 1165.015 1545.135 1165.345 1545.465 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1148.690 3199.980 1149.010 3200.040 ;
        RECT 2390.230 3199.980 2390.550 3200.040 ;
        RECT 1148.690 3199.840 2390.550 3199.980 ;
        RECT 1148.690 3199.780 1149.010 3199.840 ;
        RECT 2390.230 3199.780 2390.550 3199.840 ;
        RECT 16.630 1331.680 16.950 1331.740 ;
        RECT 1148.690 1331.680 1149.010 1331.740 ;
        RECT 16.630 1331.540 1149.010 1331.680 ;
        RECT 16.630 1331.480 16.950 1331.540 ;
        RECT 1148.690 1331.480 1149.010 1331.540 ;
      LAYER via ;
        RECT 1148.720 3199.780 1148.980 3200.040 ;
        RECT 2390.260 3199.780 2390.520 3200.040 ;
        RECT 16.660 1331.480 16.920 1331.740 ;
        RECT 1148.720 1331.480 1148.980 1331.740 ;
      LAYER met2 ;
        RECT 1148.720 3199.750 1148.980 3200.070 ;
        RECT 2390.260 3199.810 2390.520 3200.070 ;
        RECT 2391.560 3199.810 2391.840 3200.000 ;
        RECT 2390.260 3199.750 2391.840 3199.810 ;
        RECT 1148.780 1331.770 1148.920 3199.750 ;
        RECT 2390.320 3199.670 2391.840 3199.750 ;
        RECT 2391.560 3197.600 2391.840 3199.670 ;
        RECT 16.660 1331.450 16.920 1331.770 ;
        RECT 1148.720 1331.450 1148.980 1331.770 ;
        RECT 16.720 1328.565 16.860 1331.450 ;
        RECT 16.650 1328.195 16.930 1328.565 ;
      LAYER via2 ;
        RECT 16.650 1328.240 16.930 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 16.625 1328.530 16.955 1328.545 ;
        RECT -4.800 1328.230 16.955 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 16.625 1328.215 16.955 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2041.625 3198.125 2042.715 3198.295 ;
      LAYER mcon ;
        RECT 2042.545 3198.125 2042.715 3198.295 ;
      LAYER met1 ;
        RECT 2234.290 3210.520 2234.610 3210.580 ;
        RECT 2431.170 3210.520 2431.490 3210.580 ;
        RECT 2234.290 3210.380 2431.490 3210.520 ;
        RECT 2234.290 3210.320 2234.610 3210.380 ;
        RECT 2431.170 3210.320 2431.490 3210.380 ;
        RECT 20.310 3198.280 20.630 3198.340 ;
        RECT 2041.565 3198.280 2041.855 3198.325 ;
        RECT 20.310 3198.140 2041.855 3198.280 ;
        RECT 20.310 3198.080 20.630 3198.140 ;
        RECT 2041.565 3198.095 2041.855 3198.140 ;
        RECT 2042.485 3198.280 2042.775 3198.325 ;
        RECT 2234.290 3198.280 2234.610 3198.340 ;
        RECT 2042.485 3198.140 2234.610 3198.280 ;
        RECT 2042.485 3198.095 2042.775 3198.140 ;
        RECT 2234.290 3198.080 2234.610 3198.140 ;
      LAYER via ;
        RECT 2234.320 3210.320 2234.580 3210.580 ;
        RECT 2431.200 3210.320 2431.460 3210.580 ;
        RECT 20.340 3198.080 20.600 3198.340 ;
        RECT 2234.320 3198.080 2234.580 3198.340 ;
      LAYER met2 ;
        RECT 2234.320 3210.290 2234.580 3210.610 ;
        RECT 2431.200 3210.290 2431.460 3210.610 ;
        RECT 2234.380 3198.370 2234.520 3210.290 ;
        RECT 2431.260 3200.000 2431.400 3210.290 ;
        RECT 20.340 3198.050 20.600 3198.370 ;
        RECT 2234.320 3198.050 2234.580 3198.370 ;
        RECT 20.400 1113.005 20.540 3198.050 ;
        RECT 2431.120 3197.600 2431.400 3200.000 ;
        RECT 20.330 1112.635 20.610 1113.005 ;
      LAYER via2 ;
        RECT 20.330 1112.680 20.610 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 20.305 1112.970 20.635 1112.985 ;
        RECT -4.800 1112.670 20.635 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 20.305 1112.655 20.635 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 897.500 14.190 897.560 ;
        RECT 24.450 897.500 24.770 897.560 ;
        RECT 13.870 897.360 24.770 897.500 ;
        RECT 13.870 897.300 14.190 897.360 ;
        RECT 24.450 897.300 24.770 897.360 ;
      LAYER via ;
        RECT 13.900 897.300 14.160 897.560 ;
        RECT 24.480 897.300 24.740 897.560 ;
      LAYER met2 ;
        RECT 24.470 3209.755 24.750 3210.125 ;
        RECT 2470.750 3209.755 2471.030 3210.125 ;
        RECT 24.540 897.590 24.680 3209.755 ;
        RECT 2470.820 3200.000 2470.960 3209.755 ;
        RECT 2470.680 3197.600 2470.960 3200.000 ;
        RECT 13.900 897.445 14.160 897.590 ;
        RECT 13.890 897.075 14.170 897.445 ;
        RECT 24.480 897.270 24.740 897.590 ;
      LAYER via2 ;
        RECT 24.470 3209.800 24.750 3210.080 ;
        RECT 2470.750 3209.800 2471.030 3210.080 ;
        RECT 13.890 897.120 14.170 897.400 ;
      LAYER met3 ;
        RECT 24.445 3210.090 24.775 3210.105 ;
        RECT 2470.725 3210.090 2471.055 3210.105 ;
        RECT 24.445 3209.790 2471.055 3210.090 ;
        RECT 24.445 3209.775 24.775 3209.790 ;
        RECT 2470.725 3209.775 2471.055 3209.790 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 13.865 897.410 14.195 897.425 ;
        RECT -4.800 897.110 14.195 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 13.865 897.095 14.195 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2314.790 3209.840 2315.110 3209.900 ;
        RECT 2510.290 3209.840 2510.610 3209.900 ;
        RECT 2314.790 3209.700 2510.610 3209.840 ;
        RECT 2314.790 3209.640 2315.110 3209.700 ;
        RECT 2510.290 3209.640 2510.610 3209.700 ;
      LAYER via ;
        RECT 2314.820 3209.640 2315.080 3209.900 ;
        RECT 2510.320 3209.640 2510.580 3209.900 ;
      LAYER met2 ;
        RECT 2314.820 3209.610 2315.080 3209.930 ;
        RECT 2510.320 3209.610 2510.580 3209.930 ;
        RECT 2314.880 3198.565 2315.020 3209.610 ;
        RECT 2510.380 3200.000 2510.520 3209.610 ;
        RECT 19.410 3198.195 19.690 3198.565 ;
        RECT 1703.930 3198.450 1704.210 3198.565 ;
        RECT 1704.850 3198.450 1705.130 3198.565 ;
        RECT 1703.930 3198.310 1705.130 3198.450 ;
        RECT 1703.930 3198.195 1704.210 3198.310 ;
        RECT 1704.850 3198.195 1705.130 3198.310 ;
        RECT 2314.810 3198.195 2315.090 3198.565 ;
        RECT 19.480 681.885 19.620 3198.195 ;
        RECT 2510.240 3197.600 2510.520 3200.000 ;
        RECT 19.410 681.515 19.690 681.885 ;
      LAYER via2 ;
        RECT 19.410 3198.240 19.690 3198.520 ;
        RECT 1703.930 3198.240 1704.210 3198.520 ;
        RECT 1704.850 3198.240 1705.130 3198.520 ;
        RECT 2314.810 3198.240 2315.090 3198.520 ;
        RECT 19.410 681.560 19.690 681.840 ;
      LAYER met3 ;
        RECT 19.385 3198.530 19.715 3198.545 ;
        RECT 1703.905 3198.530 1704.235 3198.545 ;
        RECT 19.385 3198.230 1704.235 3198.530 ;
        RECT 19.385 3198.215 19.715 3198.230 ;
        RECT 1703.905 3198.215 1704.235 3198.230 ;
        RECT 1704.825 3198.530 1705.155 3198.545 ;
        RECT 2314.785 3198.530 2315.115 3198.545 ;
        RECT 1704.825 3198.230 2315.115 3198.530 ;
        RECT 1704.825 3198.215 1705.155 3198.230 ;
        RECT 2314.785 3198.215 2315.115 3198.230 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 19.385 681.850 19.715 681.865 ;
        RECT -4.800 681.550 19.715 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 19.385 681.535 19.715 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 3209.075 18.770 3209.445 ;
        RECT 2549.870 3209.075 2550.150 3209.445 ;
        RECT 18.560 466.325 18.700 3209.075 ;
        RECT 2549.940 3200.000 2550.080 3209.075 ;
        RECT 2549.800 3197.600 2550.080 3200.000 ;
        RECT 18.490 465.955 18.770 466.325 ;
      LAYER via2 ;
        RECT 18.490 3209.120 18.770 3209.400 ;
        RECT 2549.870 3209.120 2550.150 3209.400 ;
        RECT 18.490 466.000 18.770 466.280 ;
      LAYER met3 ;
        RECT 18.465 3209.410 18.795 3209.425 ;
        RECT 2549.845 3209.410 2550.175 3209.425 ;
        RECT 18.465 3209.110 2550.175 3209.410 ;
        RECT 18.465 3209.095 18.795 3209.110 ;
        RECT 2549.845 3209.095 2550.175 3209.110 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 18.465 466.290 18.795 466.305 ;
        RECT -4.800 465.990 18.795 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 18.465 465.975 18.795 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2425.650 3209.160 2425.970 3209.220 ;
        RECT 2588.950 3209.160 2589.270 3209.220 ;
        RECT 2425.650 3209.020 2589.270 3209.160 ;
        RECT 2425.650 3208.960 2425.970 3209.020 ;
        RECT 2588.950 3208.960 2589.270 3209.020 ;
        RECT 1104.530 3199.640 1104.850 3199.700 ;
        RECT 1176.290 3199.640 1176.610 3199.700 ;
        RECT 1104.530 3199.500 1176.610 3199.640 ;
        RECT 1104.530 3199.440 1104.850 3199.500 ;
        RECT 1176.290 3199.440 1176.610 3199.500 ;
        RECT 27.670 3197.600 27.990 3197.660 ;
        RECT 116.450 3197.600 116.770 3197.660 ;
        RECT 27.670 3197.460 116.770 3197.600 ;
        RECT 27.670 3197.400 27.990 3197.460 ;
        RECT 116.450 3197.400 116.770 3197.460 ;
        RECT 781.610 3197.600 781.930 3197.660 ;
        RECT 813.350 3197.600 813.670 3197.660 ;
        RECT 781.610 3197.460 813.670 3197.600 ;
        RECT 781.610 3197.400 781.930 3197.460 ;
        RECT 813.350 3197.400 813.670 3197.460 ;
        RECT 1007.470 3197.600 1007.790 3197.660 ;
        RECT 1055.310 3197.600 1055.630 3197.660 ;
        RECT 1007.470 3197.460 1055.630 3197.600 ;
        RECT 1007.470 3197.400 1007.790 3197.460 ;
        RECT 1055.310 3197.400 1055.630 3197.460 ;
        RECT 303.210 3196.240 303.530 3196.300 ;
        RECT 330.810 3196.240 331.130 3196.300 ;
        RECT 303.210 3196.100 331.130 3196.240 ;
        RECT 303.210 3196.040 303.530 3196.100 ;
        RECT 330.810 3196.040 331.130 3196.100 ;
      LAYER via ;
        RECT 2425.680 3208.960 2425.940 3209.220 ;
        RECT 2588.980 3208.960 2589.240 3209.220 ;
        RECT 1104.560 3199.440 1104.820 3199.700 ;
        RECT 1176.320 3199.440 1176.580 3199.700 ;
        RECT 27.700 3197.400 27.960 3197.660 ;
        RECT 116.480 3197.400 116.740 3197.660 ;
        RECT 781.640 3197.400 781.900 3197.660 ;
        RECT 813.380 3197.400 813.640 3197.660 ;
        RECT 1007.500 3197.400 1007.760 3197.660 ;
        RECT 1055.340 3197.400 1055.600 3197.660 ;
        RECT 303.240 3196.040 303.500 3196.300 ;
        RECT 330.840 3196.040 331.100 3196.300 ;
      LAYER met2 ;
        RECT 2425.680 3208.930 2425.940 3209.250 ;
        RECT 2588.980 3208.930 2589.240 3209.250 ;
        RECT 1104.560 3199.410 1104.820 3199.730 ;
        RECT 1176.320 3199.410 1176.580 3199.730 ;
        RECT 2316.190 3199.555 2316.470 3199.925 ;
        RECT 2355.290 3199.555 2355.570 3199.925 ;
        RECT 548.410 3198.875 548.690 3199.245 ;
        RECT 596.710 3198.875 596.990 3199.245 ;
        RECT 814.290 3198.875 814.570 3199.245 ;
        RECT 886.510 3198.875 886.790 3199.245 ;
        RECT 17.110 3197.515 17.390 3197.885 ;
        RECT 27.690 3197.515 27.970 3197.885 ;
        RECT 116.930 3197.770 117.210 3197.885 ;
        RECT 116.540 3197.690 117.210 3197.770 ;
        RECT 116.480 3197.630 117.210 3197.690 ;
        RECT 17.180 250.765 17.320 3197.515 ;
        RECT 27.700 3197.370 27.960 3197.515 ;
        RECT 116.480 3197.370 116.740 3197.630 ;
        RECT 116.930 3197.515 117.210 3197.630 ;
        RECT 254.010 3197.090 254.290 3197.205 ;
        RECT 255.390 3197.090 255.670 3197.205 ;
        RECT 254.010 3196.950 255.670 3197.090 ;
        RECT 254.010 3196.835 254.290 3196.950 ;
        RECT 255.390 3196.835 255.670 3196.950 ;
        RECT 303.230 3196.835 303.510 3197.205 ;
        RECT 350.610 3197.090 350.890 3197.205 ;
        RECT 351.990 3197.090 352.270 3197.205 ;
        RECT 350.610 3196.950 352.270 3197.090 ;
        RECT 350.610 3196.835 350.890 3196.950 ;
        RECT 351.990 3196.835 352.270 3196.950 ;
        RECT 399.830 3197.090 400.110 3197.205 ;
        RECT 400.750 3197.090 401.030 3197.205 ;
        RECT 399.830 3196.950 401.030 3197.090 ;
        RECT 399.830 3196.835 400.110 3196.950 ;
        RECT 400.750 3196.835 401.030 3196.950 ;
        RECT 447.210 3197.090 447.490 3197.205 ;
        RECT 448.590 3197.090 448.870 3197.205 ;
        RECT 447.210 3196.950 448.870 3197.090 ;
        RECT 447.210 3196.835 447.490 3196.950 ;
        RECT 448.590 3196.835 448.870 3196.950 ;
        RECT 303.300 3196.330 303.440 3196.835 ;
        RECT 548.480 3196.525 548.620 3198.875 ;
        RECT 596.780 3197.205 596.920 3198.875 ;
        RECT 738.850 3197.770 739.130 3197.885 ;
        RECT 738.000 3197.630 739.130 3197.770 ;
        RECT 738.000 3197.205 738.140 3197.630 ;
        RECT 738.850 3197.515 739.130 3197.630 ;
        RECT 781.630 3197.515 781.910 3197.885 ;
        RECT 781.640 3197.370 781.900 3197.515 ;
        RECT 813.380 3197.370 813.640 3197.690 ;
        RECT 596.710 3196.835 596.990 3197.205 ;
        RECT 737.930 3196.835 738.210 3197.205 ;
        RECT 813.440 3197.090 813.580 3197.370 ;
        RECT 814.360 3197.090 814.500 3198.875 ;
        RECT 886.580 3197.205 886.720 3198.875 ;
        RECT 931.590 3197.515 931.870 3197.885 ;
        RECT 813.440 3196.950 814.500 3197.090 ;
        RECT 886.510 3196.835 886.790 3197.205 ;
        RECT 930.210 3197.090 930.490 3197.205 ;
        RECT 931.660 3197.090 931.800 3197.515 ;
        RECT 1007.500 3197.370 1007.760 3197.690 ;
        RECT 1055.340 3197.370 1055.600 3197.690 ;
        RECT 1104.090 3197.515 1104.370 3197.885 ;
        RECT 1007.560 3197.205 1007.700 3197.370 ;
        RECT 930.210 3196.950 931.800 3197.090 ;
        RECT 930.210 3196.835 930.490 3196.950 ;
        RECT 1007.490 3196.835 1007.770 3197.205 ;
        RECT 1055.400 3196.525 1055.540 3197.370 ;
        RECT 1104.160 3197.090 1104.300 3197.515 ;
        RECT 1104.620 3197.090 1104.760 3199.410 ;
        RECT 1176.380 3199.245 1176.520 3199.410 ;
        RECT 1176.310 3198.875 1176.590 3199.245 ;
        RECT 2316.260 3198.565 2316.400 3199.555 ;
        RECT 2355.360 3198.565 2355.500 3199.555 ;
        RECT 2425.740 3198.565 2425.880 3208.930 ;
        RECT 2589.040 3200.000 2589.180 3208.930 ;
        RECT 2316.190 3198.195 2316.470 3198.565 ;
        RECT 2355.290 3198.195 2355.570 3198.565 ;
        RECT 2425.670 3198.195 2425.950 3198.565 ;
        RECT 2588.900 3197.600 2589.180 3200.000 ;
        RECT 1104.160 3196.950 1104.760 3197.090 ;
        RECT 303.240 3196.010 303.500 3196.330 ;
        RECT 330.830 3196.155 331.110 3196.525 ;
        RECT 548.410 3196.155 548.690 3196.525 ;
        RECT 1055.330 3196.155 1055.610 3196.525 ;
        RECT 330.840 3196.010 331.100 3196.155 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 2316.190 3199.600 2316.470 3199.880 ;
        RECT 2355.290 3199.600 2355.570 3199.880 ;
        RECT 548.410 3198.920 548.690 3199.200 ;
        RECT 596.710 3198.920 596.990 3199.200 ;
        RECT 814.290 3198.920 814.570 3199.200 ;
        RECT 886.510 3198.920 886.790 3199.200 ;
        RECT 17.110 3197.560 17.390 3197.840 ;
        RECT 27.690 3197.560 27.970 3197.840 ;
        RECT 116.930 3197.560 117.210 3197.840 ;
        RECT 254.010 3196.880 254.290 3197.160 ;
        RECT 255.390 3196.880 255.670 3197.160 ;
        RECT 303.230 3196.880 303.510 3197.160 ;
        RECT 350.610 3196.880 350.890 3197.160 ;
        RECT 351.990 3196.880 352.270 3197.160 ;
        RECT 399.830 3196.880 400.110 3197.160 ;
        RECT 400.750 3196.880 401.030 3197.160 ;
        RECT 447.210 3196.880 447.490 3197.160 ;
        RECT 448.590 3196.880 448.870 3197.160 ;
        RECT 738.850 3197.560 739.130 3197.840 ;
        RECT 781.630 3197.560 781.910 3197.840 ;
        RECT 596.710 3196.880 596.990 3197.160 ;
        RECT 737.930 3196.880 738.210 3197.160 ;
        RECT 931.590 3197.560 931.870 3197.840 ;
        RECT 886.510 3196.880 886.790 3197.160 ;
        RECT 930.210 3196.880 930.490 3197.160 ;
        RECT 1104.090 3197.560 1104.370 3197.840 ;
        RECT 1007.490 3196.880 1007.770 3197.160 ;
        RECT 1176.310 3198.920 1176.590 3199.200 ;
        RECT 2316.190 3198.240 2316.470 3198.520 ;
        RECT 2355.290 3198.240 2355.570 3198.520 ;
        RECT 2425.670 3198.240 2425.950 3198.520 ;
        RECT 330.830 3196.200 331.110 3196.480 ;
        RECT 548.410 3196.200 548.690 3196.480 ;
        RECT 1055.330 3196.200 1055.610 3196.480 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 1728.950 3200.570 1729.330 3200.580 ;
        RECT 1703.230 3200.270 1729.330 3200.570 ;
        RECT 1676.510 3199.890 1676.890 3199.900 ;
        RECT 1703.230 3199.890 1703.530 3200.270 ;
        RECT 1728.950 3200.260 1729.330 3200.270 ;
        RECT 1676.510 3199.590 1703.530 3199.890 ;
        RECT 2316.165 3199.890 2316.495 3199.905 ;
        RECT 2355.265 3199.890 2355.595 3199.905 ;
        RECT 2316.165 3199.590 2355.595 3199.890 ;
        RECT 1676.510 3199.580 1676.890 3199.590 ;
        RECT 2316.165 3199.575 2316.495 3199.590 ;
        RECT 2355.265 3199.575 2355.595 3199.590 ;
        RECT 548.385 3199.210 548.715 3199.225 ;
        RECT 596.685 3199.210 597.015 3199.225 ;
        RECT 548.385 3198.910 597.015 3199.210 ;
        RECT 548.385 3198.895 548.715 3198.910 ;
        RECT 596.685 3198.895 597.015 3198.910 ;
        RECT 814.265 3199.210 814.595 3199.225 ;
        RECT 886.485 3199.210 886.815 3199.225 ;
        RECT 814.265 3198.910 886.815 3199.210 ;
        RECT 814.265 3198.895 814.595 3198.910 ;
        RECT 886.485 3198.895 886.815 3198.910 ;
        RECT 1176.285 3199.210 1176.615 3199.225 ;
        RECT 1177.870 3199.210 1178.250 3199.220 ;
        RECT 1176.285 3198.910 1178.250 3199.210 ;
        RECT 1176.285 3198.895 1176.615 3198.910 ;
        RECT 1177.870 3198.900 1178.250 3198.910 ;
        RECT 2316.165 3198.530 2316.495 3198.545 ;
        RECT 2315.950 3198.215 2316.495 3198.530 ;
        RECT 2355.265 3198.530 2355.595 3198.545 ;
        RECT 2425.645 3198.530 2425.975 3198.545 ;
        RECT 2355.265 3198.215 2355.810 3198.530 ;
        RECT 17.085 3197.850 17.415 3197.865 ;
        RECT 27.665 3197.850 27.995 3197.865 ;
        RECT 17.085 3197.550 27.995 3197.850 ;
        RECT 17.085 3197.535 17.415 3197.550 ;
        RECT 27.665 3197.535 27.995 3197.550 ;
        RECT 116.905 3197.850 117.235 3197.865 ;
        RECT 164.950 3197.850 165.330 3197.860 ;
        RECT 165.870 3197.850 166.250 3197.860 ;
        RECT 116.905 3197.535 117.450 3197.850 ;
        RECT 164.950 3197.550 166.250 3197.850 ;
        RECT 164.950 3197.540 165.330 3197.550 ;
        RECT 165.870 3197.540 166.250 3197.550 ;
        RECT 738.825 3197.850 739.155 3197.865 ;
        RECT 781.605 3197.850 781.935 3197.865 ;
        RECT 738.825 3197.550 781.935 3197.850 ;
        RECT 738.825 3197.535 739.155 3197.550 ;
        RECT 781.605 3197.535 781.935 3197.550 ;
        RECT 931.565 3197.850 931.895 3197.865 ;
        RECT 1104.065 3197.850 1104.395 3197.865 ;
        RECT 931.565 3197.550 990.530 3197.850 ;
        RECT 931.565 3197.535 931.895 3197.550 ;
        RECT 117.150 3196.490 117.450 3197.535 ;
        RECT 165.870 3197.170 166.250 3197.180 ;
        RECT 253.985 3197.170 254.315 3197.185 ;
        RECT 165.870 3196.870 254.315 3197.170 ;
        RECT 165.870 3196.860 166.250 3196.870 ;
        RECT 253.985 3196.855 254.315 3196.870 ;
        RECT 255.365 3197.170 255.695 3197.185 ;
        RECT 303.205 3197.170 303.535 3197.185 ;
        RECT 350.585 3197.170 350.915 3197.185 ;
        RECT 255.365 3196.870 303.535 3197.170 ;
        RECT 255.365 3196.855 255.695 3196.870 ;
        RECT 303.205 3196.855 303.535 3196.870 ;
        RECT 330.590 3196.870 350.915 3197.170 ;
        RECT 330.590 3196.505 330.890 3196.870 ;
        RECT 350.585 3196.855 350.915 3196.870 ;
        RECT 351.965 3197.170 352.295 3197.185 ;
        RECT 399.805 3197.170 400.135 3197.185 ;
        RECT 351.965 3196.870 400.135 3197.170 ;
        RECT 351.965 3196.855 352.295 3196.870 ;
        RECT 399.805 3196.855 400.135 3196.870 ;
        RECT 400.725 3197.170 401.055 3197.185 ;
        RECT 447.185 3197.170 447.515 3197.185 ;
        RECT 400.725 3196.870 447.515 3197.170 ;
        RECT 400.725 3196.855 401.055 3196.870 ;
        RECT 447.185 3196.855 447.515 3196.870 ;
        RECT 448.565 3197.170 448.895 3197.185 ;
        RECT 596.685 3197.170 597.015 3197.185 ;
        RECT 737.905 3197.170 738.235 3197.185 ;
        RECT 448.565 3196.870 496.490 3197.170 ;
        RECT 448.565 3196.855 448.895 3196.870 ;
        RECT 164.950 3196.490 165.330 3196.500 ;
        RECT 117.150 3196.190 165.330 3196.490 ;
        RECT 330.590 3196.190 331.135 3196.505 ;
        RECT 496.190 3196.490 496.490 3196.870 ;
        RECT 596.685 3196.870 738.235 3197.170 ;
        RECT 596.685 3196.855 597.015 3196.870 ;
        RECT 737.905 3196.855 738.235 3196.870 ;
        RECT 886.485 3197.170 886.815 3197.185 ;
        RECT 930.185 3197.170 930.515 3197.185 ;
        RECT 886.485 3196.870 930.515 3197.170 ;
        RECT 990.230 3197.170 990.530 3197.550 ;
        RECT 1061.990 3197.550 1104.395 3197.850 ;
        RECT 1007.465 3197.170 1007.795 3197.185 ;
        RECT 990.230 3196.870 1007.795 3197.170 ;
        RECT 886.485 3196.855 886.815 3196.870 ;
        RECT 930.185 3196.855 930.515 3196.870 ;
        RECT 1007.465 3196.855 1007.795 3196.870 ;
        RECT 548.385 3196.490 548.715 3196.505 ;
        RECT 496.190 3196.190 548.715 3196.490 ;
        RECT 164.950 3196.180 165.330 3196.190 ;
        RECT 330.805 3196.175 331.135 3196.190 ;
        RECT 548.385 3196.175 548.715 3196.190 ;
        RECT 1055.305 3196.490 1055.635 3196.505 ;
        RECT 1061.990 3196.490 1062.290 3197.550 ;
        RECT 1104.065 3197.535 1104.395 3197.550 ;
        RECT 1177.870 3197.850 1178.250 3197.860 ;
        RECT 1245.030 3197.850 1245.410 3197.860 ;
        RECT 2315.950 3197.850 2316.250 3198.215 ;
        RECT 1177.870 3197.550 1245.410 3197.850 ;
        RECT 1177.870 3197.540 1178.250 3197.550 ;
        RECT 1245.030 3197.540 1245.410 3197.550 ;
        RECT 1288.310 3197.550 1340.130 3197.850 ;
        RECT 1288.310 3197.170 1288.610 3197.550 ;
        RECT 1259.790 3196.870 1288.610 3197.170 ;
        RECT 1339.830 3197.170 1340.130 3197.550 ;
        RECT 1385.830 3197.550 1436.730 3197.850 ;
        RECT 1385.830 3197.170 1386.130 3197.550 ;
        RECT 1339.830 3196.870 1386.130 3197.170 ;
        RECT 1436.430 3197.170 1436.730 3197.550 ;
        RECT 1486.110 3197.550 1535.170 3197.850 ;
        RECT 1486.110 3197.170 1486.410 3197.550 ;
        RECT 1436.430 3196.870 1486.410 3197.170 ;
        RECT 1534.870 3197.170 1535.170 3197.550 ;
        RECT 1582.710 3197.550 1632.690 3197.850 ;
        RECT 1582.710 3197.170 1583.010 3197.550 ;
        RECT 1534.870 3196.870 1583.010 3197.170 ;
        RECT 1632.390 3197.170 1632.690 3197.550 ;
        RECT 1859.630 3197.550 1922.490 3197.850 ;
        RECT 1676.510 3197.170 1676.890 3197.180 ;
        RECT 1632.390 3196.870 1676.890 3197.170 ;
        RECT 1055.305 3196.190 1062.290 3196.490 ;
        RECT 1245.030 3196.490 1245.410 3196.500 ;
        RECT 1259.790 3196.490 1260.090 3196.870 ;
        RECT 1676.510 3196.860 1676.890 3196.870 ;
        RECT 1728.950 3197.170 1729.330 3197.180 ;
        RECT 1859.630 3197.170 1859.930 3197.550 ;
        RECT 1728.950 3196.870 1859.930 3197.170 ;
        RECT 1922.190 3197.170 1922.490 3197.550 ;
        RECT 1964.510 3197.550 2209.530 3197.850 ;
        RECT 1964.510 3197.170 1964.810 3197.550 ;
        RECT 1922.190 3196.870 1964.810 3197.170 ;
        RECT 2209.230 3197.170 2209.530 3197.550 ;
        RECT 2258.910 3197.550 2316.250 3197.850 ;
        RECT 2355.510 3197.850 2355.810 3198.215 ;
        RECT 2403.350 3198.230 2425.975 3198.530 ;
        RECT 2403.350 3197.850 2403.650 3198.230 ;
        RECT 2425.645 3198.215 2425.975 3198.230 ;
        RECT 2355.510 3197.550 2403.650 3197.850 ;
        RECT 2258.910 3197.170 2259.210 3197.550 ;
        RECT 2209.230 3196.870 2259.210 3197.170 ;
        RECT 1728.950 3196.860 1729.330 3196.870 ;
        RECT 1245.030 3196.190 1260.090 3196.490 ;
        RECT 1055.305 3196.175 1055.635 3196.190 ;
        RECT 1245.030 3196.180 1245.410 3196.190 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
      LAYER via3 ;
        RECT 1676.540 3199.580 1676.860 3199.900 ;
        RECT 1728.980 3200.260 1729.300 3200.580 ;
        RECT 1177.900 3198.900 1178.220 3199.220 ;
        RECT 164.980 3197.540 165.300 3197.860 ;
        RECT 165.900 3197.540 166.220 3197.860 ;
        RECT 165.900 3196.860 166.220 3197.180 ;
        RECT 164.980 3196.180 165.300 3196.500 ;
        RECT 1177.900 3197.540 1178.220 3197.860 ;
        RECT 1245.060 3197.540 1245.380 3197.860 ;
        RECT 1245.060 3196.180 1245.380 3196.500 ;
        RECT 1676.540 3196.860 1676.860 3197.180 ;
        RECT 1728.980 3196.860 1729.300 3197.180 ;
      LAYER met4 ;
        RECT 1728.975 3200.255 1729.305 3200.585 ;
        RECT 1676.535 3199.575 1676.865 3199.905 ;
        RECT 1177.895 3198.895 1178.225 3199.225 ;
        RECT 1177.910 3197.865 1178.210 3198.895 ;
        RECT 164.975 3197.535 165.305 3197.865 ;
        RECT 165.895 3197.535 166.225 3197.865 ;
        RECT 1177.895 3197.535 1178.225 3197.865 ;
        RECT 1245.055 3197.535 1245.385 3197.865 ;
        RECT 164.990 3196.505 165.290 3197.535 ;
        RECT 165.910 3197.185 166.210 3197.535 ;
        RECT 165.895 3196.855 166.225 3197.185 ;
        RECT 1245.070 3196.505 1245.370 3197.535 ;
        RECT 1676.550 3197.185 1676.850 3199.575 ;
        RECT 1728.990 3197.185 1729.290 3200.255 ;
        RECT 1676.535 3196.855 1676.865 3197.185 ;
        RECT 1728.975 3196.855 1729.305 3197.185 ;
        RECT 164.975 3196.175 165.305 3196.505 ;
        RECT 1245.055 3196.175 1245.385 3196.505 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2579.310 3208.395 2579.590 3208.765 ;
        RECT 2628.530 3208.395 2628.810 3208.765 ;
        RECT 208.010 3207.715 208.290 3208.085 ;
        RECT 265.510 3207.715 265.790 3208.085 ;
        RECT 304.610 3207.715 304.890 3208.085 ;
        RECT 342.330 3207.715 342.610 3208.085 ;
        RECT 458.710 3207.715 458.990 3208.085 ;
        RECT 497.810 3207.715 498.090 3208.085 ;
        RECT 594.410 3207.715 594.690 3208.085 ;
        RECT 651.910 3207.715 652.190 3208.085 ;
        RECT 730.570 3207.715 730.850 3208.085 ;
        RECT 787.610 3207.715 787.890 3208.085 ;
        RECT 884.210 3207.715 884.490 3208.085 ;
        RECT 941.710 3207.715 941.990 3208.085 ;
        RECT 969.770 3207.715 970.050 3208.085 ;
        RECT 1038.310 3207.715 1038.590 3208.085 ;
        RECT 1217.710 3207.715 1217.990 3208.085 ;
        RECT 1376.410 3207.715 1376.690 3208.085 ;
        RECT 208.080 3204.685 208.220 3207.715 ;
        RECT 265.580 3204.685 265.720 3207.715 ;
        RECT 304.680 3204.685 304.820 3207.715 ;
        RECT 342.400 3204.685 342.540 3207.715 ;
        RECT 458.780 3204.685 458.920 3207.715 ;
        RECT 497.880 3204.685 498.020 3207.715 ;
        RECT 594.480 3204.685 594.620 3207.715 ;
        RECT 651.980 3204.685 652.120 3207.715 ;
        RECT 730.640 3204.685 730.780 3207.715 ;
        RECT 787.680 3204.685 787.820 3207.715 ;
        RECT 884.280 3204.685 884.420 3207.715 ;
        RECT 941.780 3204.685 941.920 3207.715 ;
        RECT 969.840 3204.685 969.980 3207.715 ;
        RECT 1038.380 3204.685 1038.520 3207.715 ;
        RECT 1217.780 3204.685 1217.920 3207.715 ;
        RECT 1376.480 3204.685 1376.620 3207.715 ;
        RECT 208.010 3204.315 208.290 3204.685 ;
        RECT 265.510 3204.315 265.790 3204.685 ;
        RECT 304.610 3204.315 304.890 3204.685 ;
        RECT 342.330 3204.315 342.610 3204.685 ;
        RECT 458.710 3204.315 458.990 3204.685 ;
        RECT 497.810 3204.315 498.090 3204.685 ;
        RECT 594.410 3204.315 594.690 3204.685 ;
        RECT 651.910 3204.315 652.190 3204.685 ;
        RECT 730.570 3204.315 730.850 3204.685 ;
        RECT 787.610 3204.315 787.890 3204.685 ;
        RECT 884.210 3204.315 884.490 3204.685 ;
        RECT 941.710 3204.315 941.990 3204.685 ;
        RECT 969.770 3204.315 970.050 3204.685 ;
        RECT 1038.310 3204.315 1038.590 3204.685 ;
        RECT 1217.710 3204.315 1217.990 3204.685 ;
        RECT 1376.410 3204.315 1376.690 3204.685 ;
        RECT 2579.380 3201.285 2579.520 3208.395 ;
        RECT 2579.310 3200.915 2579.590 3201.285 ;
        RECT 2628.600 3200.000 2628.740 3208.395 ;
        RECT 20.790 3198.875 21.070 3199.245 ;
        RECT 20.330 35.770 20.610 35.885 ;
        RECT 20.860 35.770 21.000 3198.875 ;
        RECT 2628.460 3197.600 2628.740 3200.000 ;
        RECT 20.330 35.630 21.000 35.770 ;
        RECT 20.330 35.515 20.610 35.630 ;
      LAYER via2 ;
        RECT 2579.310 3208.440 2579.590 3208.720 ;
        RECT 2628.530 3208.440 2628.810 3208.720 ;
        RECT 208.010 3207.760 208.290 3208.040 ;
        RECT 265.510 3207.760 265.790 3208.040 ;
        RECT 304.610 3207.760 304.890 3208.040 ;
        RECT 342.330 3207.760 342.610 3208.040 ;
        RECT 458.710 3207.760 458.990 3208.040 ;
        RECT 497.810 3207.760 498.090 3208.040 ;
        RECT 594.410 3207.760 594.690 3208.040 ;
        RECT 651.910 3207.760 652.190 3208.040 ;
        RECT 730.570 3207.760 730.850 3208.040 ;
        RECT 787.610 3207.760 787.890 3208.040 ;
        RECT 884.210 3207.760 884.490 3208.040 ;
        RECT 941.710 3207.760 941.990 3208.040 ;
        RECT 969.770 3207.760 970.050 3208.040 ;
        RECT 1038.310 3207.760 1038.590 3208.040 ;
        RECT 1217.710 3207.760 1217.990 3208.040 ;
        RECT 1376.410 3207.760 1376.690 3208.040 ;
        RECT 208.010 3204.360 208.290 3204.640 ;
        RECT 265.510 3204.360 265.790 3204.640 ;
        RECT 304.610 3204.360 304.890 3204.640 ;
        RECT 342.330 3204.360 342.610 3204.640 ;
        RECT 458.710 3204.360 458.990 3204.640 ;
        RECT 497.810 3204.360 498.090 3204.640 ;
        RECT 594.410 3204.360 594.690 3204.640 ;
        RECT 651.910 3204.360 652.190 3204.640 ;
        RECT 730.570 3204.360 730.850 3204.640 ;
        RECT 787.610 3204.360 787.890 3204.640 ;
        RECT 884.210 3204.360 884.490 3204.640 ;
        RECT 941.710 3204.360 941.990 3204.640 ;
        RECT 969.770 3204.360 970.050 3204.640 ;
        RECT 1038.310 3204.360 1038.590 3204.640 ;
        RECT 1217.710 3204.360 1217.990 3204.640 ;
        RECT 1376.410 3204.360 1376.690 3204.640 ;
        RECT 2579.310 3200.960 2579.590 3201.240 ;
        RECT 20.790 3198.920 21.070 3199.200 ;
        RECT 20.330 35.560 20.610 35.840 ;
      LAYER met3 ;
        RECT 2579.285 3208.730 2579.615 3208.745 ;
        RECT 2628.505 3208.730 2628.835 3208.745 ;
        RECT 2579.285 3208.430 2628.835 3208.730 ;
        RECT 2579.285 3208.415 2579.615 3208.430 ;
        RECT 2628.505 3208.415 2628.835 3208.430 ;
        RECT 37.070 3208.050 37.450 3208.060 ;
        RECT 64.670 3208.050 65.050 3208.060 ;
        RECT 37.070 3207.750 65.050 3208.050 ;
        RECT 37.070 3207.740 37.450 3207.750 ;
        RECT 64.670 3207.740 65.050 3207.750 ;
        RECT 138.270 3208.050 138.650 3208.060 ;
        RECT 207.985 3208.050 208.315 3208.065 ;
        RECT 138.270 3207.750 208.315 3208.050 ;
        RECT 138.270 3207.740 138.650 3207.750 ;
        RECT 207.985 3207.735 208.315 3207.750 ;
        RECT 265.485 3208.050 265.815 3208.065 ;
        RECT 304.585 3208.050 304.915 3208.065 ;
        RECT 265.485 3207.750 304.915 3208.050 ;
        RECT 265.485 3207.735 265.815 3207.750 ;
        RECT 304.585 3207.735 304.915 3207.750 ;
        RECT 342.305 3208.050 342.635 3208.065 ;
        RECT 398.630 3208.050 399.010 3208.060 ;
        RECT 342.305 3207.750 399.010 3208.050 ;
        RECT 342.305 3207.735 342.635 3207.750 ;
        RECT 398.630 3207.740 399.010 3207.750 ;
        RECT 458.685 3208.050 459.015 3208.065 ;
        RECT 497.785 3208.050 498.115 3208.065 ;
        RECT 458.685 3207.750 498.115 3208.050 ;
        RECT 458.685 3207.735 459.015 3207.750 ;
        RECT 497.785 3207.735 498.115 3207.750 ;
        RECT 548.590 3208.050 548.970 3208.060 ;
        RECT 594.385 3208.050 594.715 3208.065 ;
        RECT 548.590 3207.750 594.715 3208.050 ;
        RECT 548.590 3207.740 548.970 3207.750 ;
        RECT 594.385 3207.735 594.715 3207.750 ;
        RECT 651.885 3208.050 652.215 3208.065 ;
        RECT 686.590 3208.050 686.970 3208.060 ;
        RECT 651.885 3207.750 686.970 3208.050 ;
        RECT 651.885 3207.735 652.215 3207.750 ;
        RECT 686.590 3207.740 686.970 3207.750 ;
        RECT 730.545 3208.050 730.875 3208.065 ;
        RECT 787.585 3208.050 787.915 3208.065 ;
        RECT 730.545 3207.750 787.915 3208.050 ;
        RECT 730.545 3207.735 730.875 3207.750 ;
        RECT 787.585 3207.735 787.915 3207.750 ;
        RECT 836.550 3208.050 836.930 3208.060 ;
        RECT 884.185 3208.050 884.515 3208.065 ;
        RECT 836.550 3207.750 884.515 3208.050 ;
        RECT 836.550 3207.740 836.930 3207.750 ;
        RECT 884.185 3207.735 884.515 3207.750 ;
        RECT 941.685 3208.050 942.015 3208.065 ;
        RECT 969.745 3208.050 970.075 3208.065 ;
        RECT 941.685 3207.750 970.075 3208.050 ;
        RECT 941.685 3207.735 942.015 3207.750 ;
        RECT 969.745 3207.735 970.075 3207.750 ;
        RECT 1038.285 3208.050 1038.615 3208.065 ;
        RECT 1075.750 3208.050 1076.130 3208.060 ;
        RECT 1038.285 3207.750 1076.130 3208.050 ;
        RECT 1038.285 3207.735 1038.615 3207.750 ;
        RECT 1075.750 3207.740 1076.130 3207.750 ;
        RECT 1110.710 3208.050 1111.090 3208.060 ;
        RECT 1130.030 3208.050 1130.410 3208.060 ;
        RECT 1110.710 3207.750 1130.410 3208.050 ;
        RECT 1110.710 3207.740 1111.090 3207.750 ;
        RECT 1130.030 3207.740 1130.410 3207.750 ;
        RECT 1159.470 3208.050 1159.850 3208.060 ;
        RECT 1217.685 3208.050 1218.015 3208.065 ;
        RECT 1159.470 3207.750 1218.015 3208.050 ;
        RECT 1159.470 3207.740 1159.850 3207.750 ;
        RECT 1217.685 3207.735 1218.015 3207.750 ;
        RECT 1376.385 3208.050 1376.715 3208.065 ;
        RECT 1413.390 3208.050 1413.770 3208.060 ;
        RECT 1376.385 3207.750 1413.770 3208.050 ;
        RECT 1376.385 3207.735 1376.715 3207.750 ;
        RECT 1413.390 3207.740 1413.770 3207.750 ;
        RECT 1508.150 3208.050 1508.530 3208.060 ;
        RECT 1514.590 3208.050 1514.970 3208.060 ;
        RECT 1508.150 3207.750 1514.970 3208.050 ;
        RECT 1508.150 3207.740 1508.530 3207.750 ;
        RECT 1514.590 3207.740 1514.970 3207.750 ;
        RECT 1546.790 3208.050 1547.170 3208.060 ;
        RECT 1591.870 3208.050 1592.250 3208.060 ;
        RECT 1546.790 3207.750 1592.250 3208.050 ;
        RECT 1546.790 3207.740 1547.170 3207.750 ;
        RECT 1591.870 3207.740 1592.250 3207.750 ;
        RECT 1635.110 3208.050 1635.490 3208.060 ;
        RECT 1682.950 3208.050 1683.330 3208.060 ;
        RECT 1635.110 3207.750 1683.330 3208.050 ;
        RECT 1635.110 3207.740 1635.490 3207.750 ;
        RECT 1682.950 3207.740 1683.330 3207.750 ;
        RECT 1741.830 3208.050 1742.210 3208.060 ;
        RECT 1755.630 3208.050 1756.010 3208.060 ;
        RECT 1741.830 3207.750 1756.010 3208.050 ;
        RECT 1741.830 3207.740 1742.210 3207.750 ;
        RECT 1755.630 3207.740 1756.010 3207.750 ;
        RECT 1883.510 3208.050 1883.890 3208.060 ;
        RECT 1898.230 3208.050 1898.610 3208.060 ;
        RECT 1883.510 3207.750 1898.610 3208.050 ;
        RECT 1883.510 3207.740 1883.890 3207.750 ;
        RECT 1898.230 3207.740 1898.610 3207.750 ;
        RECT 2118.110 3208.050 2118.490 3208.060 ;
        RECT 2162.270 3208.050 2162.650 3208.060 ;
        RECT 2118.110 3207.750 2162.650 3208.050 ;
        RECT 2118.110 3207.740 2118.490 3207.750 ;
        RECT 2162.270 3207.740 2162.650 3207.750 ;
        RECT 2269.910 3208.050 2270.290 3208.060 ;
        RECT 2317.750 3208.050 2318.130 3208.060 ;
        RECT 2269.910 3207.750 2318.130 3208.050 ;
        RECT 2269.910 3207.740 2270.290 3207.750 ;
        RECT 2317.750 3207.740 2318.130 3207.750 ;
        RECT 207.985 3204.650 208.315 3204.665 ;
        RECT 265.485 3204.650 265.815 3204.665 ;
        RECT 207.985 3204.350 265.815 3204.650 ;
        RECT 207.985 3204.335 208.315 3204.350 ;
        RECT 265.485 3204.335 265.815 3204.350 ;
        RECT 304.585 3204.650 304.915 3204.665 ;
        RECT 342.305 3204.650 342.635 3204.665 ;
        RECT 304.585 3204.350 342.635 3204.650 ;
        RECT 304.585 3204.335 304.915 3204.350 ;
        RECT 342.305 3204.335 342.635 3204.350 ;
        RECT 404.150 3204.650 404.530 3204.660 ;
        RECT 458.685 3204.650 459.015 3204.665 ;
        RECT 404.150 3204.350 459.015 3204.650 ;
        RECT 404.150 3204.340 404.530 3204.350 ;
        RECT 458.685 3204.335 459.015 3204.350 ;
        RECT 497.785 3204.650 498.115 3204.665 ;
        RECT 542.150 3204.650 542.530 3204.660 ;
        RECT 497.785 3204.350 542.530 3204.650 ;
        RECT 497.785 3204.335 498.115 3204.350 ;
        RECT 542.150 3204.340 542.530 3204.350 ;
        RECT 594.385 3204.650 594.715 3204.665 ;
        RECT 651.885 3204.650 652.215 3204.665 ;
        RECT 594.385 3204.350 652.215 3204.650 ;
        RECT 594.385 3204.335 594.715 3204.350 ;
        RECT 651.885 3204.335 652.215 3204.350 ;
        RECT 692.110 3204.650 692.490 3204.660 ;
        RECT 730.545 3204.650 730.875 3204.665 ;
        RECT 692.110 3204.350 730.875 3204.650 ;
        RECT 692.110 3204.340 692.490 3204.350 ;
        RECT 730.545 3204.335 730.875 3204.350 ;
        RECT 787.585 3204.650 787.915 3204.665 ;
        RECT 830.110 3204.650 830.490 3204.660 ;
        RECT 787.585 3204.350 830.490 3204.650 ;
        RECT 787.585 3204.335 787.915 3204.350 ;
        RECT 830.110 3204.340 830.490 3204.350 ;
        RECT 884.185 3204.650 884.515 3204.665 ;
        RECT 941.685 3204.650 942.015 3204.665 ;
        RECT 884.185 3204.350 942.015 3204.650 ;
        RECT 884.185 3204.335 884.515 3204.350 ;
        RECT 941.685 3204.335 942.015 3204.350 ;
        RECT 969.745 3204.650 970.075 3204.665 ;
        RECT 1038.285 3204.650 1038.615 3204.665 ;
        RECT 969.745 3204.350 1038.615 3204.650 ;
        RECT 969.745 3204.335 970.075 3204.350 ;
        RECT 1038.285 3204.335 1038.615 3204.350 ;
        RECT 1217.685 3204.650 1218.015 3204.665 ;
        RECT 1258.830 3204.650 1259.210 3204.660 ;
        RECT 1217.685 3204.350 1259.210 3204.650 ;
        RECT 1217.685 3204.335 1218.015 3204.350 ;
        RECT 1258.830 3204.340 1259.210 3204.350 ;
        RECT 1322.310 3204.650 1322.690 3204.660 ;
        RECT 1376.385 3204.650 1376.715 3204.665 ;
        RECT 1322.310 3204.350 1376.715 3204.650 ;
        RECT 1322.310 3204.340 1322.690 3204.350 ;
        RECT 1376.385 3204.335 1376.715 3204.350 ;
        RECT 1449.270 3204.650 1449.650 3204.660 ;
        RECT 1496.190 3204.650 1496.570 3204.660 ;
        RECT 1449.270 3204.350 1496.570 3204.650 ;
        RECT 1449.270 3204.340 1449.650 3204.350 ;
        RECT 1496.190 3204.340 1496.570 3204.350 ;
        RECT 1593.710 3204.650 1594.090 3204.660 ;
        RECT 1610.270 3204.650 1610.650 3204.660 ;
        RECT 1593.710 3204.350 1610.650 3204.650 ;
        RECT 1593.710 3204.340 1594.090 3204.350 ;
        RECT 1610.270 3204.340 1610.650 3204.350 ;
        RECT 1786.910 3204.650 1787.290 3204.660 ;
        RECT 1834.750 3204.650 1835.130 3204.660 ;
        RECT 1786.910 3204.350 1835.130 3204.650 ;
        RECT 1786.910 3204.340 1787.290 3204.350 ;
        RECT 1834.750 3204.340 1835.130 3204.350 ;
        RECT 1835.670 3204.650 1836.050 3204.660 ;
        RECT 1882.590 3204.650 1882.970 3204.660 ;
        RECT 1835.670 3204.350 1882.970 3204.650 ;
        RECT 1835.670 3204.340 1836.050 3204.350 ;
        RECT 1882.590 3204.340 1882.970 3204.350 ;
        RECT 1945.150 3204.650 1945.530 3204.660 ;
        RECT 1978.270 3204.650 1978.650 3204.660 ;
        RECT 1945.150 3204.350 1978.650 3204.650 ;
        RECT 1945.150 3204.340 1945.530 3204.350 ;
        RECT 1978.270 3204.340 1978.650 3204.350 ;
        RECT 1980.110 3204.650 1980.490 3204.660 ;
        RECT 1996.670 3204.650 1997.050 3204.660 ;
        RECT 1980.110 3204.350 1997.050 3204.650 ;
        RECT 1980.110 3204.340 1980.490 3204.350 ;
        RECT 1996.670 3204.340 1997.050 3204.350 ;
        RECT 2180.670 3204.650 2181.050 3204.660 ;
        RECT 2192.630 3204.650 2193.010 3204.660 ;
        RECT 2180.670 3204.350 2193.010 3204.650 ;
        RECT 2180.670 3204.340 2181.050 3204.350 ;
        RECT 2192.630 3204.340 2193.010 3204.350 ;
        RECT 2319.590 3201.250 2319.970 3201.260 ;
        RECT 2404.230 3201.250 2404.610 3201.260 ;
        RECT 2319.590 3200.950 2404.610 3201.250 ;
        RECT 2319.590 3200.940 2319.970 3200.950 ;
        RECT 2404.230 3200.940 2404.610 3200.950 ;
        RECT 2545.910 3201.250 2546.290 3201.260 ;
        RECT 2579.285 3201.250 2579.615 3201.265 ;
        RECT 2545.910 3200.950 2579.615 3201.250 ;
        RECT 2545.910 3200.940 2546.290 3200.950 ;
        RECT 2579.285 3200.935 2579.615 3200.950 ;
        RECT 20.765 3199.210 21.095 3199.225 ;
        RECT 26.950 3199.210 27.330 3199.220 ;
        RECT 20.765 3198.910 27.330 3199.210 ;
        RECT 20.765 3198.895 21.095 3198.910 ;
        RECT 26.950 3198.900 27.330 3198.910 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 20.305 35.850 20.635 35.865 ;
        RECT -4.800 35.550 20.635 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 20.305 35.535 20.635 35.550 ;
      LAYER via3 ;
        RECT 37.100 3207.740 37.420 3208.060 ;
        RECT 64.700 3207.740 65.020 3208.060 ;
        RECT 138.300 3207.740 138.620 3208.060 ;
        RECT 398.660 3207.740 398.980 3208.060 ;
        RECT 548.620 3207.740 548.940 3208.060 ;
        RECT 686.620 3207.740 686.940 3208.060 ;
        RECT 836.580 3207.740 836.900 3208.060 ;
        RECT 1075.780 3207.740 1076.100 3208.060 ;
        RECT 1110.740 3207.740 1111.060 3208.060 ;
        RECT 1130.060 3207.740 1130.380 3208.060 ;
        RECT 1159.500 3207.740 1159.820 3208.060 ;
        RECT 1413.420 3207.740 1413.740 3208.060 ;
        RECT 1508.180 3207.740 1508.500 3208.060 ;
        RECT 1514.620 3207.740 1514.940 3208.060 ;
        RECT 1546.820 3207.740 1547.140 3208.060 ;
        RECT 1591.900 3207.740 1592.220 3208.060 ;
        RECT 1635.140 3207.740 1635.460 3208.060 ;
        RECT 1682.980 3207.740 1683.300 3208.060 ;
        RECT 1741.860 3207.740 1742.180 3208.060 ;
        RECT 1755.660 3207.740 1755.980 3208.060 ;
        RECT 1883.540 3207.740 1883.860 3208.060 ;
        RECT 1898.260 3207.740 1898.580 3208.060 ;
        RECT 2118.140 3207.740 2118.460 3208.060 ;
        RECT 2162.300 3207.740 2162.620 3208.060 ;
        RECT 2269.940 3207.740 2270.260 3208.060 ;
        RECT 2317.780 3207.740 2318.100 3208.060 ;
        RECT 404.180 3204.340 404.500 3204.660 ;
        RECT 542.180 3204.340 542.500 3204.660 ;
        RECT 692.140 3204.340 692.460 3204.660 ;
        RECT 830.140 3204.340 830.460 3204.660 ;
        RECT 1258.860 3204.340 1259.180 3204.660 ;
        RECT 1322.340 3204.340 1322.660 3204.660 ;
        RECT 1449.300 3204.340 1449.620 3204.660 ;
        RECT 1496.220 3204.340 1496.540 3204.660 ;
        RECT 1593.740 3204.340 1594.060 3204.660 ;
        RECT 1610.300 3204.340 1610.620 3204.660 ;
        RECT 1786.940 3204.340 1787.260 3204.660 ;
        RECT 1834.780 3204.340 1835.100 3204.660 ;
        RECT 1835.700 3204.340 1836.020 3204.660 ;
        RECT 1882.620 3204.340 1882.940 3204.660 ;
        RECT 1945.180 3204.340 1945.500 3204.660 ;
        RECT 1978.300 3204.340 1978.620 3204.660 ;
        RECT 1980.140 3204.340 1980.460 3204.660 ;
        RECT 1996.700 3204.340 1997.020 3204.660 ;
        RECT 2180.700 3204.340 2181.020 3204.660 ;
        RECT 2192.660 3204.340 2192.980 3204.660 ;
        RECT 2319.620 3200.940 2319.940 3201.260 ;
        RECT 2404.260 3200.940 2404.580 3201.260 ;
        RECT 2545.940 3200.940 2546.260 3201.260 ;
        RECT 26.980 3198.900 27.300 3199.220 ;
      LAYER met4 ;
        RECT 26.550 3207.310 27.730 3208.490 ;
        RECT 36.670 3207.310 37.850 3208.490 ;
        RECT 64.695 3207.735 65.025 3208.065 ;
        RECT 26.990 3199.225 27.290 3207.310 ;
        RECT 64.710 3205.090 65.010 3207.735 ;
        RECT 137.870 3207.310 139.050 3208.490 ;
        RECT 398.230 3207.310 399.410 3208.490 ;
        RECT 403.750 3207.310 404.930 3208.490 ;
        RECT 548.615 3207.735 548.945 3208.065 ;
        RECT 64.270 3203.910 65.450 3205.090 ;
        RECT 404.190 3204.665 404.490 3207.310 ;
        RECT 548.630 3205.090 548.930 3207.735 ;
        RECT 686.190 3207.310 687.370 3208.490 ;
        RECT 691.710 3207.310 692.890 3208.490 ;
        RECT 836.575 3207.735 836.905 3208.065 ;
        RECT 404.175 3204.335 404.505 3204.665 ;
        RECT 541.750 3203.910 542.930 3205.090 ;
        RECT 548.190 3203.910 549.370 3205.090 ;
        RECT 692.150 3204.665 692.450 3207.310 ;
        RECT 836.590 3205.090 836.890 3207.735 ;
        RECT 1075.350 3207.310 1076.530 3208.490 ;
        RECT 1110.310 3207.310 1111.490 3208.490 ;
        RECT 1130.055 3207.735 1130.385 3208.065 ;
        RECT 1159.495 3207.735 1159.825 3208.065 ;
        RECT 1130.070 3205.090 1130.370 3207.735 ;
        RECT 1159.510 3205.090 1159.810 3207.735 ;
        RECT 1321.910 3207.310 1323.090 3208.490 ;
        RECT 1412.990 3207.310 1414.170 3208.490 ;
        RECT 1495.790 3207.310 1496.970 3208.490 ;
        RECT 1507.750 3207.310 1508.930 3208.490 ;
        RECT 1514.190 3207.310 1515.370 3208.490 ;
        RECT 1546.390 3207.310 1547.570 3208.490 ;
        RECT 1591.895 3207.735 1592.225 3208.065 ;
        RECT 692.135 3204.335 692.465 3204.665 ;
        RECT 829.710 3203.910 830.890 3205.090 ;
        RECT 836.150 3203.910 837.330 3205.090 ;
        RECT 1129.630 3203.910 1130.810 3205.090 ;
        RECT 1159.070 3203.910 1160.250 3205.090 ;
        RECT 1258.430 3203.910 1259.610 3205.090 ;
        RECT 1322.350 3204.665 1322.650 3207.310 ;
        RECT 1322.335 3204.335 1322.665 3204.665 ;
        RECT 1448.870 3203.910 1450.050 3205.090 ;
        RECT 1496.230 3204.665 1496.530 3207.310 ;
        RECT 1591.910 3205.090 1592.210 3207.735 ;
        RECT 1609.870 3207.310 1611.050 3208.490 ;
        RECT 1634.710 3207.310 1635.890 3208.490 ;
        RECT 1682.975 3207.735 1683.305 3208.065 ;
        RECT 1496.215 3204.335 1496.545 3204.665 ;
        RECT 1591.470 3203.910 1592.650 3205.090 ;
        RECT 1593.310 3203.910 1594.490 3205.090 ;
        RECT 1610.310 3204.665 1610.610 3207.310 ;
        RECT 1682.990 3205.090 1683.290 3207.735 ;
        RECT 1741.430 3207.310 1742.610 3208.490 ;
        RECT 1755.655 3207.735 1755.985 3208.065 ;
        RECT 1834.790 3207.750 1836.010 3208.050 ;
        RECT 1755.670 3205.090 1755.970 3207.735 ;
        RECT 1610.295 3204.335 1610.625 3204.665 ;
        RECT 1682.550 3203.910 1683.730 3205.090 ;
        RECT 1755.230 3203.910 1756.410 3205.090 ;
        RECT 1786.510 3203.910 1787.690 3205.090 ;
        RECT 1834.790 3204.665 1835.090 3207.750 ;
        RECT 1835.710 3204.665 1836.010 3207.750 ;
        RECT 1883.110 3207.310 1884.290 3208.490 ;
        RECT 1898.255 3207.735 1898.585 3208.065 ;
        RECT 1898.270 3205.090 1898.570 3207.735 ;
        RECT 2117.710 3207.310 2118.890 3208.490 ;
        RECT 2162.295 3207.735 2162.625 3208.065 ;
        RECT 2162.310 3205.090 2162.610 3207.735 ;
        RECT 2192.230 3207.310 2193.410 3208.490 ;
        RECT 2269.510 3207.310 2270.690 3208.490 ;
        RECT 2317.775 3207.735 2318.105 3208.065 ;
        RECT 1834.775 3204.335 1835.105 3204.665 ;
        RECT 1835.695 3204.335 1836.025 3204.665 ;
        RECT 1882.190 3203.910 1883.370 3205.090 ;
        RECT 1897.830 3203.910 1899.010 3205.090 ;
        RECT 1944.750 3203.910 1945.930 3205.090 ;
        RECT 1977.870 3203.910 1979.050 3205.090 ;
        RECT 1979.710 3203.910 1980.890 3205.090 ;
        RECT 1996.270 3203.910 1997.450 3205.090 ;
        RECT 2161.870 3203.910 2163.050 3205.090 ;
        RECT 2180.270 3203.910 2181.450 3205.090 ;
        RECT 2192.670 3204.665 2192.970 3207.310 ;
        RECT 2317.790 3205.090 2318.090 3207.735 ;
        RECT 2403.830 3207.310 2405.010 3208.490 ;
        RECT 2192.655 3204.335 2192.985 3204.665 ;
        RECT 2317.350 3203.910 2318.530 3205.090 ;
        RECT 2319.190 3203.910 2320.370 3205.090 ;
        RECT 2319.630 3201.265 2319.930 3203.910 ;
        RECT 2404.270 3201.265 2404.570 3207.310 ;
        RECT 2319.615 3200.935 2319.945 3201.265 ;
        RECT 2404.255 3200.935 2404.585 3201.265 ;
        RECT 2545.510 3200.510 2546.690 3201.690 ;
        RECT 26.975 3198.895 27.305 3199.225 ;
      LAYER met5 ;
        RECT 26.340 3207.100 38.060 3208.700 ;
        RECT 99.020 3207.100 139.260 3208.700 ;
        RECT 398.020 3207.100 405.140 3208.700 ;
        RECT 685.980 3207.100 693.100 3208.700 ;
        RECT 1075.140 3207.100 1111.700 3208.700 ;
        RECT 1315.260 3207.100 1323.300 3208.700 ;
        RECT 1412.000 3207.100 1415.300 3208.700 ;
        RECT 1495.580 3207.100 1509.140 3208.700 ;
        RECT 1513.980 3207.100 1547.780 3208.700 ;
        RECT 1609.660 3207.100 1636.100 3208.700 ;
        RECT 1704.420 3207.100 1742.820 3208.700 ;
        RECT 99.020 3205.300 100.620 3207.100 ;
        RECT 1315.260 3205.300 1316.860 3207.100 ;
        RECT 64.060 3203.700 100.620 3205.300 ;
        RECT 541.540 3203.700 549.580 3205.300 ;
        RECT 829.500 3203.700 837.540 3205.300 ;
        RECT 1129.420 3203.700 1160.460 3205.300 ;
        RECT 1258.220 3203.700 1316.860 3205.300 ;
        RECT 1413.700 3205.300 1415.300 3207.100 ;
        RECT 1413.700 3203.700 1450.260 3205.300 ;
        RECT 1591.260 3203.700 1594.700 3205.300 ;
        RECT 1682.340 3203.700 1701.420 3205.300 ;
        RECT 1699.820 3201.900 1701.420 3203.700 ;
        RECT 1704.420 3201.900 1706.020 3207.100 ;
        RECT 1882.900 3205.300 1884.500 3208.700 ;
        RECT 1930.740 3205.300 1933.260 3208.700 ;
        RECT 2088.980 3207.100 2119.100 3208.700 ;
        RECT 2192.020 3207.100 2224.900 3208.700 ;
        RECT 2088.980 3205.300 2090.580 3207.100 ;
        RECT 1755.020 3203.700 1787.900 3205.300 ;
        RECT 1881.980 3203.700 1884.500 3205.300 ;
        RECT 1897.620 3203.700 1946.140 3205.300 ;
        RECT 1977.660 3203.700 1981.100 3205.300 ;
        RECT 1996.060 3203.700 2090.580 3205.300 ;
        RECT 2161.660 3203.700 2181.660 3205.300 ;
        RECT 1699.820 3200.300 1706.020 3201.900 ;
        RECT 2223.300 3201.900 2224.900 3207.100 ;
        RECT 2267.460 3207.100 2270.900 3208.700 ;
        RECT 2403.620 3207.100 2478.820 3208.700 ;
        RECT 2267.460 3201.900 2269.060 3207.100 ;
        RECT 2477.220 3205.300 2478.820 3207.100 ;
        RECT 2317.140 3203.700 2320.580 3205.300 ;
        RECT 2477.220 3203.700 2546.900 3205.300 ;
        RECT 2223.300 3200.300 2269.060 3201.900 ;
        RECT 2545.300 3200.300 2546.900 3203.700 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1286.690 3211.880 1287.010 3211.940 ;
        RECT 2903.130 3211.880 2903.450 3211.940 ;
        RECT 1286.690 3211.740 2903.450 3211.880 ;
        RECT 1286.690 3211.680 1287.010 3211.740 ;
        RECT 2903.130 3211.680 2903.450 3211.740 ;
      LAYER via ;
        RECT 1286.720 3211.680 1286.980 3211.940 ;
        RECT 2903.160 3211.680 2903.420 3211.940 ;
      LAYER met2 ;
        RECT 1286.720 3211.650 1286.980 3211.970 ;
        RECT 2903.160 3211.650 2903.420 3211.970 ;
        RECT 1286.780 3200.000 1286.920 3211.650 ;
        RECT 1286.640 3197.600 1286.920 3200.000 ;
        RECT 2903.220 909.685 2903.360 3211.650 ;
        RECT 2903.150 909.315 2903.430 909.685 ;
      LAYER via2 ;
        RECT 2903.150 909.360 2903.430 909.640 ;
      LAYER met3 ;
        RECT 2903.125 909.650 2903.455 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2903.125 909.350 2924.800 909.650 ;
        RECT 2903.125 909.335 2903.455 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1325.790 3214.260 1326.110 3214.320 ;
        RECT 1604.090 3214.260 1604.410 3214.320 ;
        RECT 1325.790 3214.120 1604.410 3214.260 ;
        RECT 1325.790 3214.060 1326.110 3214.120 ;
        RECT 1604.090 3214.060 1604.410 3214.120 ;
        RECT 1604.090 3201.340 1604.410 3201.400 ;
        RECT 2903.590 3201.340 2903.910 3201.400 ;
        RECT 1604.090 3201.200 2903.910 3201.340 ;
        RECT 1604.090 3201.140 1604.410 3201.200 ;
        RECT 2903.590 3201.140 2903.910 3201.200 ;
      LAYER via ;
        RECT 1325.820 3214.060 1326.080 3214.320 ;
        RECT 1604.120 3214.060 1604.380 3214.320 ;
        RECT 1604.120 3201.140 1604.380 3201.400 ;
        RECT 2903.620 3201.140 2903.880 3201.400 ;
      LAYER met2 ;
        RECT 1325.820 3214.030 1326.080 3214.350 ;
        RECT 1604.120 3214.030 1604.380 3214.350 ;
        RECT 1325.880 3200.000 1326.020 3214.030 ;
        RECT 1604.180 3201.430 1604.320 3214.030 ;
        RECT 1604.120 3201.110 1604.380 3201.430 ;
        RECT 2903.620 3201.110 2903.880 3201.430 ;
        RECT 1325.740 3197.600 1326.020 3200.000 ;
        RECT 2903.680 1144.285 2903.820 3201.110 ;
        RECT 2903.610 1143.915 2903.890 1144.285 ;
      LAYER via2 ;
        RECT 2903.610 1143.960 2903.890 1144.240 ;
      LAYER met3 ;
        RECT 2903.585 1144.250 2903.915 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2903.585 1143.950 2924.800 1144.250 ;
        RECT 2903.585 1143.935 2903.915 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1365.810 3198.960 1366.130 3199.020 ;
        RECT 2904.050 3198.960 2904.370 3199.020 ;
        RECT 1365.810 3198.820 2904.370 3198.960 ;
        RECT 1365.810 3198.760 1366.130 3198.820 ;
        RECT 2904.050 3198.760 2904.370 3198.820 ;
      LAYER via ;
        RECT 1365.840 3198.760 1366.100 3199.020 ;
        RECT 2904.080 3198.760 2904.340 3199.020 ;
      LAYER met2 ;
        RECT 1365.300 3199.130 1365.580 3200.000 ;
        RECT 1365.300 3199.050 1366.040 3199.130 ;
        RECT 1365.300 3198.990 1366.100 3199.050 ;
        RECT 1365.300 3197.600 1365.580 3198.990 ;
        RECT 1365.840 3198.730 1366.100 3198.990 ;
        RECT 2904.080 3198.730 2904.340 3199.050 ;
        RECT 2904.140 1378.885 2904.280 3198.730 ;
        RECT 2904.070 1378.515 2904.350 1378.885 ;
      LAYER via2 ;
        RECT 2904.070 1378.560 2904.350 1378.840 ;
      LAYER met3 ;
        RECT 2904.045 1378.850 2904.375 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2904.045 1378.550 2924.800 1378.850 ;
        RECT 2904.045 1378.535 2904.375 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1406.290 3199.300 1406.610 3199.360 ;
        RECT 2654.270 3199.300 2654.590 3199.360 ;
        RECT 1406.290 3199.160 2654.590 3199.300 ;
        RECT 1406.290 3199.100 1406.610 3199.160 ;
        RECT 2654.270 3199.100 2654.590 3199.160 ;
        RECT 2654.270 1614.560 2654.590 1614.620 ;
        RECT 2900.370 1614.560 2900.690 1614.620 ;
        RECT 2654.270 1614.420 2900.690 1614.560 ;
        RECT 2654.270 1614.360 2654.590 1614.420 ;
        RECT 2900.370 1614.360 2900.690 1614.420 ;
      LAYER via ;
        RECT 1406.320 3199.100 1406.580 3199.360 ;
        RECT 2654.300 3199.100 2654.560 3199.360 ;
        RECT 2654.300 1614.360 2654.560 1614.620 ;
        RECT 2900.400 1614.360 2900.660 1614.620 ;
      LAYER met2 ;
        RECT 1404.860 3199.130 1405.140 3200.000 ;
        RECT 1406.320 3199.130 1406.580 3199.390 ;
        RECT 1404.860 3199.070 1406.580 3199.130 ;
        RECT 2654.300 3199.070 2654.560 3199.390 ;
        RECT 1404.860 3198.990 1406.520 3199.070 ;
        RECT 1404.860 3197.600 1405.140 3198.990 ;
        RECT 2654.360 1614.650 2654.500 3199.070 ;
        RECT 2654.300 1614.330 2654.560 1614.650 ;
        RECT 2900.400 1614.330 2900.660 1614.650 ;
        RECT 2900.460 1613.485 2900.600 1614.330 ;
        RECT 2900.390 1613.115 2900.670 1613.485 ;
      LAYER via2 ;
        RECT 2900.390 1613.160 2900.670 1613.440 ;
      LAYER met3 ;
        RECT 2900.365 1613.450 2900.695 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.365 1613.150 2924.800 1613.450 ;
        RECT 2900.365 1613.135 2900.695 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1444.470 3213.580 1444.790 3213.640 ;
        RECT 1538.310 3213.580 1538.630 3213.640 ;
        RECT 1444.470 3213.440 1538.630 3213.580 ;
        RECT 1444.470 3213.380 1444.790 3213.440 ;
        RECT 1538.310 3213.380 1538.630 3213.440 ;
        RECT 1538.310 3201.000 1538.630 3201.060 ;
        RECT 2899.910 3201.000 2900.230 3201.060 ;
        RECT 1538.310 3200.860 2900.230 3201.000 ;
        RECT 1538.310 3200.800 1538.630 3200.860 ;
        RECT 2899.910 3200.800 2900.230 3200.860 ;
      LAYER via ;
        RECT 1444.500 3213.380 1444.760 3213.640 ;
        RECT 1538.340 3213.380 1538.600 3213.640 ;
        RECT 1538.340 3200.800 1538.600 3201.060 ;
        RECT 2899.940 3200.800 2900.200 3201.060 ;
      LAYER met2 ;
        RECT 1444.500 3213.350 1444.760 3213.670 ;
        RECT 1538.340 3213.350 1538.600 3213.670 ;
        RECT 1444.560 3200.000 1444.700 3213.350 ;
        RECT 1538.400 3201.090 1538.540 3213.350 ;
        RECT 1538.340 3200.770 1538.600 3201.090 ;
        RECT 2899.940 3200.770 2900.200 3201.090 ;
        RECT 1444.420 3197.600 1444.700 3200.000 ;
        RECT 2900.000 1848.085 2900.140 3200.770 ;
        RECT 2899.930 1847.715 2900.210 1848.085 ;
      LAYER via2 ;
        RECT 2899.930 1847.760 2900.210 1848.040 ;
      LAYER met3 ;
        RECT 2899.905 1848.050 2900.235 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2899.905 1847.750 2924.800 1848.050 ;
        RECT 2899.905 1847.735 2900.235 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1484.030 3200.660 1484.350 3200.720 ;
        RECT 2655.650 3200.660 2655.970 3200.720 ;
        RECT 1484.030 3200.520 2655.970 3200.660 ;
        RECT 1484.030 3200.460 1484.350 3200.520 ;
        RECT 2655.650 3200.460 2655.970 3200.520 ;
        RECT 2655.650 2083.760 2655.970 2083.820 ;
        RECT 2899.450 2083.760 2899.770 2083.820 ;
        RECT 2655.650 2083.620 2899.770 2083.760 ;
        RECT 2655.650 2083.560 2655.970 2083.620 ;
        RECT 2899.450 2083.560 2899.770 2083.620 ;
      LAYER via ;
        RECT 1484.060 3200.460 1484.320 3200.720 ;
        RECT 2655.680 3200.460 2655.940 3200.720 ;
        RECT 2655.680 2083.560 2655.940 2083.820 ;
        RECT 2899.480 2083.560 2899.740 2083.820 ;
      LAYER met2 ;
        RECT 1484.060 3200.430 1484.320 3200.750 ;
        RECT 2655.680 3200.430 2655.940 3200.750 ;
        RECT 1484.120 3200.000 1484.260 3200.430 ;
        RECT 1483.980 3197.600 1484.260 3200.000 ;
        RECT 2655.740 2083.850 2655.880 3200.430 ;
        RECT 2655.680 2083.530 2655.940 2083.850 ;
        RECT 2899.480 2083.530 2899.740 2083.850 ;
        RECT 2899.540 2082.685 2899.680 2083.530 ;
        RECT 2899.470 2082.315 2899.750 2082.685 ;
      LAYER via2 ;
        RECT 2899.470 2082.360 2899.750 2082.640 ;
      LAYER met3 ;
        RECT 2899.445 2082.650 2899.775 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2899.445 2082.350 2924.800 2082.650 ;
        RECT 2899.445 2082.335 2899.775 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1523.130 3213.240 1523.450 3213.300 ;
        RECT 2660.250 3213.240 2660.570 3213.300 ;
        RECT 1523.130 3213.100 2660.570 3213.240 ;
        RECT 1523.130 3213.040 1523.450 3213.100 ;
        RECT 2660.250 3213.040 2660.570 3213.100 ;
        RECT 2660.250 2318.360 2660.570 2318.420 ;
        RECT 2898.990 2318.360 2899.310 2318.420 ;
        RECT 2660.250 2318.220 2899.310 2318.360 ;
        RECT 2660.250 2318.160 2660.570 2318.220 ;
        RECT 2898.990 2318.160 2899.310 2318.220 ;
      LAYER via ;
        RECT 1523.160 3213.040 1523.420 3213.300 ;
        RECT 2660.280 3213.040 2660.540 3213.300 ;
        RECT 2660.280 2318.160 2660.540 2318.420 ;
        RECT 2899.020 2318.160 2899.280 2318.420 ;
      LAYER met2 ;
        RECT 1523.160 3213.010 1523.420 3213.330 ;
        RECT 2660.280 3213.010 2660.540 3213.330 ;
        RECT 1523.220 3200.000 1523.360 3213.010 ;
        RECT 1523.080 3197.600 1523.360 3200.000 ;
        RECT 2660.340 2318.450 2660.480 3213.010 ;
        RECT 2660.280 2318.130 2660.540 2318.450 ;
        RECT 2899.020 2318.130 2899.280 2318.450 ;
        RECT 2899.080 2317.285 2899.220 2318.130 ;
        RECT 2899.010 2316.915 2899.290 2317.285 ;
      LAYER via2 ;
        RECT 2899.010 2316.960 2899.290 2317.240 ;
      LAYER met3 ;
        RECT 2898.985 2317.250 2899.315 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2898.985 2316.950 2924.800 2317.250 ;
        RECT 2898.985 2316.935 2899.315 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1181.350 3212.900 1181.670 3212.960 ;
        RECT 1449.990 3212.900 1450.310 3212.960 ;
        RECT 1181.350 3212.760 1450.310 3212.900 ;
        RECT 1181.350 3212.700 1181.670 3212.760 ;
        RECT 1449.990 3212.700 1450.310 3212.760 ;
      LAYER via ;
        RECT 1181.380 3212.700 1181.640 3212.960 ;
        RECT 1450.020 3212.700 1450.280 3212.960 ;
      LAYER met2 ;
        RECT 1181.380 3212.670 1181.640 3212.990 ;
        RECT 1450.020 3212.670 1450.280 3212.990 ;
        RECT 1181.440 3200.000 1181.580 3212.670 ;
        RECT 1181.300 3197.600 1181.580 3200.000 ;
        RECT 1450.080 3199.245 1450.220 3212.670 ;
        RECT 1450.010 3198.875 1450.290 3199.245 ;
        RECT 1703.930 3199.130 1704.210 3199.245 ;
        RECT 1704.850 3199.130 1705.130 3199.245 ;
        RECT 1703.930 3198.990 1705.130 3199.130 ;
        RECT 1703.930 3198.875 1704.210 3198.990 ;
        RECT 1704.850 3198.875 1705.130 3198.990 ;
        RECT 2898.090 3198.875 2898.370 3199.245 ;
        RECT 2898.160 3195.845 2898.300 3198.875 ;
        RECT 2898.090 3195.475 2898.370 3195.845 ;
        RECT 2901.310 3195.475 2901.590 3195.845 ;
        RECT 2901.380 146.725 2901.520 3195.475 ;
        RECT 2901.310 146.355 2901.590 146.725 ;
      LAYER via2 ;
        RECT 1450.010 3198.920 1450.290 3199.200 ;
        RECT 1703.930 3198.920 1704.210 3199.200 ;
        RECT 1704.850 3198.920 1705.130 3199.200 ;
        RECT 2898.090 3198.920 2898.370 3199.200 ;
        RECT 2898.090 3195.520 2898.370 3195.800 ;
        RECT 2901.310 3195.520 2901.590 3195.800 ;
        RECT 2901.310 146.400 2901.590 146.680 ;
      LAYER met3 ;
        RECT 1449.985 3199.210 1450.315 3199.225 ;
        RECT 1703.905 3199.210 1704.235 3199.225 ;
        RECT 1449.985 3198.910 1704.235 3199.210 ;
        RECT 1449.985 3198.895 1450.315 3198.910 ;
        RECT 1703.905 3198.895 1704.235 3198.910 ;
        RECT 1704.825 3199.210 1705.155 3199.225 ;
        RECT 2898.065 3199.210 2898.395 3199.225 ;
        RECT 1704.825 3198.910 2898.395 3199.210 ;
        RECT 1704.825 3198.895 1705.155 3198.910 ;
        RECT 2898.065 3198.895 2898.395 3198.910 ;
        RECT 2898.065 3195.810 2898.395 3195.825 ;
        RECT 2901.285 3195.810 2901.615 3195.825 ;
        RECT 2898.065 3195.510 2901.615 3195.810 ;
        RECT 2898.065 3195.495 2898.395 3195.510 ;
        RECT 2901.285 3195.495 2901.615 3195.510 ;
        RECT 2901.285 146.690 2901.615 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2901.285 146.390 2924.800 146.690 ;
        RECT 2901.285 146.375 2901.615 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1576.030 3213.580 1576.350 3213.640 ;
        RECT 2660.710 3213.580 2661.030 3213.640 ;
        RECT 1576.030 3213.440 2661.030 3213.580 ;
        RECT 1576.030 3213.380 1576.350 3213.440 ;
        RECT 2660.710 3213.380 2661.030 3213.440 ;
        RECT 2660.710 2497.540 2661.030 2497.600 ;
        RECT 2898.990 2497.540 2899.310 2497.600 ;
        RECT 2660.710 2497.400 2899.310 2497.540 ;
        RECT 2660.710 2497.340 2661.030 2497.400 ;
        RECT 2898.990 2497.340 2899.310 2497.400 ;
      LAYER via ;
        RECT 1576.060 3213.380 1576.320 3213.640 ;
        RECT 2660.740 3213.380 2661.000 3213.640 ;
        RECT 2660.740 2497.340 2661.000 2497.600 ;
        RECT 2899.020 2497.340 2899.280 2497.600 ;
      LAYER met2 ;
        RECT 1576.060 3213.350 1576.320 3213.670 ;
        RECT 2660.740 3213.350 2661.000 3213.670 ;
        RECT 1576.120 3200.000 1576.260 3213.350 ;
        RECT 1575.980 3197.600 1576.260 3200.000 ;
        RECT 2660.800 2497.630 2660.940 3213.350 ;
        RECT 2660.740 2497.310 2661.000 2497.630 ;
        RECT 2899.020 2497.310 2899.280 2497.630 ;
        RECT 2899.080 2493.405 2899.220 2497.310 ;
        RECT 2899.010 2493.035 2899.290 2493.405 ;
      LAYER via2 ;
        RECT 2899.010 2493.080 2899.290 2493.360 ;
      LAYER met3 ;
        RECT 2898.985 2493.370 2899.315 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2898.985 2493.070 2924.800 2493.370 ;
        RECT 2898.985 2493.055 2899.315 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1615.590 3214.260 1615.910 3214.320 ;
        RECT 2661.170 3214.260 2661.490 3214.320 ;
        RECT 1615.590 3214.120 2661.490 3214.260 ;
        RECT 1615.590 3214.060 1615.910 3214.120 ;
        RECT 2661.170 3214.060 2661.490 3214.120 ;
        RECT 2661.170 2732.140 2661.490 2732.200 ;
        RECT 2898.990 2732.140 2899.310 2732.200 ;
        RECT 2661.170 2732.000 2899.310 2732.140 ;
        RECT 2661.170 2731.940 2661.490 2732.000 ;
        RECT 2898.990 2731.940 2899.310 2732.000 ;
      LAYER via ;
        RECT 1615.620 3214.060 1615.880 3214.320 ;
        RECT 2661.200 3214.060 2661.460 3214.320 ;
        RECT 2661.200 2731.940 2661.460 2732.200 ;
        RECT 2899.020 2731.940 2899.280 2732.200 ;
      LAYER met2 ;
        RECT 1615.620 3214.030 1615.880 3214.350 ;
        RECT 2661.200 3214.030 2661.460 3214.350 ;
        RECT 1615.680 3200.000 1615.820 3214.030 ;
        RECT 1615.540 3197.600 1615.820 3200.000 ;
        RECT 2661.260 2732.230 2661.400 3214.030 ;
        RECT 2661.200 2731.910 2661.460 2732.230 ;
        RECT 2899.020 2731.910 2899.280 2732.230 ;
        RECT 2899.080 2728.005 2899.220 2731.910 ;
        RECT 2899.010 2727.635 2899.290 2728.005 ;
      LAYER via2 ;
        RECT 2899.010 2727.680 2899.290 2727.960 ;
      LAYER met3 ;
        RECT 2898.985 2727.970 2899.315 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2898.985 2727.670 2924.800 2727.970 ;
        RECT 2898.985 2727.655 2899.315 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1655.150 3214.600 1655.470 3214.660 ;
        RECT 2661.630 3214.600 2661.950 3214.660 ;
        RECT 1655.150 3214.460 2661.950 3214.600 ;
        RECT 1655.150 3214.400 1655.470 3214.460 ;
        RECT 2661.630 3214.400 2661.950 3214.460 ;
        RECT 2661.630 2966.740 2661.950 2966.800 ;
        RECT 2898.990 2966.740 2899.310 2966.800 ;
        RECT 2661.630 2966.600 2899.310 2966.740 ;
        RECT 2661.630 2966.540 2661.950 2966.600 ;
        RECT 2898.990 2966.540 2899.310 2966.600 ;
      LAYER via ;
        RECT 1655.180 3214.400 1655.440 3214.660 ;
        RECT 2661.660 3214.400 2661.920 3214.660 ;
        RECT 2661.660 2966.540 2661.920 2966.800 ;
        RECT 2899.020 2966.540 2899.280 2966.800 ;
      LAYER met2 ;
        RECT 1655.180 3214.370 1655.440 3214.690 ;
        RECT 2661.660 3214.370 2661.920 3214.690 ;
        RECT 1655.240 3200.000 1655.380 3214.370 ;
        RECT 1655.100 3197.600 1655.380 3200.000 ;
        RECT 2661.720 2966.830 2661.860 3214.370 ;
        RECT 2661.660 2966.510 2661.920 2966.830 ;
        RECT 2899.020 2966.510 2899.280 2966.830 ;
        RECT 2899.080 2962.605 2899.220 2966.510 ;
        RECT 2899.010 2962.235 2899.290 2962.605 ;
      LAYER via2 ;
        RECT 2899.010 2962.280 2899.290 2962.560 ;
      LAYER met3 ;
        RECT 2898.985 2962.570 2899.315 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2898.985 2962.270 2924.800 2962.570 ;
        RECT 2898.985 2962.255 2899.315 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1696.090 3200.320 1696.410 3200.380 ;
        RECT 2900.830 3200.320 2901.150 3200.380 ;
        RECT 1696.090 3200.180 2901.150 3200.320 ;
        RECT 1696.090 3200.120 1696.410 3200.180 ;
        RECT 2900.830 3200.120 2901.150 3200.180 ;
      LAYER via ;
        RECT 1696.120 3200.120 1696.380 3200.380 ;
        RECT 2900.860 3200.120 2901.120 3200.380 ;
      LAYER met2 ;
        RECT 1696.120 3200.090 1696.380 3200.410 ;
        RECT 2900.860 3200.090 2901.120 3200.410 ;
        RECT 1694.200 3199.810 1694.480 3200.000 ;
        RECT 1696.180 3199.810 1696.320 3200.090 ;
        RECT 1694.200 3199.670 1696.320 3199.810 ;
        RECT 1694.200 3197.600 1694.480 3199.670 ;
        RECT 2900.920 3197.205 2901.060 3200.090 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2146.060 3429.680 2149.880 3429.820 ;
        RECT 1738.410 3429.480 1738.730 3429.540 ;
        RECT 2146.060 3429.480 2146.200 3429.680 ;
        RECT 1738.410 3429.340 2146.200 3429.480 ;
        RECT 2149.740 3429.480 2149.880 3429.680 ;
        RECT 2762.920 3429.680 2798.940 3429.820 ;
        RECT 2762.920 3429.480 2763.060 3429.680 ;
        RECT 2149.740 3429.340 2763.060 3429.480 ;
        RECT 2798.800 3429.480 2798.940 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2798.800 3429.340 2901.150 3429.480 ;
        RECT 1738.410 3429.280 1738.730 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 1738.440 3429.280 1738.700 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1738.440 3429.250 1738.700 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1738.500 3200.490 1738.640 3429.250 ;
        RECT 1736.660 3200.350 1738.640 3200.490 ;
        RECT 1733.760 3199.130 1734.040 3200.000 ;
        RECT 1736.660 3199.130 1736.800 3200.350 ;
        RECT 1733.760 3198.990 1736.800 3199.130 ;
        RECT 1733.760 3197.600 1734.040 3198.990 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1779.810 3504.620 1780.130 3504.680 ;
        RECT 2717.290 3504.620 2717.610 3504.680 ;
        RECT 1779.810 3504.480 2717.610 3504.620 ;
        RECT 1779.810 3504.420 1780.130 3504.480 ;
        RECT 2717.290 3504.420 2717.610 3504.480 ;
      LAYER via ;
        RECT 1779.840 3504.420 1780.100 3504.680 ;
        RECT 2717.320 3504.420 2717.580 3504.680 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3504.710 2717.520 3517.600 ;
        RECT 1779.840 3504.390 1780.100 3504.710 ;
        RECT 2717.320 3504.390 2717.580 3504.710 ;
        RECT 1779.900 3200.490 1780.040 3504.390 ;
        RECT 1776.680 3200.350 1780.040 3200.490 ;
        RECT 1773.320 3199.810 1773.600 3200.000 ;
        RECT 1776.680 3199.810 1776.820 3200.350 ;
        RECT 1773.320 3199.670 1776.820 3199.810 ;
        RECT 1773.320 3197.600 1773.600 3199.670 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1814.310 3500.540 1814.630 3500.600 ;
        RECT 2392.530 3500.540 2392.850 3500.600 ;
        RECT 1814.310 3500.400 2392.850 3500.540 ;
        RECT 1814.310 3500.340 1814.630 3500.400 ;
        RECT 2392.530 3500.340 2392.850 3500.400 ;
      LAYER via ;
        RECT 1814.340 3500.340 1814.600 3500.600 ;
        RECT 2392.560 3500.340 2392.820 3500.600 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3500.630 2392.760 3517.600 ;
        RECT 1814.340 3500.310 1814.600 3500.630 ;
        RECT 2392.560 3500.310 2392.820 3500.630 ;
        RECT 1812.880 3199.810 1813.160 3200.000 ;
        RECT 1814.400 3199.810 1814.540 3500.310 ;
        RECT 1812.880 3199.670 1814.540 3199.810 ;
        RECT 1812.880 3197.600 1813.160 3199.670 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.710 3499.180 1856.030 3499.240 ;
        RECT 2068.230 3499.180 2068.550 3499.240 ;
        RECT 1855.710 3499.040 2068.550 3499.180 ;
        RECT 1855.710 3498.980 1856.030 3499.040 ;
        RECT 2068.230 3498.980 2068.550 3499.040 ;
      LAYER via ;
        RECT 1855.740 3498.980 1856.000 3499.240 ;
        RECT 2068.260 3498.980 2068.520 3499.240 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3499.270 2068.460 3517.600 ;
        RECT 1855.740 3498.950 1856.000 3499.270 ;
        RECT 2068.260 3498.950 2068.520 3499.270 ;
        RECT 1852.440 3199.130 1852.720 3200.000 ;
        RECT 1855.800 3199.130 1855.940 3498.950 ;
        RECT 1852.440 3198.990 1855.940 3199.130 ;
        RECT 1852.440 3197.600 1852.720 3198.990 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1743.930 3498.840 1744.250 3498.900 ;
        RECT 1890.670 3498.840 1890.990 3498.900 ;
        RECT 1743.930 3498.700 1890.990 3498.840 ;
        RECT 1743.930 3498.640 1744.250 3498.700 ;
        RECT 1890.670 3498.640 1890.990 3498.700 ;
      LAYER via ;
        RECT 1743.960 3498.640 1744.220 3498.900 ;
        RECT 1890.700 3498.640 1890.960 3498.900 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3498.930 1744.160 3517.600 ;
        RECT 1743.960 3498.610 1744.220 3498.930 ;
        RECT 1890.700 3498.610 1890.960 3498.930 ;
        RECT 1890.760 3199.810 1890.900 3498.610 ;
        RECT 1891.540 3199.810 1891.820 3200.000 ;
        RECT 1890.760 3199.670 1891.820 3199.810 ;
        RECT 1891.540 3197.600 1891.820 3199.670 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3499.860 1419.490 3499.920 ;
        RECT 1925.170 3499.860 1925.490 3499.920 ;
        RECT 1419.170 3499.720 1925.490 3499.860 ;
        RECT 1419.170 3499.660 1419.490 3499.720 ;
        RECT 1925.170 3499.660 1925.490 3499.720 ;
      LAYER via ;
        RECT 1419.200 3499.660 1419.460 3499.920 ;
        RECT 1925.200 3499.660 1925.460 3499.920 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3499.950 1419.400 3517.600 ;
        RECT 1419.200 3499.630 1419.460 3499.950 ;
        RECT 1925.200 3499.630 1925.460 3499.950 ;
        RECT 1925.260 3200.490 1925.400 3499.630 ;
        RECT 1925.260 3200.350 1928.620 3200.490 ;
        RECT 1928.480 3199.130 1928.620 3200.350 ;
        RECT 1931.100 3199.130 1931.380 3200.000 ;
        RECT 1928.480 3198.990 1931.380 3199.130 ;
        RECT 1931.100 3197.600 1931.380 3198.990 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1220.930 3200.235 1221.210 3200.605 ;
        RECT 1221.000 3200.000 1221.140 3200.235 ;
        RECT 1220.860 3197.600 1221.140 3200.000 ;
        RECT 2902.230 3196.155 2902.510 3196.525 ;
        RECT 2902.300 381.325 2902.440 3196.155 ;
        RECT 2902.230 380.955 2902.510 381.325 ;
      LAYER via2 ;
        RECT 1220.930 3200.280 1221.210 3200.560 ;
        RECT 2902.230 3196.200 2902.510 3196.480 ;
        RECT 2902.230 381.000 2902.510 381.280 ;
      LAYER met3 ;
        RECT 1220.905 3200.570 1221.235 3200.585 ;
        RECT 1260.670 3200.570 1261.050 3200.580 ;
        RECT 1220.905 3200.270 1261.050 3200.570 ;
        RECT 1220.905 3200.255 1221.235 3200.270 ;
        RECT 1260.670 3200.260 1261.050 3200.270 ;
        RECT 1260.670 3196.490 1261.050 3196.500 ;
        RECT 2902.205 3196.490 2902.535 3196.505 ;
        RECT 1260.670 3196.190 2902.535 3196.490 ;
        RECT 1260.670 3196.180 1261.050 3196.190 ;
        RECT 2902.205 3196.175 2902.535 3196.190 ;
        RECT 2902.205 381.290 2902.535 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2902.205 380.990 2924.800 381.290 ;
        RECT 2902.205 380.975 2902.535 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
      LAYER via3 ;
        RECT 1260.700 3200.260 1261.020 3200.580 ;
        RECT 1260.700 3196.180 1261.020 3196.500 ;
      LAYER met4 ;
        RECT 1260.695 3200.255 1261.025 3200.585 ;
        RECT 1260.710 3196.505 1261.010 3200.255 ;
        RECT 1260.695 3196.175 1261.025 3196.505 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3504.960 1095.190 3505.020 ;
        RECT 1966.570 3504.960 1966.890 3505.020 ;
        RECT 1094.870 3504.820 1966.890 3504.960 ;
        RECT 1094.870 3504.760 1095.190 3504.820 ;
        RECT 1966.570 3504.760 1966.890 3504.820 ;
      LAYER via ;
        RECT 1094.900 3504.760 1095.160 3505.020 ;
        RECT 1966.600 3504.760 1966.860 3505.020 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3505.050 1095.100 3517.600 ;
        RECT 1094.900 3504.730 1095.160 3505.050 ;
        RECT 1966.600 3504.730 1966.860 3505.050 ;
        RECT 1966.660 3199.130 1966.800 3504.730 ;
        RECT 1970.660 3199.130 1970.940 3200.000 ;
        RECT 1966.660 3198.990 1970.940 3199.130 ;
        RECT 1970.660 3197.600 1970.940 3198.990 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3503.600 770.890 3503.660 ;
        RECT 2007.970 3503.600 2008.290 3503.660 ;
        RECT 770.570 3503.460 2008.290 3503.600 ;
        RECT 770.570 3503.400 770.890 3503.460 ;
        RECT 2007.970 3503.400 2008.290 3503.460 ;
      LAYER via ;
        RECT 770.600 3503.400 770.860 3503.660 ;
        RECT 2008.000 3503.400 2008.260 3503.660 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3503.690 770.800 3517.600 ;
        RECT 770.600 3503.370 770.860 3503.690 ;
        RECT 2008.000 3503.370 2008.260 3503.690 ;
        RECT 2008.060 3199.810 2008.200 3503.370 ;
        RECT 2010.220 3199.810 2010.500 3200.000 ;
        RECT 2008.060 3199.670 2010.500 3199.810 ;
        RECT 2010.220 3197.600 2010.500 3199.670 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3502.580 446.130 3502.640 ;
        RECT 2049.370 3502.580 2049.690 3502.640 ;
        RECT 445.810 3502.440 2049.690 3502.580 ;
        RECT 445.810 3502.380 446.130 3502.440 ;
        RECT 2049.370 3502.380 2049.690 3502.440 ;
      LAYER via ;
        RECT 445.840 3502.380 446.100 3502.640 ;
        RECT 2049.400 3502.380 2049.660 3502.640 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3502.670 446.040 3517.600 ;
        RECT 445.840 3502.350 446.100 3502.670 ;
        RECT 2049.400 3502.350 2049.660 3502.670 ;
        RECT 2049.460 3199.810 2049.600 3502.350 ;
        RECT 2049.780 3199.810 2050.060 3200.000 ;
        RECT 2049.460 3199.670 2050.060 3199.810 ;
        RECT 2049.780 3197.600 2050.060 3199.670 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 2083.870 3501.560 2084.190 3501.620 ;
        RECT 121.510 3501.420 2084.190 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 2083.870 3501.360 2084.190 3501.420 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 2083.900 3501.360 2084.160 3501.620 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 2083.900 3501.330 2084.160 3501.650 ;
        RECT 2083.960 3199.130 2084.100 3501.330 ;
        RECT 2088.880 3199.130 2089.160 3200.000 ;
        RECT 2083.960 3198.990 2089.160 3199.130 ;
        RECT 2088.880 3197.600 2089.160 3198.990 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 2125.270 3339.720 2125.590 3339.780 ;
        RECT 17.090 3339.580 2125.590 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 2125.270 3339.520 2125.590 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 2125.300 3339.520 2125.560 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 2125.300 3339.490 2125.560 3339.810 ;
        RECT 2125.360 3201.170 2125.500 3339.490 ;
        RECT 2125.360 3201.030 2126.880 3201.170 ;
        RECT 2126.740 3199.810 2126.880 3201.030 ;
        RECT 2128.440 3199.810 2128.720 3200.000 ;
        RECT 2126.740 3199.670 2128.720 3199.810 ;
        RECT 2128.440 3197.600 2128.720 3199.670 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 27.210 3211.200 27.530 3211.260 ;
        RECT 2168.050 3211.200 2168.370 3211.260 ;
        RECT 27.210 3211.060 2168.370 3211.200 ;
        RECT 27.210 3211.000 27.530 3211.060 ;
        RECT 2168.050 3211.000 2168.370 3211.060 ;
        RECT 13.870 3053.100 14.190 3053.160 ;
        RECT 27.210 3053.100 27.530 3053.160 ;
        RECT 13.870 3052.960 27.530 3053.100 ;
        RECT 13.870 3052.900 14.190 3052.960 ;
        RECT 27.210 3052.900 27.530 3052.960 ;
      LAYER via ;
        RECT 27.240 3211.000 27.500 3211.260 ;
        RECT 2168.080 3211.000 2168.340 3211.260 ;
        RECT 13.900 3052.900 14.160 3053.160 ;
        RECT 27.240 3052.900 27.500 3053.160 ;
      LAYER met2 ;
        RECT 27.240 3210.970 27.500 3211.290 ;
        RECT 2168.080 3210.970 2168.340 3211.290 ;
        RECT 27.300 3053.190 27.440 3210.970 ;
        RECT 2168.140 3200.000 2168.280 3210.970 ;
        RECT 2168.000 3197.600 2168.280 3200.000 ;
        RECT 13.900 3052.870 14.160 3053.190 ;
        RECT 27.240 3052.870 27.500 3053.190 ;
        RECT 13.960 3052.365 14.100 3052.870 ;
        RECT 13.890 3051.995 14.170 3052.365 ;
      LAYER via2 ;
        RECT 13.890 3052.040 14.170 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 13.865 3052.330 14.195 3052.345 ;
        RECT -4.800 3052.030 14.195 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 13.865 3052.015 14.195 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.750 3210.860 27.070 3210.920 ;
        RECT 2207.610 3210.860 2207.930 3210.920 ;
        RECT 26.750 3210.720 2207.930 3210.860 ;
        RECT 26.750 3210.660 27.070 3210.720 ;
        RECT 2207.610 3210.660 2207.930 3210.720 ;
        RECT 13.870 2765.460 14.190 2765.520 ;
        RECT 26.750 2765.460 27.070 2765.520 ;
        RECT 13.870 2765.320 27.070 2765.460 ;
        RECT 13.870 2765.260 14.190 2765.320 ;
        RECT 26.750 2765.260 27.070 2765.320 ;
      LAYER via ;
        RECT 26.780 3210.660 27.040 3210.920 ;
        RECT 2207.640 3210.660 2207.900 3210.920 ;
        RECT 13.900 2765.260 14.160 2765.520 ;
        RECT 26.780 2765.260 27.040 2765.520 ;
      LAYER met2 ;
        RECT 26.780 3210.630 27.040 3210.950 ;
        RECT 2207.640 3210.630 2207.900 3210.950 ;
        RECT 26.840 2765.550 26.980 3210.630 ;
        RECT 2207.700 3200.000 2207.840 3210.630 ;
        RECT 2207.560 3197.600 2207.840 3200.000 ;
        RECT 13.900 2765.405 14.160 2765.550 ;
        RECT 13.890 2765.035 14.170 2765.405 ;
        RECT 26.780 2765.230 27.040 2765.550 ;
      LAYER via2 ;
        RECT 13.890 2765.080 14.170 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 13.865 2765.370 14.195 2765.385 ;
        RECT -4.800 2765.070 14.195 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 13.865 2765.055 14.195 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.290 3210.180 26.610 3210.240 ;
        RECT 2247.170 3210.180 2247.490 3210.240 ;
        RECT 26.290 3210.040 2247.490 3210.180 ;
        RECT 26.290 3209.980 26.610 3210.040 ;
        RECT 2247.170 3209.980 2247.490 3210.040 ;
        RECT 13.870 2483.600 14.190 2483.660 ;
        RECT 26.290 2483.600 26.610 2483.660 ;
        RECT 13.870 2483.460 26.610 2483.600 ;
        RECT 13.870 2483.400 14.190 2483.460 ;
        RECT 26.290 2483.400 26.610 2483.460 ;
      LAYER via ;
        RECT 26.320 3209.980 26.580 3210.240 ;
        RECT 2247.200 3209.980 2247.460 3210.240 ;
        RECT 13.900 2483.400 14.160 2483.660 ;
        RECT 26.320 2483.400 26.580 2483.660 ;
      LAYER met2 ;
        RECT 26.320 3209.950 26.580 3210.270 ;
        RECT 2247.200 3209.950 2247.460 3210.270 ;
        RECT 26.380 2483.690 26.520 3209.950 ;
        RECT 2247.260 3200.000 2247.400 3209.950 ;
        RECT 2247.120 3197.600 2247.400 3200.000 ;
        RECT 13.900 2483.370 14.160 2483.690 ;
        RECT 26.320 2483.370 26.580 2483.690 ;
        RECT 13.960 2477.765 14.100 2483.370 ;
        RECT 13.890 2477.395 14.170 2477.765 ;
      LAYER via2 ;
        RECT 13.890 2477.440 14.170 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 13.865 2477.730 14.195 2477.745 ;
        RECT -4.800 2477.430 14.195 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 13.865 2477.415 14.195 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 186.905 3197.785 187.535 3197.955 ;
        RECT 966.145 3197.785 967.235 3197.955 ;
        RECT 1063.205 3197.785 1063.835 3197.955 ;
        RECT 1148.765 3197.785 1148.935 3198.975 ;
        RECT 1197.065 3197.785 1197.235 3198.975 ;
        RECT 1238.005 3197.785 1238.175 3198.975 ;
        RECT 1289.985 3197.785 1290.155 3198.975 ;
        RECT 1338.745 3197.785 1338.915 3199.315 ;
        RECT 1386.585 3197.785 1386.755 3199.315 ;
        RECT 1435.345 3197.785 1435.515 3200.335 ;
        RECT 1462.945 3197.785 1463.115 3200.335 ;
        RECT 1535.165 3197.785 1535.335 3200.335 ;
        RECT 1559.545 3197.785 1559.715 3200.335 ;
        RECT 1629.005 3197.785 1629.175 3200.335 ;
        RECT 1680.065 3197.785 1680.235 3200.335 ;
        RECT 1725.145 3197.785 1725.315 3208.495 ;
        RECT 1772.985 3197.785 1773.155 3208.495 ;
        RECT 1821.745 3197.785 1821.915 3208.495 ;
        RECT 1869.585 3197.785 1869.755 3208.495 ;
        RECT 1918.345 3197.785 1918.515 3208.495 ;
        RECT 1966.185 3197.785 1966.355 3208.495 ;
        RECT 2014.945 3197.785 2015.115 3208.495 ;
        RECT 2062.785 3197.785 2062.955 3208.495 ;
        RECT 2208.145 3197.785 2208.315 3198.635 ;
      LAYER mcon ;
        RECT 1725.145 3208.325 1725.315 3208.495 ;
        RECT 1435.345 3200.165 1435.515 3200.335 ;
        RECT 1338.745 3199.145 1338.915 3199.315 ;
        RECT 1148.765 3198.805 1148.935 3198.975 ;
        RECT 187.365 3197.785 187.535 3197.955 ;
        RECT 967.065 3197.785 967.235 3197.955 ;
        RECT 1063.665 3197.785 1063.835 3197.955 ;
        RECT 1197.065 3198.805 1197.235 3198.975 ;
        RECT 1238.005 3198.805 1238.175 3198.975 ;
        RECT 1289.985 3198.805 1290.155 3198.975 ;
        RECT 1386.585 3199.145 1386.755 3199.315 ;
        RECT 1462.945 3200.165 1463.115 3200.335 ;
        RECT 1535.165 3200.165 1535.335 3200.335 ;
        RECT 1559.545 3200.165 1559.715 3200.335 ;
        RECT 1629.005 3200.165 1629.175 3200.335 ;
        RECT 1680.065 3200.165 1680.235 3200.335 ;
        RECT 1772.985 3208.325 1773.155 3208.495 ;
        RECT 1821.745 3208.325 1821.915 3208.495 ;
        RECT 1869.585 3208.325 1869.755 3208.495 ;
        RECT 1918.345 3208.325 1918.515 3208.495 ;
        RECT 1966.185 3208.325 1966.355 3208.495 ;
        RECT 2014.945 3208.325 2015.115 3208.495 ;
        RECT 2062.785 3208.325 2062.955 3208.495 ;
        RECT 2208.145 3198.465 2208.315 3198.635 ;
      LAYER met1 ;
        RECT 1725.085 3208.480 1725.375 3208.525 ;
        RECT 1772.925 3208.480 1773.215 3208.525 ;
        RECT 1725.085 3208.340 1773.215 3208.480 ;
        RECT 1725.085 3208.295 1725.375 3208.340 ;
        RECT 1772.925 3208.295 1773.215 3208.340 ;
        RECT 1821.685 3208.480 1821.975 3208.525 ;
        RECT 1869.525 3208.480 1869.815 3208.525 ;
        RECT 1821.685 3208.340 1869.815 3208.480 ;
        RECT 1821.685 3208.295 1821.975 3208.340 ;
        RECT 1869.525 3208.295 1869.815 3208.340 ;
        RECT 1918.285 3208.480 1918.575 3208.525 ;
        RECT 1966.125 3208.480 1966.415 3208.525 ;
        RECT 1918.285 3208.340 1966.415 3208.480 ;
        RECT 1918.285 3208.295 1918.575 3208.340 ;
        RECT 1966.125 3208.295 1966.415 3208.340 ;
        RECT 2014.885 3208.480 2015.175 3208.525 ;
        RECT 2062.725 3208.480 2063.015 3208.525 ;
        RECT 2014.885 3208.340 2063.015 3208.480 ;
        RECT 2014.885 3208.295 2015.175 3208.340 ;
        RECT 2062.725 3208.295 2063.015 3208.340 ;
        RECT 1435.285 3200.320 1435.575 3200.365 ;
        RECT 1462.885 3200.320 1463.175 3200.365 ;
        RECT 1435.285 3200.180 1463.175 3200.320 ;
        RECT 1435.285 3200.135 1435.575 3200.180 ;
        RECT 1462.885 3200.135 1463.175 3200.180 ;
        RECT 1535.105 3200.320 1535.395 3200.365 ;
        RECT 1559.485 3200.320 1559.775 3200.365 ;
        RECT 1535.105 3200.180 1559.775 3200.320 ;
        RECT 1535.105 3200.135 1535.395 3200.180 ;
        RECT 1559.485 3200.135 1559.775 3200.180 ;
        RECT 1628.945 3200.320 1629.235 3200.365 ;
        RECT 1680.005 3200.320 1680.295 3200.365 ;
        RECT 1628.945 3200.180 1680.295 3200.320 ;
        RECT 1628.945 3200.135 1629.235 3200.180 ;
        RECT 1680.005 3200.135 1680.295 3200.180 ;
        RECT 1338.685 3199.300 1338.975 3199.345 ;
        RECT 1386.525 3199.300 1386.815 3199.345 ;
        RECT 1338.685 3199.160 1386.815 3199.300 ;
        RECT 1338.685 3199.115 1338.975 3199.160 ;
        RECT 1386.525 3199.115 1386.815 3199.160 ;
        RECT 1148.705 3198.960 1148.995 3199.005 ;
        RECT 1197.005 3198.960 1197.295 3199.005 ;
        RECT 1148.705 3198.820 1197.295 3198.960 ;
        RECT 1148.705 3198.775 1148.995 3198.820 ;
        RECT 1197.005 3198.775 1197.295 3198.820 ;
        RECT 1237.945 3198.960 1238.235 3199.005 ;
        RECT 1289.925 3198.960 1290.215 3199.005 ;
        RECT 1237.945 3198.820 1290.215 3198.960 ;
        RECT 1237.945 3198.775 1238.235 3198.820 ;
        RECT 1289.925 3198.775 1290.215 3198.820 ;
        RECT 2208.085 3198.620 2208.375 3198.665 ;
        RECT 2285.350 3198.620 2285.670 3198.680 ;
        RECT 2208.085 3198.480 2285.670 3198.620 ;
        RECT 2208.085 3198.435 2208.375 3198.480 ;
        RECT 2285.350 3198.420 2285.670 3198.480 ;
        RECT 39.170 3197.940 39.490 3198.000 ;
        RECT 186.845 3197.940 187.135 3197.985 ;
        RECT 39.170 3197.800 187.135 3197.940 ;
        RECT 39.170 3197.740 39.490 3197.800 ;
        RECT 186.845 3197.755 187.135 3197.800 ;
        RECT 187.305 3197.940 187.595 3197.985 ;
        RECT 966.085 3197.940 966.375 3197.985 ;
        RECT 187.305 3197.800 966.375 3197.940 ;
        RECT 187.305 3197.755 187.595 3197.800 ;
        RECT 966.085 3197.755 966.375 3197.800 ;
        RECT 967.005 3197.940 967.295 3197.985 ;
        RECT 1063.145 3197.940 1063.435 3197.985 ;
        RECT 967.005 3197.800 1063.435 3197.940 ;
        RECT 967.005 3197.755 967.295 3197.800 ;
        RECT 1063.145 3197.755 1063.435 3197.800 ;
        RECT 1063.605 3197.940 1063.895 3197.985 ;
        RECT 1148.705 3197.940 1148.995 3197.985 ;
        RECT 1063.605 3197.800 1148.995 3197.940 ;
        RECT 1063.605 3197.755 1063.895 3197.800 ;
        RECT 1148.705 3197.755 1148.995 3197.800 ;
        RECT 1197.005 3197.940 1197.295 3197.985 ;
        RECT 1237.945 3197.940 1238.235 3197.985 ;
        RECT 1197.005 3197.800 1238.235 3197.940 ;
        RECT 1197.005 3197.755 1197.295 3197.800 ;
        RECT 1237.945 3197.755 1238.235 3197.800 ;
        RECT 1289.925 3197.940 1290.215 3197.985 ;
        RECT 1338.685 3197.940 1338.975 3197.985 ;
        RECT 1289.925 3197.800 1338.975 3197.940 ;
        RECT 1289.925 3197.755 1290.215 3197.800 ;
        RECT 1338.685 3197.755 1338.975 3197.800 ;
        RECT 1386.525 3197.940 1386.815 3197.985 ;
        RECT 1435.285 3197.940 1435.575 3197.985 ;
        RECT 1386.525 3197.800 1435.575 3197.940 ;
        RECT 1386.525 3197.755 1386.815 3197.800 ;
        RECT 1435.285 3197.755 1435.575 3197.800 ;
        RECT 1462.885 3197.940 1463.175 3197.985 ;
        RECT 1535.105 3197.940 1535.395 3197.985 ;
        RECT 1462.885 3197.800 1535.395 3197.940 ;
        RECT 1462.885 3197.755 1463.175 3197.800 ;
        RECT 1535.105 3197.755 1535.395 3197.800 ;
        RECT 1559.485 3197.940 1559.775 3197.985 ;
        RECT 1628.945 3197.940 1629.235 3197.985 ;
        RECT 1559.485 3197.800 1629.235 3197.940 ;
        RECT 1559.485 3197.755 1559.775 3197.800 ;
        RECT 1628.945 3197.755 1629.235 3197.800 ;
        RECT 1680.005 3197.940 1680.295 3197.985 ;
        RECT 1725.085 3197.940 1725.375 3197.985 ;
        RECT 1680.005 3197.800 1725.375 3197.940 ;
        RECT 1680.005 3197.755 1680.295 3197.800 ;
        RECT 1725.085 3197.755 1725.375 3197.800 ;
        RECT 1772.925 3197.940 1773.215 3197.985 ;
        RECT 1821.685 3197.940 1821.975 3197.985 ;
        RECT 1772.925 3197.800 1821.975 3197.940 ;
        RECT 1772.925 3197.755 1773.215 3197.800 ;
        RECT 1821.685 3197.755 1821.975 3197.800 ;
        RECT 1869.525 3197.940 1869.815 3197.985 ;
        RECT 1918.285 3197.940 1918.575 3197.985 ;
        RECT 1869.525 3197.800 1918.575 3197.940 ;
        RECT 1869.525 3197.755 1869.815 3197.800 ;
        RECT 1918.285 3197.755 1918.575 3197.800 ;
        RECT 1966.125 3197.940 1966.415 3197.985 ;
        RECT 2014.885 3197.940 2015.175 3197.985 ;
        RECT 1966.125 3197.800 2015.175 3197.940 ;
        RECT 1966.125 3197.755 1966.415 3197.800 ;
        RECT 2014.885 3197.755 2015.175 3197.800 ;
        RECT 2062.725 3197.940 2063.015 3197.985 ;
        RECT 2208.085 3197.940 2208.375 3197.985 ;
        RECT 2062.725 3197.800 2208.375 3197.940 ;
        RECT 2062.725 3197.755 2063.015 3197.800 ;
        RECT 2208.085 3197.755 2208.375 3197.800 ;
        RECT 15.710 2193.920 16.030 2193.980 ;
        RECT 39.170 2193.920 39.490 2193.980 ;
        RECT 15.710 2193.780 39.490 2193.920 ;
        RECT 15.710 2193.720 16.030 2193.780 ;
        RECT 39.170 2193.720 39.490 2193.780 ;
      LAYER via ;
        RECT 2285.380 3198.420 2285.640 3198.680 ;
        RECT 39.200 3197.740 39.460 3198.000 ;
        RECT 15.740 2193.720 16.000 2193.980 ;
        RECT 39.200 2193.720 39.460 2193.980 ;
      LAYER met2 ;
        RECT 2285.380 3198.450 2285.640 3198.710 ;
        RECT 2286.680 3198.450 2286.960 3200.000 ;
        RECT 2285.380 3198.390 2286.960 3198.450 ;
        RECT 2285.440 3198.310 2286.960 3198.390 ;
        RECT 39.200 3197.710 39.460 3198.030 ;
        RECT 39.260 2194.010 39.400 3197.710 ;
        RECT 2286.680 3197.600 2286.960 3198.310 ;
        RECT 15.740 2193.690 16.000 2194.010 ;
        RECT 39.200 2193.690 39.460 2194.010 ;
        RECT 15.800 2190.125 15.940 2193.690 ;
        RECT 15.730 2189.755 16.010 2190.125 ;
      LAYER via2 ;
        RECT 15.730 2189.800 16.010 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 15.705 2190.090 16.035 2190.105 ;
        RECT -4.800 2189.790 16.035 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 15.705 2189.775 16.035 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.830 3209.500 26.150 3209.560 ;
        RECT 2325.830 3209.500 2326.150 3209.560 ;
        RECT 25.830 3209.360 2326.150 3209.500 ;
        RECT 25.830 3209.300 26.150 3209.360 ;
        RECT 2325.830 3209.300 2326.150 3209.360 ;
        RECT 13.870 1903.220 14.190 1903.280 ;
        RECT 25.830 1903.220 26.150 1903.280 ;
        RECT 13.870 1903.080 26.150 1903.220 ;
        RECT 13.870 1903.020 14.190 1903.080 ;
        RECT 25.830 1903.020 26.150 1903.080 ;
      LAYER via ;
        RECT 25.860 3209.300 26.120 3209.560 ;
        RECT 2325.860 3209.300 2326.120 3209.560 ;
        RECT 13.900 1903.020 14.160 1903.280 ;
        RECT 25.860 1903.020 26.120 1903.280 ;
      LAYER met2 ;
        RECT 25.860 3209.270 26.120 3209.590 ;
        RECT 2325.860 3209.270 2326.120 3209.590 ;
        RECT 25.920 1903.310 26.060 3209.270 ;
        RECT 2325.920 3200.000 2326.060 3209.270 ;
        RECT 2325.780 3197.600 2326.060 3200.000 ;
        RECT 13.900 1903.165 14.160 1903.310 ;
        RECT 13.890 1902.795 14.170 1903.165 ;
        RECT 25.860 1902.990 26.120 1903.310 ;
      LAYER via2 ;
        RECT 13.890 1902.840 14.170 1903.120 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 13.865 1903.130 14.195 1903.145 ;
        RECT -4.800 1902.830 14.195 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 13.865 1902.815 14.195 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1260.010 3212.220 1260.330 3212.280 ;
        RECT 1317.970 3212.220 1318.290 3212.280 ;
        RECT 1260.010 3212.080 1318.290 3212.220 ;
        RECT 1260.010 3212.020 1260.330 3212.080 ;
        RECT 1317.970 3212.020 1318.290 3212.080 ;
        RECT 1317.970 3199.640 1318.290 3199.700 ;
        RECT 2902.670 3199.640 2902.990 3199.700 ;
        RECT 1317.970 3199.500 2902.990 3199.640 ;
        RECT 1317.970 3199.440 1318.290 3199.500 ;
        RECT 2902.670 3199.440 2902.990 3199.500 ;
      LAYER via ;
        RECT 1260.040 3212.020 1260.300 3212.280 ;
        RECT 1318.000 3212.020 1318.260 3212.280 ;
        RECT 1318.000 3199.440 1318.260 3199.700 ;
        RECT 2902.700 3199.440 2902.960 3199.700 ;
      LAYER met2 ;
        RECT 1260.040 3211.990 1260.300 3212.310 ;
        RECT 1318.000 3211.990 1318.260 3212.310 ;
        RECT 1260.100 3200.000 1260.240 3211.990 ;
        RECT 1259.960 3197.600 1260.240 3200.000 ;
        RECT 1318.060 3199.730 1318.200 3211.990 ;
        RECT 1318.000 3199.410 1318.260 3199.730 ;
        RECT 2902.700 3199.410 2902.960 3199.730 ;
        RECT 2902.760 615.925 2902.900 3199.410 ;
        RECT 2902.690 615.555 2902.970 615.925 ;
      LAYER via2 ;
        RECT 2902.690 615.600 2902.970 615.880 ;
      LAYER met3 ;
        RECT 2902.665 615.890 2902.995 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2902.665 615.590 2924.800 615.890 ;
        RECT 2902.665 615.575 2902.995 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.370 3209.160 25.690 3209.220 ;
        RECT 2365.390 3209.160 2365.710 3209.220 ;
        RECT 25.370 3209.020 2365.710 3209.160 ;
        RECT 25.370 3208.960 25.690 3209.020 ;
        RECT 2365.390 3208.960 2365.710 3209.020 ;
        RECT 13.870 1617.960 14.190 1618.020 ;
        RECT 25.370 1617.960 25.690 1618.020 ;
        RECT 13.870 1617.820 25.690 1617.960 ;
        RECT 13.870 1617.760 14.190 1617.820 ;
        RECT 25.370 1617.760 25.690 1617.820 ;
      LAYER via ;
        RECT 25.400 3208.960 25.660 3209.220 ;
        RECT 2365.420 3208.960 2365.680 3209.220 ;
        RECT 13.900 1617.760 14.160 1618.020 ;
        RECT 25.400 1617.760 25.660 1618.020 ;
      LAYER met2 ;
        RECT 25.400 3208.930 25.660 3209.250 ;
        RECT 2365.420 3208.930 2365.680 3209.250 ;
        RECT 25.460 1618.050 25.600 3208.930 ;
        RECT 2365.480 3200.000 2365.620 3208.930 ;
        RECT 2365.340 3197.600 2365.620 3200.000 ;
        RECT 13.900 1617.730 14.160 1618.050 ;
        RECT 25.400 1617.730 25.660 1618.050 ;
        RECT 13.960 1615.525 14.100 1617.730 ;
        RECT 13.890 1615.155 14.170 1615.525 ;
      LAYER via2 ;
        RECT 13.890 1615.200 14.170 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 13.865 1615.490 14.195 1615.505 ;
        RECT -4.800 1615.190 14.195 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 13.865 1615.175 14.195 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 76.045 3196.425 76.215 3197.275 ;
        RECT 123.885 3196.425 124.055 3197.615 ;
        RECT 138.145 3196.425 138.315 3197.615 ;
        RECT 185.985 3196.425 186.155 3197.615 ;
        RECT 186.445 3196.425 186.615 3197.615 ;
        RECT 234.745 3196.425 234.915 3197.615 ;
        RECT 303.285 3197.275 303.455 3197.615 ;
        RECT 303.285 3197.105 304.375 3197.275 ;
        RECT 338.245 3196.765 338.415 3197.615 ;
        RECT 379.645 3196.425 379.815 3197.615 ;
        RECT 427.485 3196.425 427.655 3197.275 ;
        RECT 434.845 3196.765 435.015 3197.615 ;
        RECT 496.485 3197.275 496.655 3197.615 ;
        RECT 496.485 3197.105 497.575 3197.275 ;
        RECT 531.445 3196.765 531.615 3197.615 ;
        RECT 593.085 3197.275 593.255 3197.615 ;
        RECT 593.085 3197.105 594.175 3197.275 ;
        RECT 628.045 3196.765 628.215 3197.615 ;
        RECT 766.045 3197.445 768.055 3197.615 ;
        RECT 767.885 3197.105 768.055 3197.445 ;
        RECT 717.745 3196.765 718.375 3196.935 ;
        RECT 821.245 3196.765 821.415 3197.615 ;
        RECT 882.885 3197.275 883.055 3197.615 ;
        RECT 882.885 3197.105 883.975 3197.275 ;
        RECT 917.845 3196.765 918.015 3197.615 ;
        RECT 979.485 3197.445 980.115 3197.615 ;
        RECT 979.945 3197.105 980.115 3197.445 ;
        RECT 1062.745 3197.275 1062.915 3197.615 ;
        RECT 1014.445 3196.425 1014.615 3197.275 ;
        RECT 1062.285 3196.425 1062.455 3197.275 ;
        RECT 1062.745 3197.105 1063.375 3197.275 ;
        RECT 1148.305 3197.105 1148.475 3199.315 ;
        RECT 1196.605 3197.785 1196.775 3199.315 ;
        RECT 1259.165 3197.785 1259.335 3199.315 ;
        RECT 1289.525 3197.785 1289.695 3199.315 ;
        RECT 1339.205 3197.785 1339.375 3200.335 ;
        RECT 1386.125 3197.785 1386.295 3200.335 ;
        RECT 1435.805 3197.785 1435.975 3200.675 ;
        RECT 1452.825 3197.785 1452.995 3200.675 ;
        RECT 1535.625 3197.785 1535.795 3201.355 ;
        RECT 1559.085 3197.785 1559.255 3201.355 ;
        RECT 1629.005 3201.015 1629.175 3208.495 ;
        RECT 1629.005 3200.845 1629.635 3201.015 ;
        RECT 1629.465 3197.785 1629.635 3200.845 ;
        RECT 1675.925 3197.785 1676.095 3208.495 ;
        RECT 2208.605 3197.785 2208.775 3203.395 ;
        RECT 2226.085 3197.785 2226.255 3203.395 ;
        RECT 2318.545 3197.785 2318.715 3198.635 ;
        RECT 2366.385 3197.785 2366.555 3198.635 ;
      LAYER mcon ;
        RECT 1629.005 3208.325 1629.175 3208.495 ;
        RECT 1535.625 3201.185 1535.795 3201.355 ;
        RECT 1435.805 3200.505 1435.975 3200.675 ;
        RECT 1339.205 3200.165 1339.375 3200.335 ;
        RECT 1148.305 3199.145 1148.475 3199.315 ;
        RECT 123.885 3197.445 124.055 3197.615 ;
        RECT 76.045 3197.105 76.215 3197.275 ;
        RECT 138.145 3197.445 138.315 3197.615 ;
        RECT 185.985 3197.445 186.155 3197.615 ;
        RECT 186.445 3197.445 186.615 3197.615 ;
        RECT 234.745 3197.445 234.915 3197.615 ;
        RECT 303.285 3197.445 303.455 3197.615 ;
        RECT 338.245 3197.445 338.415 3197.615 ;
        RECT 304.205 3197.105 304.375 3197.275 ;
        RECT 379.645 3197.445 379.815 3197.615 ;
        RECT 434.845 3197.445 435.015 3197.615 ;
        RECT 427.485 3197.105 427.655 3197.275 ;
        RECT 496.485 3197.445 496.655 3197.615 ;
        RECT 531.445 3197.445 531.615 3197.615 ;
        RECT 497.405 3197.105 497.575 3197.275 ;
        RECT 593.085 3197.445 593.255 3197.615 ;
        RECT 628.045 3197.445 628.215 3197.615 ;
        RECT 594.005 3197.105 594.175 3197.275 ;
        RECT 821.245 3197.445 821.415 3197.615 ;
        RECT 882.885 3197.445 883.055 3197.615 ;
        RECT 917.845 3197.445 918.015 3197.615 ;
        RECT 883.805 3197.105 883.975 3197.275 ;
        RECT 718.205 3196.765 718.375 3196.935 ;
        RECT 1062.745 3197.445 1062.915 3197.615 ;
        RECT 1196.605 3199.145 1196.775 3199.315 ;
        RECT 1259.165 3199.145 1259.335 3199.315 ;
        RECT 1289.525 3199.145 1289.695 3199.315 ;
        RECT 1386.125 3200.165 1386.295 3200.335 ;
        RECT 1452.825 3200.505 1452.995 3200.675 ;
        RECT 1559.085 3201.185 1559.255 3201.355 ;
        RECT 1675.925 3208.325 1676.095 3208.495 ;
        RECT 2208.605 3203.225 2208.775 3203.395 ;
        RECT 2226.085 3203.225 2226.255 3203.395 ;
        RECT 2318.545 3198.465 2318.715 3198.635 ;
        RECT 2366.385 3198.465 2366.555 3198.635 ;
        RECT 1014.445 3197.105 1014.615 3197.275 ;
        RECT 1062.285 3197.105 1062.455 3197.275 ;
        RECT 1063.205 3197.105 1063.375 3197.275 ;
      LAYER met1 ;
        RECT 1628.945 3208.480 1629.235 3208.525 ;
        RECT 1675.865 3208.480 1676.155 3208.525 ;
        RECT 1628.945 3208.340 1676.155 3208.480 ;
        RECT 1628.945 3208.295 1629.235 3208.340 ;
        RECT 1675.865 3208.295 1676.155 3208.340 ;
        RECT 2208.545 3203.380 2208.835 3203.425 ;
        RECT 2226.025 3203.380 2226.315 3203.425 ;
        RECT 2208.545 3203.240 2226.315 3203.380 ;
        RECT 2208.545 3203.195 2208.835 3203.240 ;
        RECT 2226.025 3203.195 2226.315 3203.240 ;
        RECT 1535.565 3201.340 1535.855 3201.385 ;
        RECT 1559.025 3201.340 1559.315 3201.385 ;
        RECT 1535.565 3201.200 1559.315 3201.340 ;
        RECT 1535.565 3201.155 1535.855 3201.200 ;
        RECT 1559.025 3201.155 1559.315 3201.200 ;
        RECT 1435.745 3200.660 1436.035 3200.705 ;
        RECT 1452.765 3200.660 1453.055 3200.705 ;
        RECT 1435.745 3200.520 1453.055 3200.660 ;
        RECT 1435.745 3200.475 1436.035 3200.520 ;
        RECT 1452.765 3200.475 1453.055 3200.520 ;
        RECT 1339.145 3200.320 1339.435 3200.365 ;
        RECT 1386.065 3200.320 1386.355 3200.365 ;
        RECT 1339.145 3200.180 1386.355 3200.320 ;
        RECT 1339.145 3200.135 1339.435 3200.180 ;
        RECT 1386.065 3200.135 1386.355 3200.180 ;
        RECT 1148.245 3199.300 1148.535 3199.345 ;
        RECT 1196.545 3199.300 1196.835 3199.345 ;
        RECT 1148.245 3199.160 1196.835 3199.300 ;
        RECT 1148.245 3199.115 1148.535 3199.160 ;
        RECT 1196.545 3199.115 1196.835 3199.160 ;
        RECT 1259.105 3199.300 1259.395 3199.345 ;
        RECT 1289.465 3199.300 1289.755 3199.345 ;
        RECT 1259.105 3199.160 1289.755 3199.300 ;
        RECT 1259.105 3199.115 1259.395 3199.160 ;
        RECT 1289.465 3199.115 1289.755 3199.160 ;
        RECT 2318.485 3198.620 2318.775 3198.665 ;
        RECT 2366.325 3198.620 2366.615 3198.665 ;
        RECT 2318.485 3198.480 2366.615 3198.620 ;
        RECT 2318.485 3198.435 2318.775 3198.480 ;
        RECT 2366.325 3198.435 2366.615 3198.480 ;
        RECT 2403.110 3198.280 2403.430 3198.340 ;
        RECT 2380.200 3198.140 2403.430 3198.280 ;
        RECT 1196.545 3197.755 1196.835 3197.985 ;
        RECT 1259.105 3197.755 1259.395 3197.985 ;
        RECT 1289.465 3197.755 1289.755 3197.985 ;
        RECT 1339.145 3197.755 1339.435 3197.985 ;
        RECT 1386.065 3197.755 1386.355 3197.985 ;
        RECT 1435.745 3197.755 1436.035 3197.985 ;
        RECT 1452.765 3197.755 1453.055 3197.985 ;
        RECT 1535.565 3197.755 1535.855 3197.985 ;
        RECT 1559.025 3197.755 1559.315 3197.985 ;
        RECT 1629.405 3197.755 1629.695 3197.985 ;
        RECT 1675.865 3197.755 1676.155 3197.985 ;
        RECT 1725.620 3197.800 1772.680 3197.940 ;
        RECT 123.825 3197.600 124.115 3197.645 ;
        RECT 138.085 3197.600 138.375 3197.645 ;
        RECT 123.825 3197.460 138.375 3197.600 ;
        RECT 123.825 3197.415 124.115 3197.460 ;
        RECT 138.085 3197.415 138.375 3197.460 ;
        RECT 185.925 3197.600 186.215 3197.645 ;
        RECT 186.385 3197.600 186.675 3197.645 ;
        RECT 185.925 3197.460 186.675 3197.600 ;
        RECT 185.925 3197.415 186.215 3197.460 ;
        RECT 186.385 3197.415 186.675 3197.460 ;
        RECT 234.685 3197.600 234.975 3197.645 ;
        RECT 303.225 3197.600 303.515 3197.645 ;
        RECT 234.685 3197.460 303.515 3197.600 ;
        RECT 234.685 3197.415 234.975 3197.460 ;
        RECT 303.225 3197.415 303.515 3197.460 ;
        RECT 338.185 3197.600 338.475 3197.645 ;
        RECT 379.585 3197.600 379.875 3197.645 ;
        RECT 338.185 3197.460 379.875 3197.600 ;
        RECT 338.185 3197.415 338.475 3197.460 ;
        RECT 379.585 3197.415 379.875 3197.460 ;
        RECT 434.785 3197.600 435.075 3197.645 ;
        RECT 496.425 3197.600 496.715 3197.645 ;
        RECT 434.785 3197.460 496.715 3197.600 ;
        RECT 434.785 3197.415 435.075 3197.460 ;
        RECT 496.425 3197.415 496.715 3197.460 ;
        RECT 531.385 3197.600 531.675 3197.645 ;
        RECT 593.025 3197.600 593.315 3197.645 ;
        RECT 531.385 3197.460 593.315 3197.600 ;
        RECT 531.385 3197.415 531.675 3197.460 ;
        RECT 593.025 3197.415 593.315 3197.460 ;
        RECT 627.985 3197.600 628.275 3197.645 ;
        RECT 765.985 3197.600 766.275 3197.645 ;
        RECT 627.985 3197.460 717.440 3197.600 ;
        RECT 627.985 3197.415 628.275 3197.460 ;
        RECT 31.350 3197.260 31.670 3197.320 ;
        RECT 75.985 3197.260 76.275 3197.305 ;
        RECT 31.350 3197.120 76.275 3197.260 ;
        RECT 31.350 3197.060 31.670 3197.120 ;
        RECT 75.985 3197.075 76.275 3197.120 ;
        RECT 304.145 3197.260 304.435 3197.305 ;
        RECT 427.425 3197.260 427.715 3197.305 ;
        RECT 497.345 3197.260 497.635 3197.305 ;
        RECT 593.945 3197.260 594.235 3197.305 ;
        RECT 717.300 3197.260 717.440 3197.460 ;
        RECT 741.220 3197.460 766.275 3197.600 ;
        RECT 304.145 3197.120 338.400 3197.260 ;
        RECT 304.145 3197.075 304.435 3197.120 ;
        RECT 338.260 3196.965 338.400 3197.120 ;
        RECT 427.425 3197.120 435.000 3197.260 ;
        RECT 427.425 3197.075 427.715 3197.120 ;
        RECT 434.860 3196.965 435.000 3197.120 ;
        RECT 497.345 3197.120 531.600 3197.260 ;
        RECT 497.345 3197.075 497.635 3197.120 ;
        RECT 531.460 3196.965 531.600 3197.120 ;
        RECT 593.945 3197.120 628.200 3197.260 ;
        RECT 717.300 3197.120 717.900 3197.260 ;
        RECT 593.945 3197.075 594.235 3197.120 ;
        RECT 628.060 3196.965 628.200 3197.120 ;
        RECT 717.760 3196.965 717.900 3197.120 ;
        RECT 338.185 3196.735 338.475 3196.965 ;
        RECT 434.785 3196.735 435.075 3196.965 ;
        RECT 531.385 3196.735 531.675 3196.965 ;
        RECT 627.985 3196.735 628.275 3196.965 ;
        RECT 717.685 3196.735 717.975 3196.965 ;
        RECT 718.145 3196.920 718.435 3196.965 ;
        RECT 741.220 3196.920 741.360 3197.460 ;
        RECT 765.985 3197.415 766.275 3197.460 ;
        RECT 821.185 3197.600 821.475 3197.645 ;
        RECT 882.825 3197.600 883.115 3197.645 ;
        RECT 821.185 3197.460 883.115 3197.600 ;
        RECT 821.185 3197.415 821.475 3197.460 ;
        RECT 882.825 3197.415 883.115 3197.460 ;
        RECT 917.785 3197.600 918.075 3197.645 ;
        RECT 979.425 3197.600 979.715 3197.645 ;
        RECT 1062.685 3197.600 1062.975 3197.645 ;
        RECT 917.785 3197.460 979.715 3197.600 ;
        RECT 917.785 3197.415 918.075 3197.460 ;
        RECT 979.425 3197.415 979.715 3197.460 ;
        RECT 1062.300 3197.460 1062.975 3197.600 ;
        RECT 1196.620 3197.600 1196.760 3197.755 ;
        RECT 1259.180 3197.600 1259.320 3197.755 ;
        RECT 1196.620 3197.460 1259.320 3197.600 ;
        RECT 1289.540 3197.600 1289.680 3197.755 ;
        RECT 1339.220 3197.600 1339.360 3197.755 ;
        RECT 1289.540 3197.460 1339.360 3197.600 ;
        RECT 1386.140 3197.600 1386.280 3197.755 ;
        RECT 1435.820 3197.600 1435.960 3197.755 ;
        RECT 1386.140 3197.460 1435.960 3197.600 ;
        RECT 1452.840 3197.600 1452.980 3197.755 ;
        RECT 1535.640 3197.600 1535.780 3197.755 ;
        RECT 1452.840 3197.460 1535.780 3197.600 ;
        RECT 1559.100 3197.600 1559.240 3197.755 ;
        RECT 1629.480 3197.600 1629.620 3197.755 ;
        RECT 1559.100 3197.460 1629.620 3197.600 ;
        RECT 1675.940 3197.600 1676.080 3197.755 ;
        RECT 1725.620 3197.600 1725.760 3197.800 ;
        RECT 1675.940 3197.460 1725.760 3197.600 ;
        RECT 1772.540 3197.600 1772.680 3197.800 ;
        RECT 1824.980 3197.800 1869.280 3197.940 ;
        RECT 1824.980 3197.600 1825.120 3197.800 ;
        RECT 1772.540 3197.460 1825.120 3197.600 ;
        RECT 1869.140 3197.600 1869.280 3197.800 ;
        RECT 1921.580 3197.800 1965.880 3197.940 ;
        RECT 1921.580 3197.600 1921.720 3197.800 ;
        RECT 1869.140 3197.460 1921.720 3197.600 ;
        RECT 1965.740 3197.600 1965.880 3197.800 ;
        RECT 2208.545 3197.755 2208.835 3197.985 ;
        RECT 2226.025 3197.755 2226.315 3197.985 ;
        RECT 2318.485 3197.755 2318.775 3197.985 ;
        RECT 2366.325 3197.940 2366.615 3197.985 ;
        RECT 2380.200 3197.940 2380.340 3198.140 ;
        RECT 2403.110 3198.080 2403.430 3198.140 ;
        RECT 2366.325 3197.800 2380.340 3197.940 ;
        RECT 2366.325 3197.755 2366.615 3197.800 ;
        RECT 2208.620 3197.600 2208.760 3197.755 ;
        RECT 1965.740 3197.460 2208.760 3197.600 ;
        RECT 2226.100 3197.600 2226.240 3197.755 ;
        RECT 2318.560 3197.600 2318.700 3197.755 ;
        RECT 2226.100 3197.460 2318.700 3197.600 ;
        RECT 1062.300 3197.305 1062.440 3197.460 ;
        RECT 1062.685 3197.415 1062.975 3197.460 ;
        RECT 767.825 3197.260 768.115 3197.305 ;
        RECT 883.745 3197.260 884.035 3197.305 ;
        RECT 979.885 3197.260 980.175 3197.305 ;
        RECT 1014.385 3197.260 1014.675 3197.305 ;
        RECT 767.825 3197.120 821.400 3197.260 ;
        RECT 767.825 3197.075 768.115 3197.120 ;
        RECT 821.260 3196.965 821.400 3197.120 ;
        RECT 883.745 3197.120 918.000 3197.260 ;
        RECT 883.745 3197.075 884.035 3197.120 ;
        RECT 917.860 3196.965 918.000 3197.120 ;
        RECT 979.885 3197.120 1014.675 3197.260 ;
        RECT 979.885 3197.075 980.175 3197.120 ;
        RECT 1014.385 3197.075 1014.675 3197.120 ;
        RECT 1062.225 3197.075 1062.515 3197.305 ;
        RECT 1063.145 3197.260 1063.435 3197.305 ;
        RECT 1148.245 3197.260 1148.535 3197.305 ;
        RECT 1063.145 3197.120 1148.535 3197.260 ;
        RECT 1063.145 3197.075 1063.435 3197.120 ;
        RECT 1148.245 3197.075 1148.535 3197.120 ;
        RECT 718.145 3196.780 741.360 3196.920 ;
        RECT 718.145 3196.735 718.435 3196.780 ;
        RECT 821.185 3196.735 821.475 3196.965 ;
        RECT 917.785 3196.735 918.075 3196.965 ;
        RECT 75.985 3196.580 76.275 3196.625 ;
        RECT 123.825 3196.580 124.115 3196.625 ;
        RECT 75.985 3196.440 124.115 3196.580 ;
        RECT 75.985 3196.395 76.275 3196.440 ;
        RECT 123.825 3196.395 124.115 3196.440 ;
        RECT 138.085 3196.580 138.375 3196.625 ;
        RECT 185.925 3196.580 186.215 3196.625 ;
        RECT 138.085 3196.440 186.215 3196.580 ;
        RECT 138.085 3196.395 138.375 3196.440 ;
        RECT 185.925 3196.395 186.215 3196.440 ;
        RECT 186.385 3196.580 186.675 3196.625 ;
        RECT 234.685 3196.580 234.975 3196.625 ;
        RECT 186.385 3196.440 234.975 3196.580 ;
        RECT 186.385 3196.395 186.675 3196.440 ;
        RECT 234.685 3196.395 234.975 3196.440 ;
        RECT 379.585 3196.580 379.875 3196.625 ;
        RECT 427.425 3196.580 427.715 3196.625 ;
        RECT 379.585 3196.440 427.715 3196.580 ;
        RECT 379.585 3196.395 379.875 3196.440 ;
        RECT 427.425 3196.395 427.715 3196.440 ;
        RECT 1014.385 3196.580 1014.675 3196.625 ;
        RECT 1062.225 3196.580 1062.515 3196.625 ;
        RECT 1014.385 3196.440 1062.515 3196.580 ;
        RECT 1014.385 3196.395 1014.675 3196.440 ;
        RECT 1062.225 3196.395 1062.515 3196.440 ;
        RECT 15.710 1400.700 16.030 1400.760 ;
        RECT 31.350 1400.700 31.670 1400.760 ;
        RECT 15.710 1400.560 31.670 1400.700 ;
        RECT 15.710 1400.500 16.030 1400.560 ;
        RECT 31.350 1400.500 31.670 1400.560 ;
      LAYER via ;
        RECT 31.380 3197.060 31.640 3197.320 ;
        RECT 2403.140 3198.080 2403.400 3198.340 ;
        RECT 15.740 1400.500 16.000 1400.760 ;
        RECT 31.380 1400.500 31.640 1400.760 ;
      LAYER met2 ;
        RECT 2404.900 3198.450 2405.180 3200.000 ;
        RECT 2403.200 3198.370 2405.180 3198.450 ;
        RECT 2403.140 3198.310 2405.180 3198.370 ;
        RECT 2403.140 3198.050 2403.400 3198.310 ;
        RECT 2404.900 3197.600 2405.180 3198.310 ;
        RECT 31.380 3197.030 31.640 3197.350 ;
        RECT 31.440 1400.790 31.580 3197.030 ;
        RECT 15.740 1400.645 16.000 1400.790 ;
        RECT 15.730 1400.275 16.010 1400.645 ;
        RECT 31.380 1400.470 31.640 1400.790 ;
      LAYER via2 ;
        RECT 15.730 1400.320 16.010 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 15.705 1400.610 16.035 1400.625 ;
        RECT -4.800 1400.310 16.035 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 15.705 1400.295 16.035 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 24.910 3208.820 25.230 3208.880 ;
        RECT 2444.510 3208.820 2444.830 3208.880 ;
        RECT 24.910 3208.680 2444.830 3208.820 ;
        RECT 24.910 3208.620 25.230 3208.680 ;
        RECT 2444.510 3208.620 2444.830 3208.680 ;
        RECT 13.870 1186.500 14.190 1186.560 ;
        RECT 24.910 1186.500 25.230 1186.560 ;
        RECT 13.870 1186.360 25.230 1186.500 ;
        RECT 13.870 1186.300 14.190 1186.360 ;
        RECT 24.910 1186.300 25.230 1186.360 ;
      LAYER via ;
        RECT 24.940 3208.620 25.200 3208.880 ;
        RECT 2444.540 3208.620 2444.800 3208.880 ;
        RECT 13.900 1186.300 14.160 1186.560 ;
        RECT 24.940 1186.300 25.200 1186.560 ;
      LAYER met2 ;
        RECT 24.940 3208.590 25.200 3208.910 ;
        RECT 2444.540 3208.590 2444.800 3208.910 ;
        RECT 25.000 1186.590 25.140 3208.590 ;
        RECT 2444.600 3200.000 2444.740 3208.590 ;
        RECT 2444.460 3197.600 2444.740 3200.000 ;
        RECT 13.900 1186.270 14.160 1186.590 ;
        RECT 24.940 1186.270 25.200 1186.590 ;
        RECT 13.960 1185.085 14.100 1186.270 ;
        RECT 13.890 1184.715 14.170 1185.085 ;
      LAYER via2 ;
        RECT 13.890 1184.760 14.170 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 13.865 1185.050 14.195 1185.065 ;
        RECT -4.800 1184.750 14.195 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 13.865 1184.735 14.195 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 971.620 16.030 971.680 ;
        RECT 30.890 971.620 31.210 971.680 ;
        RECT 15.710 971.480 31.210 971.620 ;
        RECT 15.710 971.420 16.030 971.480 ;
        RECT 30.890 971.420 31.210 971.480 ;
      LAYER via ;
        RECT 15.740 971.420 16.000 971.680 ;
        RECT 30.920 971.420 31.180 971.680 ;
      LAYER met2 ;
        RECT 2483.170 3198.450 2483.450 3198.565 ;
        RECT 2484.020 3198.450 2484.300 3200.000 ;
        RECT 2483.170 3198.310 2484.300 3198.450 ;
        RECT 2483.170 3198.195 2483.450 3198.310 ;
        RECT 2484.020 3197.600 2484.300 3198.310 ;
        RECT 30.910 3195.475 31.190 3195.845 ;
        RECT 30.980 971.710 31.120 3195.475 ;
        RECT 15.740 971.390 16.000 971.710 ;
        RECT 30.920 971.390 31.180 971.710 ;
        RECT 15.800 969.525 15.940 971.390 ;
        RECT 15.730 969.155 16.010 969.525 ;
      LAYER via2 ;
        RECT 2483.170 3198.240 2483.450 3198.520 ;
        RECT 30.910 3195.520 31.190 3195.800 ;
        RECT 15.730 969.200 16.010 969.480 ;
      LAYER met3 ;
        RECT 2466.790 3198.530 2467.170 3198.540 ;
        RECT 2483.145 3198.530 2483.475 3198.545 ;
        RECT 2466.790 3198.230 2483.475 3198.530 ;
        RECT 2466.790 3198.220 2467.170 3198.230 ;
        RECT 2483.145 3198.215 2483.475 3198.230 ;
        RECT 30.885 3195.810 31.215 3195.825 ;
        RECT 2466.790 3195.810 2467.170 3195.820 ;
        RECT 30.885 3195.510 2467.170 3195.810 ;
        RECT 30.885 3195.495 31.215 3195.510 ;
        RECT 2466.790 3195.500 2467.170 3195.510 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.705 969.490 16.035 969.505 ;
        RECT -4.800 969.190 16.035 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.705 969.175 16.035 969.190 ;
      LAYER via3 ;
        RECT 2466.820 3198.220 2467.140 3198.540 ;
        RECT 2466.820 3195.500 2467.140 3195.820 ;
      LAYER met4 ;
        RECT 2466.815 3198.215 2467.145 3198.545 ;
        RECT 2466.830 3195.825 2467.130 3198.215 ;
        RECT 2466.815 3195.495 2467.145 3195.825 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 3205.080 20.170 3205.140 ;
        RECT 1293.590 3205.080 1293.910 3205.140 ;
        RECT 19.850 3204.940 1293.910 3205.080 ;
        RECT 19.850 3204.880 20.170 3204.940 ;
        RECT 1293.590 3204.880 1293.910 3204.940 ;
      LAYER via ;
        RECT 19.880 3204.880 20.140 3205.140 ;
        RECT 1293.620 3204.880 1293.880 3205.140 ;
      LAYER met2 ;
        RECT 1293.610 3213.835 1293.890 3214.205 ;
        RECT 2523.190 3213.835 2523.470 3214.205 ;
        RECT 1293.680 3205.170 1293.820 3213.835 ;
        RECT 19.880 3204.850 20.140 3205.170 ;
        RECT 1293.620 3204.850 1293.880 3205.170 ;
        RECT 19.940 753.965 20.080 3204.850 ;
        RECT 2523.260 3200.000 2523.400 3213.835 ;
        RECT 2523.120 3197.600 2523.400 3200.000 ;
        RECT 19.870 753.595 20.150 753.965 ;
      LAYER via2 ;
        RECT 1293.610 3213.880 1293.890 3214.160 ;
        RECT 2523.190 3213.880 2523.470 3214.160 ;
        RECT 19.870 753.640 20.150 753.920 ;
      LAYER met3 ;
        RECT 1293.585 3214.170 1293.915 3214.185 ;
        RECT 2523.165 3214.170 2523.495 3214.185 ;
        RECT 1293.585 3213.870 2523.495 3214.170 ;
        RECT 1293.585 3213.855 1293.915 3213.870 ;
        RECT 2523.165 3213.855 2523.495 3213.870 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 19.845 753.930 20.175 753.945 ;
        RECT -4.800 753.630 20.175 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 19.845 753.615 20.175 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2561.370 3198.450 2561.650 3198.565 ;
        RECT 2562.680 3198.450 2562.960 3200.000 ;
        RECT 2561.370 3198.310 2562.960 3198.450 ;
        RECT 2561.370 3198.195 2561.650 3198.310 ;
        RECT 2562.680 3197.600 2562.960 3198.310 ;
        RECT 18.030 3194.795 18.310 3195.165 ;
        RECT 18.100 538.405 18.240 3194.795 ;
        RECT 18.030 538.035 18.310 538.405 ;
      LAYER via2 ;
        RECT 2561.370 3198.240 2561.650 3198.520 ;
        RECT 18.030 3194.840 18.310 3195.120 ;
        RECT 18.030 538.080 18.310 538.360 ;
      LAYER met3 ;
        RECT 2545.910 3198.530 2546.290 3198.540 ;
        RECT 2561.345 3198.530 2561.675 3198.545 ;
        RECT 2545.910 3198.230 2561.675 3198.530 ;
        RECT 2545.910 3198.220 2546.290 3198.230 ;
        RECT 2561.345 3198.215 2561.675 3198.230 ;
        RECT 18.005 3195.130 18.335 3195.145 ;
        RECT 2545.910 3195.130 2546.290 3195.140 ;
        RECT 18.005 3194.830 2546.290 3195.130 ;
        RECT 18.005 3194.815 18.335 3194.830 ;
        RECT 2545.910 3194.820 2546.290 3194.830 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 18.005 538.370 18.335 538.385 ;
        RECT -4.800 538.070 18.335 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 18.005 538.055 18.335 538.070 ;
      LAYER via3 ;
        RECT 2545.940 3198.220 2546.260 3198.540 ;
        RECT 2545.940 3194.820 2546.260 3195.140 ;
      LAYER met4 ;
        RECT 2545.935 3198.215 2546.265 3198.545 ;
        RECT 2545.950 3195.145 2546.250 3198.215 ;
        RECT 2545.935 3194.815 2546.265 3195.145 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 3215.195 17.850 3215.565 ;
        RECT 2602.310 3215.195 2602.590 3215.565 ;
        RECT 17.640 322.845 17.780 3215.195 ;
        RECT 2602.380 3200.000 2602.520 3215.195 ;
        RECT 2602.240 3197.600 2602.520 3200.000 ;
        RECT 17.570 322.475 17.850 322.845 ;
      LAYER via2 ;
        RECT 17.570 3215.240 17.850 3215.520 ;
        RECT 2602.310 3215.240 2602.590 3215.520 ;
        RECT 17.570 322.520 17.850 322.800 ;
      LAYER met3 ;
        RECT 17.545 3215.530 17.875 3215.545 ;
        RECT 2602.285 3215.530 2602.615 3215.545 ;
        RECT 17.545 3215.230 2602.615 3215.530 ;
        RECT 17.545 3215.215 17.875 3215.230 ;
        RECT 2602.285 3215.215 2602.615 3215.230 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 17.545 322.810 17.875 322.825 ;
        RECT -4.800 322.510 17.875 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 17.545 322.495 17.875 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2640.490 3198.450 2640.770 3198.565 ;
        RECT 2641.800 3198.450 2642.080 3200.000 ;
        RECT 2640.490 3198.310 2642.080 3198.450 ;
        RECT 2640.490 3198.195 2640.770 3198.310 ;
        RECT 2641.800 3197.600 2642.080 3198.310 ;
        RECT 2637.270 1682.475 2637.550 1682.845 ;
        RECT 2637.340 1595.125 2637.480 1682.475 ;
        RECT 2637.270 1594.755 2637.550 1595.125 ;
        RECT 2638.190 1545.115 2638.470 1545.485 ;
        RECT 2638.260 1510.805 2638.400 1545.115 ;
        RECT 2638.190 1510.435 2638.470 1510.805 ;
        RECT 2638.190 1448.555 2638.470 1448.925 ;
        RECT 2638.260 1402.005 2638.400 1448.555 ;
        RECT 2638.190 1401.635 2638.470 1402.005 ;
        RECT 2637.270 1351.995 2637.550 1352.365 ;
        RECT 2637.340 1305.445 2637.480 1351.995 ;
        RECT 2637.270 1305.075 2637.550 1305.445 ;
        RECT 2637.270 1255.435 2637.550 1255.805 ;
        RECT 2637.340 1208.885 2637.480 1255.435 ;
        RECT 2637.270 1208.515 2637.550 1208.885 ;
        RECT 2638.190 1158.875 2638.470 1159.245 ;
        RECT 2638.260 1111.645 2638.400 1158.875 ;
        RECT 2638.190 1111.275 2638.470 1111.645 ;
        RECT 2637.270 1062.315 2637.550 1062.685 ;
        RECT 2637.340 1015.765 2637.480 1062.315 ;
        RECT 2637.270 1015.395 2637.550 1015.765 ;
        RECT 2637.270 965.755 2637.550 966.125 ;
        RECT 2637.340 919.205 2637.480 965.755 ;
        RECT 2637.270 918.835 2637.550 919.205 ;
        RECT 2636.350 869.195 2636.630 869.565 ;
        RECT 2636.420 821.285 2636.560 869.195 ;
        RECT 2636.350 820.915 2636.630 821.285 ;
        RECT 2636.350 771.275 2636.630 771.645 ;
        RECT 2636.420 724.725 2636.560 771.275 ;
        RECT 2636.350 724.355 2636.630 724.725 ;
        RECT 2639.110 675.395 2639.390 675.765 ;
        RECT 2639.180 628.165 2639.320 675.395 ;
        RECT 2639.110 627.795 2639.390 628.165 ;
        RECT 2637.270 482.275 2637.550 482.645 ;
        RECT 2637.340 435.045 2637.480 482.275 ;
        RECT 2637.270 434.675 2637.550 435.045 ;
        RECT 2636.350 288.475 2636.630 288.845 ;
        RECT 2636.420 241.925 2636.560 288.475 ;
        RECT 2636.350 241.555 2636.630 241.925 ;
        RECT 2637.270 192.595 2637.550 192.965 ;
        RECT 2637.340 146.045 2637.480 192.595 ;
        RECT 2637.270 145.675 2637.550 146.045 ;
        RECT 2608.290 110.995 2608.570 111.365 ;
        RECT 2608.360 110.005 2608.500 110.995 ;
        RECT 2608.290 109.635 2608.570 110.005 ;
      LAYER via2 ;
        RECT 2640.490 3198.240 2640.770 3198.520 ;
        RECT 2637.270 1682.520 2637.550 1682.800 ;
        RECT 2637.270 1594.800 2637.550 1595.080 ;
        RECT 2638.190 1545.160 2638.470 1545.440 ;
        RECT 2638.190 1510.480 2638.470 1510.760 ;
        RECT 2638.190 1448.600 2638.470 1448.880 ;
        RECT 2638.190 1401.680 2638.470 1401.960 ;
        RECT 2637.270 1352.040 2637.550 1352.320 ;
        RECT 2637.270 1305.120 2637.550 1305.400 ;
        RECT 2637.270 1255.480 2637.550 1255.760 ;
        RECT 2637.270 1208.560 2637.550 1208.840 ;
        RECT 2638.190 1158.920 2638.470 1159.200 ;
        RECT 2638.190 1111.320 2638.470 1111.600 ;
        RECT 2637.270 1062.360 2637.550 1062.640 ;
        RECT 2637.270 1015.440 2637.550 1015.720 ;
        RECT 2637.270 965.800 2637.550 966.080 ;
        RECT 2637.270 918.880 2637.550 919.160 ;
        RECT 2636.350 869.240 2636.630 869.520 ;
        RECT 2636.350 820.960 2636.630 821.240 ;
        RECT 2636.350 771.320 2636.630 771.600 ;
        RECT 2636.350 724.400 2636.630 724.680 ;
        RECT 2639.110 675.440 2639.390 675.720 ;
        RECT 2639.110 627.840 2639.390 628.120 ;
        RECT 2637.270 482.320 2637.550 482.600 ;
        RECT 2637.270 434.720 2637.550 435.000 ;
        RECT 2636.350 288.520 2636.630 288.800 ;
        RECT 2636.350 241.600 2636.630 241.880 ;
        RECT 2637.270 192.640 2637.550 192.920 ;
        RECT 2637.270 145.720 2637.550 146.000 ;
        RECT 2608.290 111.040 2608.570 111.320 ;
        RECT 2608.290 109.680 2608.570 109.960 ;
      LAYER met3 ;
        RECT 2636.990 3198.530 2637.370 3198.540 ;
        RECT 2640.465 3198.530 2640.795 3198.545 ;
        RECT 2636.990 3198.230 2640.795 3198.530 ;
        RECT 2636.990 3198.220 2637.370 3198.230 ;
        RECT 2640.465 3198.215 2640.795 3198.230 ;
        RECT 2636.990 3171.330 2637.370 3171.340 ;
        RECT 2636.110 3171.030 2637.370 3171.330 ;
        RECT 2636.110 3169.980 2636.410 3171.030 ;
        RECT 2636.990 3171.020 2637.370 3171.030 ;
        RECT 2636.070 3169.660 2636.450 3169.980 ;
        RECT 2636.070 3115.570 2636.450 3115.580 ;
        RECT 2640.670 3115.570 2641.050 3115.580 ;
        RECT 2636.070 3115.270 2641.050 3115.570 ;
        RECT 2636.070 3115.260 2636.450 3115.270 ;
        RECT 2640.670 3115.260 2641.050 3115.270 ;
        RECT 2640.670 3091.090 2641.050 3091.100 ;
        RECT 2643.430 3091.090 2643.810 3091.100 ;
        RECT 2640.670 3090.790 2643.810 3091.090 ;
        RECT 2640.670 3090.780 2641.050 3090.790 ;
        RECT 2643.430 3090.780 2643.810 3090.790 ;
        RECT 2641.590 3043.490 2641.970 3043.500 ;
        RECT 2643.430 3043.490 2643.810 3043.500 ;
        RECT 2641.590 3043.190 2643.810 3043.490 ;
        RECT 2641.590 3043.180 2641.970 3043.190 ;
        RECT 2643.430 3043.180 2643.810 3043.190 ;
        RECT 2637.910 3019.010 2638.290 3019.020 ;
        RECT 2641.590 3019.010 2641.970 3019.020 ;
        RECT 2637.910 3018.710 2641.970 3019.010 ;
        RECT 2637.910 3018.700 2638.290 3018.710 ;
        RECT 2641.590 3018.700 2641.970 3018.710 ;
        RECT 2636.070 2936.050 2636.450 2936.060 ;
        RECT 2639.750 2936.050 2640.130 2936.060 ;
        RECT 2636.070 2935.750 2640.130 2936.050 ;
        RECT 2636.070 2935.740 2636.450 2935.750 ;
        RECT 2639.750 2935.740 2640.130 2935.750 ;
        RECT 2639.750 2897.970 2640.130 2897.980 ;
        RECT 2641.590 2897.970 2641.970 2897.980 ;
        RECT 2639.750 2897.670 2641.970 2897.970 ;
        RECT 2639.750 2897.660 2640.130 2897.670 ;
        RECT 2641.590 2897.660 2641.970 2897.670 ;
        RECT 2641.590 2851.050 2641.970 2851.060 ;
        RECT 2638.870 2850.750 2641.970 2851.050 ;
        RECT 2638.870 2850.380 2639.170 2850.750 ;
        RECT 2641.590 2850.740 2641.970 2850.750 ;
        RECT 2638.830 2850.060 2639.210 2850.380 ;
        RECT 2638.830 2815.380 2639.210 2815.700 ;
        RECT 2638.870 2814.330 2639.170 2815.380 ;
        RECT 2639.750 2814.330 2640.130 2814.340 ;
        RECT 2638.870 2814.030 2640.130 2814.330 ;
        RECT 2639.750 2814.020 2640.130 2814.030 ;
        RECT 2636.990 2801.410 2637.370 2801.420 ;
        RECT 2639.750 2801.410 2640.130 2801.420 ;
        RECT 2636.990 2801.110 2640.130 2801.410 ;
        RECT 2636.990 2801.100 2637.370 2801.110 ;
        RECT 2639.750 2801.100 2640.130 2801.110 ;
        RECT 2636.990 2754.490 2637.370 2754.500 ;
        RECT 2636.990 2754.190 2639.170 2754.490 ;
        RECT 2636.990 2754.180 2637.370 2754.190 ;
        RECT 2638.870 2753.820 2639.170 2754.190 ;
        RECT 2638.830 2753.500 2639.210 2753.820 ;
        RECT 2638.830 2719.810 2639.210 2719.820 ;
        RECT 2636.110 2719.510 2639.210 2719.810 ;
        RECT 2636.110 2717.780 2636.410 2719.510 ;
        RECT 2638.830 2719.500 2639.210 2719.510 ;
        RECT 2636.070 2717.460 2636.450 2717.780 ;
        RECT 2636.070 2670.170 2636.450 2670.180 ;
        RECT 2640.670 2670.170 2641.050 2670.180 ;
        RECT 2636.070 2669.870 2641.050 2670.170 ;
        RECT 2636.070 2669.860 2636.450 2669.870 ;
        RECT 2640.670 2669.860 2641.050 2669.870 ;
        RECT 2640.670 2623.250 2641.050 2623.260 ;
        RECT 2639.790 2622.950 2641.050 2623.250 ;
        RECT 2639.790 2621.220 2640.090 2622.950 ;
        RECT 2640.670 2622.940 2641.050 2622.950 ;
        RECT 2639.750 2620.900 2640.130 2621.220 ;
        RECT 2636.070 2608.290 2636.450 2608.300 ;
        RECT 2639.750 2608.290 2640.130 2608.300 ;
        RECT 2636.070 2607.990 2640.130 2608.290 ;
        RECT 2636.070 2607.980 2636.450 2607.990 ;
        RECT 2639.750 2607.980 2640.130 2607.990 ;
        RECT 2636.070 2561.370 2636.450 2561.380 ;
        RECT 2636.070 2561.070 2638.250 2561.370 ;
        RECT 2636.070 2561.060 2636.450 2561.070 ;
        RECT 2637.950 2560.700 2638.250 2561.070 ;
        RECT 2637.910 2560.380 2638.290 2560.700 ;
        RECT 2637.910 2525.700 2638.290 2526.020 ;
        RECT 2637.950 2524.650 2638.250 2525.700 ;
        RECT 2638.830 2524.650 2639.210 2524.660 ;
        RECT 2637.950 2524.350 2639.210 2524.650 ;
        RECT 2638.830 2524.340 2639.210 2524.350 ;
        RECT 2636.990 2511.730 2637.370 2511.740 ;
        RECT 2638.830 2511.730 2639.210 2511.740 ;
        RECT 2636.990 2511.430 2639.210 2511.730 ;
        RECT 2636.990 2511.420 2637.370 2511.430 ;
        RECT 2638.830 2511.420 2639.210 2511.430 ;
        RECT 2636.990 2463.450 2637.370 2463.460 ;
        RECT 2639.750 2463.450 2640.130 2463.460 ;
        RECT 2636.990 2463.150 2640.130 2463.450 ;
        RECT 2636.990 2463.140 2637.370 2463.150 ;
        RECT 2639.750 2463.140 2640.130 2463.150 ;
        RECT 2639.750 2429.450 2640.130 2429.460 ;
        RECT 2638.870 2429.150 2640.130 2429.450 ;
        RECT 2638.870 2428.100 2639.170 2429.150 ;
        RECT 2639.750 2429.140 2640.130 2429.150 ;
        RECT 2638.830 2427.780 2639.210 2428.100 ;
        RECT 2638.830 2414.490 2639.210 2414.500 ;
        RECT 2640.670 2414.490 2641.050 2414.500 ;
        RECT 2638.830 2414.190 2641.050 2414.490 ;
        RECT 2638.830 2414.180 2639.210 2414.190 ;
        RECT 2640.670 2414.180 2641.050 2414.190 ;
        RECT 2637.910 2366.890 2638.290 2366.900 ;
        RECT 2640.670 2366.890 2641.050 2366.900 ;
        RECT 2637.910 2366.590 2641.050 2366.890 ;
        RECT 2637.910 2366.580 2638.290 2366.590 ;
        RECT 2640.670 2366.580 2641.050 2366.590 ;
        RECT 2636.070 2331.530 2636.450 2331.540 ;
        RECT 2637.910 2331.530 2638.290 2331.540 ;
        RECT 2636.070 2331.230 2638.290 2331.530 ;
        RECT 2636.070 2331.220 2636.450 2331.230 ;
        RECT 2637.910 2331.220 2638.290 2331.230 ;
        RECT 2636.070 2283.930 2636.450 2283.940 ;
        RECT 2638.830 2283.930 2639.210 2283.940 ;
        RECT 2636.070 2283.630 2639.210 2283.930 ;
        RECT 2636.070 2283.620 2636.450 2283.630 ;
        RECT 2638.830 2283.620 2639.210 2283.630 ;
        RECT 2636.070 2222.050 2636.450 2222.060 ;
        RECT 2637.910 2222.050 2638.290 2222.060 ;
        RECT 2636.070 2221.750 2638.290 2222.050 ;
        RECT 2636.070 2221.740 2636.450 2221.750 ;
        RECT 2637.910 2221.740 2638.290 2221.750 ;
        RECT 2636.070 2187.370 2636.450 2187.380 ;
        RECT 2639.750 2187.370 2640.130 2187.380 ;
        RECT 2636.070 2187.070 2640.130 2187.370 ;
        RECT 2636.070 2187.060 2636.450 2187.070 ;
        RECT 2639.750 2187.060 2640.130 2187.070 ;
        RECT 2639.750 2139.770 2640.130 2139.780 ;
        RECT 2638.870 2139.470 2640.130 2139.770 ;
        RECT 2638.870 2138.420 2639.170 2139.470 ;
        RECT 2639.750 2139.460 2640.130 2139.470 ;
        RECT 2638.830 2138.100 2639.210 2138.420 ;
        RECT 2638.830 2124.500 2639.210 2124.820 ;
        RECT 2636.990 2124.130 2637.370 2124.140 ;
        RECT 2638.870 2124.130 2639.170 2124.500 ;
        RECT 2636.990 2123.830 2639.170 2124.130 ;
        RECT 2636.990 2123.820 2637.370 2123.830 ;
        RECT 2636.990 2077.210 2637.370 2077.220 ;
        RECT 2639.750 2077.210 2640.130 2077.220 ;
        RECT 2636.990 2076.910 2640.130 2077.210 ;
        RECT 2636.990 2076.900 2637.370 2076.910 ;
        RECT 2639.750 2076.900 2640.130 2076.910 ;
        RECT 2639.750 2043.210 2640.130 2043.220 ;
        RECT 2638.870 2042.910 2640.130 2043.210 ;
        RECT 2638.870 2041.860 2639.170 2042.910 ;
        RECT 2639.750 2042.900 2640.130 2042.910 ;
        RECT 2638.830 2041.540 2639.210 2041.860 ;
        RECT 2636.070 2028.250 2636.450 2028.260 ;
        RECT 2638.830 2028.250 2639.210 2028.260 ;
        RECT 2636.070 2027.950 2639.210 2028.250 ;
        RECT 2636.070 2027.940 2636.450 2027.950 ;
        RECT 2638.830 2027.940 2639.210 2027.950 ;
        RECT 2636.070 1980.650 2636.450 1980.660 ;
        RECT 2637.910 1980.650 2638.290 1980.660 ;
        RECT 2636.070 1980.350 2638.290 1980.650 ;
        RECT 2636.070 1980.340 2636.450 1980.350 ;
        RECT 2637.910 1980.340 2638.290 1980.350 ;
        RECT 2637.910 1946.650 2638.290 1946.660 ;
        RECT 2637.030 1946.350 2638.290 1946.650 ;
        RECT 2637.030 1945.300 2637.330 1946.350 ;
        RECT 2637.910 1946.340 2638.290 1946.350 ;
        RECT 2636.990 1944.980 2637.370 1945.300 ;
        RECT 2636.990 1931.380 2637.370 1931.700 ;
        RECT 2637.030 1931.010 2637.330 1931.380 ;
        RECT 2639.750 1931.010 2640.130 1931.020 ;
        RECT 2637.030 1930.710 2640.130 1931.010 ;
        RECT 2639.750 1930.700 2640.130 1930.710 ;
        RECT 2637.910 1884.090 2638.290 1884.100 ;
        RECT 2639.750 1884.090 2640.130 1884.100 ;
        RECT 2637.910 1883.790 2640.130 1884.090 ;
        RECT 2637.910 1883.780 2638.290 1883.790 ;
        RECT 2639.750 1883.780 2640.130 1883.790 ;
        RECT 2637.910 1849.780 2638.290 1850.100 ;
        RECT 2637.950 1848.730 2638.250 1849.780 ;
        RECT 2638.830 1848.730 2639.210 1848.740 ;
        RECT 2637.950 1848.430 2639.210 1848.730 ;
        RECT 2638.830 1848.420 2639.210 1848.430 ;
        RECT 2638.830 1834.820 2639.210 1835.140 ;
        RECT 2638.870 1834.450 2639.170 1834.820 ;
        RECT 2641.590 1834.450 2641.970 1834.460 ;
        RECT 2638.870 1834.150 2641.970 1834.450 ;
        RECT 2641.590 1834.140 2641.970 1834.150 ;
        RECT 2639.750 1787.530 2640.130 1787.540 ;
        RECT 2641.590 1787.530 2641.970 1787.540 ;
        RECT 2639.750 1787.230 2641.970 1787.530 ;
        RECT 2639.750 1787.220 2640.130 1787.230 ;
        RECT 2641.590 1787.220 2641.970 1787.230 ;
        RECT 2639.750 1753.530 2640.130 1753.540 ;
        RECT 2638.870 1753.230 2640.130 1753.530 ;
        RECT 2638.870 1752.180 2639.170 1753.230 ;
        RECT 2639.750 1753.220 2640.130 1753.230 ;
        RECT 2638.830 1751.860 2639.210 1752.180 ;
        RECT 2638.830 1738.570 2639.210 1738.580 ;
        RECT 2641.590 1738.570 2641.970 1738.580 ;
        RECT 2638.830 1738.270 2641.970 1738.570 ;
        RECT 2638.830 1738.260 2639.210 1738.270 ;
        RECT 2641.590 1738.260 2641.970 1738.270 ;
        RECT 2637.910 1701.850 2638.290 1701.860 ;
        RECT 2641.590 1701.850 2641.970 1701.860 ;
        RECT 2637.910 1701.550 2641.970 1701.850 ;
        RECT 2637.910 1701.540 2638.290 1701.550 ;
        RECT 2641.590 1701.540 2641.970 1701.550 ;
        RECT 2637.910 1683.180 2638.290 1683.500 ;
        RECT 2637.245 1682.810 2637.575 1682.825 ;
        RECT 2637.950 1682.810 2638.250 1683.180 ;
        RECT 2637.245 1682.510 2638.250 1682.810 ;
        RECT 2637.245 1682.495 2637.575 1682.510 ;
        RECT 2637.245 1595.090 2637.575 1595.105 ;
        RECT 2637.030 1594.775 2637.575 1595.090 ;
        RECT 2637.030 1594.420 2637.330 1594.775 ;
        RECT 2636.990 1594.100 2637.370 1594.420 ;
        RECT 2636.990 1560.100 2637.370 1560.420 ;
        RECT 2637.030 1559.050 2637.330 1560.100 ;
        RECT 2637.910 1559.050 2638.290 1559.060 ;
        RECT 2637.030 1558.750 2638.290 1559.050 ;
        RECT 2637.910 1558.740 2638.290 1558.750 ;
        RECT 2638.165 1545.460 2638.495 1545.465 ;
        RECT 2637.910 1545.450 2638.495 1545.460 ;
        RECT 2637.910 1545.150 2638.720 1545.450 ;
        RECT 2637.910 1545.140 2638.495 1545.150 ;
        RECT 2638.165 1545.135 2638.495 1545.140 ;
        RECT 2636.990 1510.770 2637.370 1510.780 ;
        RECT 2638.165 1510.770 2638.495 1510.785 ;
        RECT 2636.990 1510.470 2638.495 1510.770 ;
        RECT 2636.990 1510.460 2637.370 1510.470 ;
        RECT 2638.165 1510.455 2638.495 1510.470 ;
        RECT 2638.165 1448.900 2638.495 1448.905 ;
        RECT 2637.910 1448.890 2638.495 1448.900 ;
        RECT 2637.910 1448.590 2638.720 1448.890 ;
        RECT 2637.910 1448.580 2638.495 1448.590 ;
        RECT 2638.165 1448.575 2638.495 1448.580 ;
        RECT 2638.165 1401.970 2638.495 1401.985 ;
        RECT 2637.030 1401.670 2638.495 1401.970 ;
        RECT 2637.030 1401.300 2637.330 1401.670 ;
        RECT 2638.165 1401.655 2638.495 1401.670 ;
        RECT 2636.990 1400.980 2637.370 1401.300 ;
        RECT 2636.990 1366.980 2637.370 1367.300 ;
        RECT 2637.030 1365.250 2637.330 1366.980 ;
        RECT 2637.910 1365.250 2638.290 1365.260 ;
        RECT 2637.030 1364.950 2638.290 1365.250 ;
        RECT 2637.910 1364.940 2638.290 1364.950 ;
        RECT 2637.245 1352.330 2637.575 1352.345 ;
        RECT 2637.910 1352.330 2638.290 1352.340 ;
        RECT 2637.245 1352.030 2638.290 1352.330 ;
        RECT 2637.245 1352.015 2637.575 1352.030 ;
        RECT 2637.910 1352.020 2638.290 1352.030 ;
        RECT 2637.245 1305.410 2637.575 1305.425 ;
        RECT 2637.030 1305.095 2637.575 1305.410 ;
        RECT 2637.030 1304.740 2637.330 1305.095 ;
        RECT 2636.990 1304.420 2637.370 1304.740 ;
        RECT 2636.990 1269.740 2637.370 1270.060 ;
        RECT 2637.030 1268.690 2637.330 1269.740 ;
        RECT 2637.910 1268.690 2638.290 1268.700 ;
        RECT 2637.030 1268.390 2638.290 1268.690 ;
        RECT 2637.910 1268.380 2638.290 1268.390 ;
        RECT 2637.245 1255.770 2637.575 1255.785 ;
        RECT 2637.910 1255.770 2638.290 1255.780 ;
        RECT 2637.245 1255.470 2638.290 1255.770 ;
        RECT 2637.245 1255.455 2637.575 1255.470 ;
        RECT 2637.910 1255.460 2638.290 1255.470 ;
        RECT 2637.245 1208.850 2637.575 1208.865 ;
        RECT 2637.030 1208.535 2637.575 1208.850 ;
        RECT 2637.030 1208.180 2637.330 1208.535 ;
        RECT 2636.990 1207.860 2637.370 1208.180 ;
        RECT 2636.990 1173.180 2637.370 1173.500 ;
        RECT 2637.030 1172.130 2637.330 1173.180 ;
        RECT 2637.910 1172.130 2638.290 1172.140 ;
        RECT 2637.030 1171.830 2638.290 1172.130 ;
        RECT 2637.910 1171.820 2638.290 1171.830 ;
        RECT 2638.165 1159.220 2638.495 1159.225 ;
        RECT 2637.910 1159.210 2638.495 1159.220 ;
        RECT 2637.710 1158.910 2638.495 1159.210 ;
        RECT 2637.910 1158.900 2638.495 1158.910 ;
        RECT 2638.165 1158.895 2638.495 1158.900 ;
        RECT 2638.165 1111.610 2638.495 1111.625 ;
        RECT 2638.830 1111.610 2639.210 1111.620 ;
        RECT 2638.165 1111.310 2639.210 1111.610 ;
        RECT 2638.165 1111.295 2638.495 1111.310 ;
        RECT 2638.830 1111.300 2639.210 1111.310 ;
        RECT 2638.830 1077.610 2639.210 1077.620 ;
        RECT 2637.950 1077.310 2639.210 1077.610 ;
        RECT 2637.950 1076.260 2638.250 1077.310 ;
        RECT 2638.830 1077.300 2639.210 1077.310 ;
        RECT 2637.910 1075.940 2638.290 1076.260 ;
        RECT 2637.245 1062.650 2637.575 1062.665 ;
        RECT 2637.910 1062.650 2638.290 1062.660 ;
        RECT 2637.245 1062.350 2638.290 1062.650 ;
        RECT 2637.245 1062.335 2637.575 1062.350 ;
        RECT 2637.910 1062.340 2638.290 1062.350 ;
        RECT 2637.245 1015.730 2637.575 1015.745 ;
        RECT 2637.030 1015.415 2637.575 1015.730 ;
        RECT 2637.030 1015.060 2637.330 1015.415 ;
        RECT 2636.990 1014.740 2637.370 1015.060 ;
        RECT 2636.990 980.060 2637.370 980.380 ;
        RECT 2637.030 979.010 2637.330 980.060 ;
        RECT 2637.910 979.010 2638.290 979.020 ;
        RECT 2637.030 978.710 2638.290 979.010 ;
        RECT 2637.910 978.700 2638.290 978.710 ;
        RECT 2637.245 966.090 2637.575 966.105 ;
        RECT 2637.910 966.090 2638.290 966.100 ;
        RECT 2637.245 965.790 2638.290 966.090 ;
        RECT 2637.245 965.775 2637.575 965.790 ;
        RECT 2637.910 965.780 2638.290 965.790 ;
        RECT 2637.245 919.170 2637.575 919.185 ;
        RECT 2637.030 918.855 2637.575 919.170 ;
        RECT 2637.030 918.500 2637.330 918.855 ;
        RECT 2636.990 918.180 2637.370 918.500 ;
        RECT 2636.990 883.810 2637.370 883.820 ;
        RECT 2636.110 883.510 2637.370 883.810 ;
        RECT 2636.110 882.460 2636.410 883.510 ;
        RECT 2636.990 883.500 2637.370 883.510 ;
        RECT 2636.070 882.140 2636.450 882.460 ;
        RECT 2636.325 869.540 2636.655 869.545 ;
        RECT 2636.070 869.530 2636.655 869.540 ;
        RECT 2635.870 869.230 2636.655 869.530 ;
        RECT 2636.070 869.220 2636.655 869.230 ;
        RECT 2636.325 869.215 2636.655 869.220 ;
        RECT 2636.325 821.250 2636.655 821.265 ;
        RECT 2636.990 821.250 2637.370 821.260 ;
        RECT 2636.325 820.950 2637.370 821.250 ;
        RECT 2636.325 820.935 2636.655 820.950 ;
        RECT 2636.990 820.940 2637.370 820.950 ;
        RECT 2636.990 787.250 2637.370 787.260 ;
        RECT 2636.110 786.950 2637.370 787.250 ;
        RECT 2636.110 785.900 2636.410 786.950 ;
        RECT 2636.990 786.940 2637.370 786.950 ;
        RECT 2636.070 785.580 2636.450 785.900 ;
        RECT 2636.070 771.980 2636.450 772.300 ;
        RECT 2636.110 771.625 2636.410 771.980 ;
        RECT 2636.110 771.310 2636.655 771.625 ;
        RECT 2636.325 771.295 2636.655 771.310 ;
        RECT 2636.325 724.690 2636.655 724.705 ;
        RECT 2636.990 724.690 2637.370 724.700 ;
        RECT 2636.325 724.390 2637.370 724.690 ;
        RECT 2636.325 724.375 2636.655 724.390 ;
        RECT 2636.990 724.380 2637.370 724.390 ;
        RECT 2636.990 700.210 2637.370 700.220 ;
        RECT 2638.830 700.210 2639.210 700.220 ;
        RECT 2636.990 699.910 2639.210 700.210 ;
        RECT 2636.990 699.900 2637.370 699.910 ;
        RECT 2638.830 699.900 2639.210 699.910 ;
        RECT 2639.085 675.740 2639.415 675.745 ;
        RECT 2638.830 675.730 2639.415 675.740 ;
        RECT 2638.830 675.430 2639.640 675.730 ;
        RECT 2638.830 675.420 2639.415 675.430 ;
        RECT 2639.085 675.415 2639.415 675.420 ;
        RECT 2636.990 628.130 2637.370 628.140 ;
        RECT 2639.085 628.130 2639.415 628.145 ;
        RECT 2636.990 627.830 2639.415 628.130 ;
        RECT 2636.990 627.820 2637.370 627.830 ;
        RECT 2639.085 627.815 2639.415 627.830 ;
        RECT 2636.990 593.820 2637.370 594.140 ;
        RECT 2637.030 592.770 2637.330 593.820 ;
        RECT 2637.910 592.770 2638.290 592.780 ;
        RECT 2637.030 592.470 2638.290 592.770 ;
        RECT 2637.910 592.460 2638.290 592.470 ;
        RECT 2636.070 545.170 2636.450 545.180 ;
        RECT 2638.830 545.170 2639.210 545.180 ;
        RECT 2636.070 544.870 2639.210 545.170 ;
        RECT 2636.070 544.860 2636.450 544.870 ;
        RECT 2638.830 544.860 2639.210 544.870 ;
        RECT 2638.830 497.570 2639.210 497.580 ;
        RECT 2637.950 497.270 2639.210 497.570 ;
        RECT 2637.950 496.220 2638.250 497.270 ;
        RECT 2638.830 497.260 2639.210 497.270 ;
        RECT 2637.910 495.900 2638.290 496.220 ;
        RECT 2637.245 482.610 2637.575 482.625 ;
        RECT 2637.910 482.610 2638.290 482.620 ;
        RECT 2637.245 482.310 2638.290 482.610 ;
        RECT 2637.245 482.295 2637.575 482.310 ;
        RECT 2637.910 482.300 2638.290 482.310 ;
        RECT 2637.245 435.020 2637.575 435.025 ;
        RECT 2636.990 435.010 2637.575 435.020 ;
        RECT 2636.790 434.710 2637.575 435.010 ;
        RECT 2636.990 434.700 2637.575 434.710 ;
        RECT 2637.245 434.695 2637.575 434.700 ;
        RECT 2636.990 401.010 2637.370 401.020 ;
        RECT 2636.110 400.710 2637.370 401.010 ;
        RECT 2636.110 399.660 2636.410 400.710 ;
        RECT 2636.990 400.700 2637.370 400.710 ;
        RECT 2636.070 399.340 2636.450 399.660 ;
        RECT 2636.070 352.420 2636.450 352.740 ;
        RECT 2636.110 351.370 2636.410 352.420 ;
        RECT 2637.910 351.370 2638.290 351.380 ;
        RECT 2636.110 351.070 2638.290 351.370 ;
        RECT 2637.910 351.060 2638.290 351.070 ;
        RECT 2636.070 313.970 2636.450 313.980 ;
        RECT 2638.830 313.970 2639.210 313.980 ;
        RECT 2636.070 313.670 2639.210 313.970 ;
        RECT 2636.070 313.660 2636.450 313.670 ;
        RECT 2638.830 313.660 2639.210 313.670 ;
        RECT 2636.070 289.180 2636.450 289.500 ;
        RECT 2636.110 288.825 2636.410 289.180 ;
        RECT 2636.110 288.510 2636.655 288.825 ;
        RECT 2636.325 288.495 2636.655 288.510 ;
        RECT 2636.325 241.890 2636.655 241.905 ;
        RECT 2636.990 241.890 2637.370 241.900 ;
        RECT 2636.325 241.590 2637.370 241.890 ;
        RECT 2636.325 241.575 2636.655 241.590 ;
        RECT 2636.990 241.580 2637.370 241.590 ;
        RECT 2636.990 207.580 2637.370 207.900 ;
        RECT 2637.030 206.530 2637.330 207.580 ;
        RECT 2637.910 206.530 2638.290 206.540 ;
        RECT 2637.030 206.230 2638.290 206.530 ;
        RECT 2637.910 206.220 2638.290 206.230 ;
        RECT 2637.245 192.930 2637.575 192.945 ;
        RECT 2637.910 192.930 2638.290 192.940 ;
        RECT 2637.245 192.630 2638.290 192.930 ;
        RECT 2637.245 192.615 2637.575 192.630 ;
        RECT 2637.910 192.620 2638.290 192.630 ;
        RECT 2637.245 146.010 2637.575 146.025 ;
        RECT 2637.030 145.695 2637.575 146.010 ;
        RECT 2637.030 145.340 2637.330 145.695 ;
        RECT 2636.990 145.020 2637.370 145.340 ;
        RECT 2608.265 111.330 2608.595 111.345 ;
        RECT 2636.990 111.330 2637.370 111.340 ;
        RECT 2608.265 111.030 2637.370 111.330 ;
        RECT 2608.265 111.015 2608.595 111.030 ;
        RECT 2636.990 111.020 2637.370 111.030 ;
        RECT 2608.265 109.970 2608.595 109.985 ;
        RECT 3.070 109.670 2608.595 109.970 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 3.070 107.250 3.370 109.670 ;
        RECT 2608.265 109.655 2608.595 109.670 ;
        RECT -4.800 106.950 3.370 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
      LAYER via3 ;
        RECT 2637.020 3198.220 2637.340 3198.540 ;
        RECT 2637.020 3171.020 2637.340 3171.340 ;
        RECT 2636.100 3169.660 2636.420 3169.980 ;
        RECT 2636.100 3115.260 2636.420 3115.580 ;
        RECT 2640.700 3115.260 2641.020 3115.580 ;
        RECT 2640.700 3090.780 2641.020 3091.100 ;
        RECT 2643.460 3090.780 2643.780 3091.100 ;
        RECT 2641.620 3043.180 2641.940 3043.500 ;
        RECT 2643.460 3043.180 2643.780 3043.500 ;
        RECT 2637.940 3018.700 2638.260 3019.020 ;
        RECT 2641.620 3018.700 2641.940 3019.020 ;
        RECT 2636.100 2935.740 2636.420 2936.060 ;
        RECT 2639.780 2935.740 2640.100 2936.060 ;
        RECT 2639.780 2897.660 2640.100 2897.980 ;
        RECT 2641.620 2897.660 2641.940 2897.980 ;
        RECT 2641.620 2850.740 2641.940 2851.060 ;
        RECT 2638.860 2850.060 2639.180 2850.380 ;
        RECT 2638.860 2815.380 2639.180 2815.700 ;
        RECT 2639.780 2814.020 2640.100 2814.340 ;
        RECT 2637.020 2801.100 2637.340 2801.420 ;
        RECT 2639.780 2801.100 2640.100 2801.420 ;
        RECT 2637.020 2754.180 2637.340 2754.500 ;
        RECT 2638.860 2753.500 2639.180 2753.820 ;
        RECT 2638.860 2719.500 2639.180 2719.820 ;
        RECT 2636.100 2717.460 2636.420 2717.780 ;
        RECT 2636.100 2669.860 2636.420 2670.180 ;
        RECT 2640.700 2669.860 2641.020 2670.180 ;
        RECT 2640.700 2622.940 2641.020 2623.260 ;
        RECT 2639.780 2620.900 2640.100 2621.220 ;
        RECT 2636.100 2607.980 2636.420 2608.300 ;
        RECT 2639.780 2607.980 2640.100 2608.300 ;
        RECT 2636.100 2561.060 2636.420 2561.380 ;
        RECT 2637.940 2560.380 2638.260 2560.700 ;
        RECT 2637.940 2525.700 2638.260 2526.020 ;
        RECT 2638.860 2524.340 2639.180 2524.660 ;
        RECT 2637.020 2511.420 2637.340 2511.740 ;
        RECT 2638.860 2511.420 2639.180 2511.740 ;
        RECT 2637.020 2463.140 2637.340 2463.460 ;
        RECT 2639.780 2463.140 2640.100 2463.460 ;
        RECT 2639.780 2429.140 2640.100 2429.460 ;
        RECT 2638.860 2427.780 2639.180 2428.100 ;
        RECT 2638.860 2414.180 2639.180 2414.500 ;
        RECT 2640.700 2414.180 2641.020 2414.500 ;
        RECT 2637.940 2366.580 2638.260 2366.900 ;
        RECT 2640.700 2366.580 2641.020 2366.900 ;
        RECT 2636.100 2331.220 2636.420 2331.540 ;
        RECT 2637.940 2331.220 2638.260 2331.540 ;
        RECT 2636.100 2283.620 2636.420 2283.940 ;
        RECT 2638.860 2283.620 2639.180 2283.940 ;
        RECT 2636.100 2221.740 2636.420 2222.060 ;
        RECT 2637.940 2221.740 2638.260 2222.060 ;
        RECT 2636.100 2187.060 2636.420 2187.380 ;
        RECT 2639.780 2187.060 2640.100 2187.380 ;
        RECT 2639.780 2139.460 2640.100 2139.780 ;
        RECT 2638.860 2138.100 2639.180 2138.420 ;
        RECT 2638.860 2124.500 2639.180 2124.820 ;
        RECT 2637.020 2123.820 2637.340 2124.140 ;
        RECT 2637.020 2076.900 2637.340 2077.220 ;
        RECT 2639.780 2076.900 2640.100 2077.220 ;
        RECT 2639.780 2042.900 2640.100 2043.220 ;
        RECT 2638.860 2041.540 2639.180 2041.860 ;
        RECT 2636.100 2027.940 2636.420 2028.260 ;
        RECT 2638.860 2027.940 2639.180 2028.260 ;
        RECT 2636.100 1980.340 2636.420 1980.660 ;
        RECT 2637.940 1980.340 2638.260 1980.660 ;
        RECT 2637.940 1946.340 2638.260 1946.660 ;
        RECT 2637.020 1944.980 2637.340 1945.300 ;
        RECT 2637.020 1931.380 2637.340 1931.700 ;
        RECT 2639.780 1930.700 2640.100 1931.020 ;
        RECT 2637.940 1883.780 2638.260 1884.100 ;
        RECT 2639.780 1883.780 2640.100 1884.100 ;
        RECT 2637.940 1849.780 2638.260 1850.100 ;
        RECT 2638.860 1848.420 2639.180 1848.740 ;
        RECT 2638.860 1834.820 2639.180 1835.140 ;
        RECT 2641.620 1834.140 2641.940 1834.460 ;
        RECT 2639.780 1787.220 2640.100 1787.540 ;
        RECT 2641.620 1787.220 2641.940 1787.540 ;
        RECT 2639.780 1753.220 2640.100 1753.540 ;
        RECT 2638.860 1751.860 2639.180 1752.180 ;
        RECT 2638.860 1738.260 2639.180 1738.580 ;
        RECT 2641.620 1738.260 2641.940 1738.580 ;
        RECT 2637.940 1701.540 2638.260 1701.860 ;
        RECT 2641.620 1701.540 2641.940 1701.860 ;
        RECT 2637.940 1683.180 2638.260 1683.500 ;
        RECT 2637.020 1594.100 2637.340 1594.420 ;
        RECT 2637.020 1560.100 2637.340 1560.420 ;
        RECT 2637.940 1558.740 2638.260 1559.060 ;
        RECT 2637.940 1545.140 2638.260 1545.460 ;
        RECT 2637.020 1510.460 2637.340 1510.780 ;
        RECT 2637.940 1448.580 2638.260 1448.900 ;
        RECT 2637.020 1400.980 2637.340 1401.300 ;
        RECT 2637.020 1366.980 2637.340 1367.300 ;
        RECT 2637.940 1364.940 2638.260 1365.260 ;
        RECT 2637.940 1352.020 2638.260 1352.340 ;
        RECT 2637.020 1304.420 2637.340 1304.740 ;
        RECT 2637.020 1269.740 2637.340 1270.060 ;
        RECT 2637.940 1268.380 2638.260 1268.700 ;
        RECT 2637.940 1255.460 2638.260 1255.780 ;
        RECT 2637.020 1207.860 2637.340 1208.180 ;
        RECT 2637.020 1173.180 2637.340 1173.500 ;
        RECT 2637.940 1171.820 2638.260 1172.140 ;
        RECT 2637.940 1158.900 2638.260 1159.220 ;
        RECT 2638.860 1111.300 2639.180 1111.620 ;
        RECT 2638.860 1077.300 2639.180 1077.620 ;
        RECT 2637.940 1075.940 2638.260 1076.260 ;
        RECT 2637.940 1062.340 2638.260 1062.660 ;
        RECT 2637.020 1014.740 2637.340 1015.060 ;
        RECT 2637.020 980.060 2637.340 980.380 ;
        RECT 2637.940 978.700 2638.260 979.020 ;
        RECT 2637.940 965.780 2638.260 966.100 ;
        RECT 2637.020 918.180 2637.340 918.500 ;
        RECT 2637.020 883.500 2637.340 883.820 ;
        RECT 2636.100 882.140 2636.420 882.460 ;
        RECT 2636.100 869.220 2636.420 869.540 ;
        RECT 2637.020 820.940 2637.340 821.260 ;
        RECT 2637.020 786.940 2637.340 787.260 ;
        RECT 2636.100 785.580 2636.420 785.900 ;
        RECT 2636.100 771.980 2636.420 772.300 ;
        RECT 2637.020 724.380 2637.340 724.700 ;
        RECT 2637.020 699.900 2637.340 700.220 ;
        RECT 2638.860 699.900 2639.180 700.220 ;
        RECT 2638.860 675.420 2639.180 675.740 ;
        RECT 2637.020 627.820 2637.340 628.140 ;
        RECT 2637.020 593.820 2637.340 594.140 ;
        RECT 2637.940 592.460 2638.260 592.780 ;
        RECT 2636.100 544.860 2636.420 545.180 ;
        RECT 2638.860 544.860 2639.180 545.180 ;
        RECT 2638.860 497.260 2639.180 497.580 ;
        RECT 2637.940 495.900 2638.260 496.220 ;
        RECT 2637.940 482.300 2638.260 482.620 ;
        RECT 2637.020 434.700 2637.340 435.020 ;
        RECT 2637.020 400.700 2637.340 401.020 ;
        RECT 2636.100 399.340 2636.420 399.660 ;
        RECT 2636.100 352.420 2636.420 352.740 ;
        RECT 2637.940 351.060 2638.260 351.380 ;
        RECT 2636.100 313.660 2636.420 313.980 ;
        RECT 2638.860 313.660 2639.180 313.980 ;
        RECT 2636.100 289.180 2636.420 289.500 ;
        RECT 2637.020 241.580 2637.340 241.900 ;
        RECT 2637.020 207.580 2637.340 207.900 ;
        RECT 2637.940 206.220 2638.260 206.540 ;
        RECT 2637.940 192.620 2638.260 192.940 ;
        RECT 2637.020 145.020 2637.340 145.340 ;
        RECT 2637.020 111.020 2637.340 111.340 ;
      LAYER met4 ;
        RECT 2637.015 3198.215 2637.345 3198.545 ;
        RECT 2637.030 3171.345 2637.330 3198.215 ;
        RECT 2637.015 3171.015 2637.345 3171.345 ;
        RECT 2636.095 3169.655 2636.425 3169.985 ;
        RECT 2636.110 3115.585 2636.410 3169.655 ;
        RECT 2636.095 3115.255 2636.425 3115.585 ;
        RECT 2640.695 3115.255 2641.025 3115.585 ;
        RECT 2640.710 3091.105 2641.010 3115.255 ;
        RECT 2640.695 3090.775 2641.025 3091.105 ;
        RECT 2643.455 3090.775 2643.785 3091.105 ;
        RECT 2643.470 3043.505 2643.770 3090.775 ;
        RECT 2641.615 3043.175 2641.945 3043.505 ;
        RECT 2643.455 3043.175 2643.785 3043.505 ;
        RECT 2641.630 3019.025 2641.930 3043.175 ;
        RECT 2637.935 3018.695 2638.265 3019.025 ;
        RECT 2641.615 3018.695 2641.945 3019.025 ;
        RECT 2637.950 2980.250 2638.250 3018.695 ;
        RECT 2636.110 2979.950 2638.250 2980.250 ;
        RECT 2636.110 2936.065 2636.410 2979.950 ;
        RECT 2636.095 2935.735 2636.425 2936.065 ;
        RECT 2639.775 2935.735 2640.105 2936.065 ;
        RECT 2639.790 2897.985 2640.090 2935.735 ;
        RECT 2639.775 2897.655 2640.105 2897.985 ;
        RECT 2641.615 2897.655 2641.945 2897.985 ;
        RECT 2641.630 2851.065 2641.930 2897.655 ;
        RECT 2641.615 2850.735 2641.945 2851.065 ;
        RECT 2638.855 2850.055 2639.185 2850.385 ;
        RECT 2638.870 2815.705 2639.170 2850.055 ;
        RECT 2638.855 2815.375 2639.185 2815.705 ;
        RECT 2639.775 2814.015 2640.105 2814.345 ;
        RECT 2639.790 2801.425 2640.090 2814.015 ;
        RECT 2637.015 2801.095 2637.345 2801.425 ;
        RECT 2639.775 2801.095 2640.105 2801.425 ;
        RECT 2637.030 2754.505 2637.330 2801.095 ;
        RECT 2637.015 2754.175 2637.345 2754.505 ;
        RECT 2638.855 2753.495 2639.185 2753.825 ;
        RECT 2638.870 2719.825 2639.170 2753.495 ;
        RECT 2638.855 2719.495 2639.185 2719.825 ;
        RECT 2636.095 2717.455 2636.425 2717.785 ;
        RECT 2636.110 2670.185 2636.410 2717.455 ;
        RECT 2636.095 2669.855 2636.425 2670.185 ;
        RECT 2640.695 2669.855 2641.025 2670.185 ;
        RECT 2640.710 2623.265 2641.010 2669.855 ;
        RECT 2640.695 2622.935 2641.025 2623.265 ;
        RECT 2639.775 2620.895 2640.105 2621.225 ;
        RECT 2639.790 2608.305 2640.090 2620.895 ;
        RECT 2636.095 2607.975 2636.425 2608.305 ;
        RECT 2639.775 2607.975 2640.105 2608.305 ;
        RECT 2636.110 2561.385 2636.410 2607.975 ;
        RECT 2636.095 2561.055 2636.425 2561.385 ;
        RECT 2637.935 2560.375 2638.265 2560.705 ;
        RECT 2637.950 2526.025 2638.250 2560.375 ;
        RECT 2637.935 2525.695 2638.265 2526.025 ;
        RECT 2638.855 2524.335 2639.185 2524.665 ;
        RECT 2638.870 2511.745 2639.170 2524.335 ;
        RECT 2637.015 2511.415 2637.345 2511.745 ;
        RECT 2638.855 2511.415 2639.185 2511.745 ;
        RECT 2637.030 2463.465 2637.330 2511.415 ;
        RECT 2637.015 2463.135 2637.345 2463.465 ;
        RECT 2639.775 2463.135 2640.105 2463.465 ;
        RECT 2639.790 2429.465 2640.090 2463.135 ;
        RECT 2639.775 2429.135 2640.105 2429.465 ;
        RECT 2638.855 2427.775 2639.185 2428.105 ;
        RECT 2638.870 2414.505 2639.170 2427.775 ;
        RECT 2638.855 2414.175 2639.185 2414.505 ;
        RECT 2640.695 2414.175 2641.025 2414.505 ;
        RECT 2640.710 2366.905 2641.010 2414.175 ;
        RECT 2637.935 2366.575 2638.265 2366.905 ;
        RECT 2640.695 2366.575 2641.025 2366.905 ;
        RECT 2637.950 2331.545 2638.250 2366.575 ;
        RECT 2636.095 2331.215 2636.425 2331.545 ;
        RECT 2637.935 2331.215 2638.265 2331.545 ;
        RECT 2636.110 2283.945 2636.410 2331.215 ;
        RECT 2636.095 2283.615 2636.425 2283.945 ;
        RECT 2638.855 2283.615 2639.185 2283.945 ;
        RECT 2638.870 2269.650 2639.170 2283.615 ;
        RECT 2637.950 2269.350 2639.170 2269.650 ;
        RECT 2637.950 2222.065 2638.250 2269.350 ;
        RECT 2636.095 2221.735 2636.425 2222.065 ;
        RECT 2637.935 2221.735 2638.265 2222.065 ;
        RECT 2636.110 2187.385 2636.410 2221.735 ;
        RECT 2636.095 2187.055 2636.425 2187.385 ;
        RECT 2639.775 2187.055 2640.105 2187.385 ;
        RECT 2639.790 2139.785 2640.090 2187.055 ;
        RECT 2639.775 2139.455 2640.105 2139.785 ;
        RECT 2638.855 2138.095 2639.185 2138.425 ;
        RECT 2638.870 2124.825 2639.170 2138.095 ;
        RECT 2638.855 2124.495 2639.185 2124.825 ;
        RECT 2637.015 2123.815 2637.345 2124.145 ;
        RECT 2637.030 2077.225 2637.330 2123.815 ;
        RECT 2637.015 2076.895 2637.345 2077.225 ;
        RECT 2639.775 2076.895 2640.105 2077.225 ;
        RECT 2639.790 2043.225 2640.090 2076.895 ;
        RECT 2639.775 2042.895 2640.105 2043.225 ;
        RECT 2638.855 2041.535 2639.185 2041.865 ;
        RECT 2638.870 2028.265 2639.170 2041.535 ;
        RECT 2636.095 2027.935 2636.425 2028.265 ;
        RECT 2638.855 2027.935 2639.185 2028.265 ;
        RECT 2636.110 1980.665 2636.410 2027.935 ;
        RECT 2636.095 1980.335 2636.425 1980.665 ;
        RECT 2637.935 1980.335 2638.265 1980.665 ;
        RECT 2637.950 1946.665 2638.250 1980.335 ;
        RECT 2637.935 1946.335 2638.265 1946.665 ;
        RECT 2637.015 1944.975 2637.345 1945.305 ;
        RECT 2637.030 1931.705 2637.330 1944.975 ;
        RECT 2637.015 1931.375 2637.345 1931.705 ;
        RECT 2639.775 1930.695 2640.105 1931.025 ;
        RECT 2639.790 1884.105 2640.090 1930.695 ;
        RECT 2637.935 1883.775 2638.265 1884.105 ;
        RECT 2639.775 1883.775 2640.105 1884.105 ;
        RECT 2637.950 1850.105 2638.250 1883.775 ;
        RECT 2637.935 1849.775 2638.265 1850.105 ;
        RECT 2638.855 1848.415 2639.185 1848.745 ;
        RECT 2638.870 1835.145 2639.170 1848.415 ;
        RECT 2638.855 1834.815 2639.185 1835.145 ;
        RECT 2641.615 1834.135 2641.945 1834.465 ;
        RECT 2641.630 1787.545 2641.930 1834.135 ;
        RECT 2639.775 1787.215 2640.105 1787.545 ;
        RECT 2641.615 1787.215 2641.945 1787.545 ;
        RECT 2639.790 1753.545 2640.090 1787.215 ;
        RECT 2639.775 1753.215 2640.105 1753.545 ;
        RECT 2638.855 1751.855 2639.185 1752.185 ;
        RECT 2638.870 1738.585 2639.170 1751.855 ;
        RECT 2638.855 1738.255 2639.185 1738.585 ;
        RECT 2641.615 1738.255 2641.945 1738.585 ;
        RECT 2641.630 1701.865 2641.930 1738.255 ;
        RECT 2637.935 1701.535 2638.265 1701.865 ;
        RECT 2641.615 1701.535 2641.945 1701.865 ;
        RECT 2637.950 1683.505 2638.250 1701.535 ;
        RECT 2637.935 1683.175 2638.265 1683.505 ;
        RECT 2637.015 1594.095 2637.345 1594.425 ;
        RECT 2637.030 1560.425 2637.330 1594.095 ;
        RECT 2637.015 1560.095 2637.345 1560.425 ;
        RECT 2637.935 1558.735 2638.265 1559.065 ;
        RECT 2637.950 1545.465 2638.250 1558.735 ;
        RECT 2637.935 1545.135 2638.265 1545.465 ;
        RECT 2637.015 1510.455 2637.345 1510.785 ;
        RECT 2637.030 1463.850 2637.330 1510.455 ;
        RECT 2637.030 1463.550 2638.250 1463.850 ;
        RECT 2637.950 1448.905 2638.250 1463.550 ;
        RECT 2637.935 1448.575 2638.265 1448.905 ;
        RECT 2637.015 1400.975 2637.345 1401.305 ;
        RECT 2637.030 1367.305 2637.330 1400.975 ;
        RECT 2637.015 1366.975 2637.345 1367.305 ;
        RECT 2637.935 1364.935 2638.265 1365.265 ;
        RECT 2637.950 1352.345 2638.250 1364.935 ;
        RECT 2637.935 1352.015 2638.265 1352.345 ;
        RECT 2637.015 1304.415 2637.345 1304.745 ;
        RECT 2637.030 1270.065 2637.330 1304.415 ;
        RECT 2637.015 1269.735 2637.345 1270.065 ;
        RECT 2637.935 1268.375 2638.265 1268.705 ;
        RECT 2637.950 1255.785 2638.250 1268.375 ;
        RECT 2637.935 1255.455 2638.265 1255.785 ;
        RECT 2637.015 1207.855 2637.345 1208.185 ;
        RECT 2637.030 1173.505 2637.330 1207.855 ;
        RECT 2637.015 1173.175 2637.345 1173.505 ;
        RECT 2637.935 1171.815 2638.265 1172.145 ;
        RECT 2637.950 1159.225 2638.250 1171.815 ;
        RECT 2637.935 1158.895 2638.265 1159.225 ;
        RECT 2638.855 1111.295 2639.185 1111.625 ;
        RECT 2638.870 1077.625 2639.170 1111.295 ;
        RECT 2638.855 1077.295 2639.185 1077.625 ;
        RECT 2637.935 1075.935 2638.265 1076.265 ;
        RECT 2637.950 1062.665 2638.250 1075.935 ;
        RECT 2637.935 1062.335 2638.265 1062.665 ;
        RECT 2637.015 1014.735 2637.345 1015.065 ;
        RECT 2637.030 980.385 2637.330 1014.735 ;
        RECT 2637.015 980.055 2637.345 980.385 ;
        RECT 2637.935 978.695 2638.265 979.025 ;
        RECT 2637.950 966.105 2638.250 978.695 ;
        RECT 2637.935 965.775 2638.265 966.105 ;
        RECT 2637.015 918.175 2637.345 918.505 ;
        RECT 2637.030 883.825 2637.330 918.175 ;
        RECT 2637.015 883.495 2637.345 883.825 ;
        RECT 2636.095 882.135 2636.425 882.465 ;
        RECT 2636.110 869.545 2636.410 882.135 ;
        RECT 2636.095 869.215 2636.425 869.545 ;
        RECT 2637.015 820.935 2637.345 821.265 ;
        RECT 2637.030 787.265 2637.330 820.935 ;
        RECT 2637.015 786.935 2637.345 787.265 ;
        RECT 2636.095 785.575 2636.425 785.905 ;
        RECT 2636.110 772.305 2636.410 785.575 ;
        RECT 2636.095 771.975 2636.425 772.305 ;
        RECT 2637.015 724.375 2637.345 724.705 ;
        RECT 2637.030 700.225 2637.330 724.375 ;
        RECT 2637.015 699.895 2637.345 700.225 ;
        RECT 2638.855 699.895 2639.185 700.225 ;
        RECT 2638.870 675.745 2639.170 699.895 ;
        RECT 2638.855 675.415 2639.185 675.745 ;
        RECT 2637.015 627.815 2637.345 628.145 ;
        RECT 2637.030 594.145 2637.330 627.815 ;
        RECT 2637.015 593.815 2637.345 594.145 ;
        RECT 2637.935 592.455 2638.265 592.785 ;
        RECT 2637.950 545.850 2638.250 592.455 ;
        RECT 2636.110 545.550 2638.250 545.850 ;
        RECT 2636.110 545.185 2636.410 545.550 ;
        RECT 2636.095 544.855 2636.425 545.185 ;
        RECT 2638.855 544.855 2639.185 545.185 ;
        RECT 2638.870 497.585 2639.170 544.855 ;
        RECT 2638.855 497.255 2639.185 497.585 ;
        RECT 2637.935 495.895 2638.265 496.225 ;
        RECT 2637.950 482.625 2638.250 495.895 ;
        RECT 2637.935 482.295 2638.265 482.625 ;
        RECT 2637.015 434.695 2637.345 435.025 ;
        RECT 2637.030 401.025 2637.330 434.695 ;
        RECT 2637.015 400.695 2637.345 401.025 ;
        RECT 2636.095 399.335 2636.425 399.665 ;
        RECT 2636.110 352.745 2636.410 399.335 ;
        RECT 2636.095 352.415 2636.425 352.745 ;
        RECT 2637.935 351.055 2638.265 351.385 ;
        RECT 2637.950 338.450 2638.250 351.055 ;
        RECT 2637.950 338.150 2639.170 338.450 ;
        RECT 2638.870 313.985 2639.170 338.150 ;
        RECT 2636.095 313.655 2636.425 313.985 ;
        RECT 2638.855 313.655 2639.185 313.985 ;
        RECT 2636.110 289.505 2636.410 313.655 ;
        RECT 2636.095 289.175 2636.425 289.505 ;
        RECT 2637.015 241.575 2637.345 241.905 ;
        RECT 2637.030 207.905 2637.330 241.575 ;
        RECT 2637.015 207.575 2637.345 207.905 ;
        RECT 2637.935 206.215 2638.265 206.545 ;
        RECT 2637.950 192.945 2638.250 206.215 ;
        RECT 2637.935 192.615 2638.265 192.945 ;
        RECT 2637.015 145.015 2637.345 145.345 ;
        RECT 2637.030 111.345 2637.330 145.015 ;
        RECT 2637.015 111.015 2637.345 111.345 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1193.770 851.600 1194.090 851.660 ;
        RECT 1241.610 851.600 1241.930 851.660 ;
        RECT 1193.770 851.460 1241.930 851.600 ;
        RECT 1193.770 851.400 1194.090 851.460 ;
        RECT 1241.610 851.400 1241.930 851.460 ;
        RECT 1448.150 849.900 1448.470 849.960 ;
        RECT 1464.710 849.900 1465.030 849.960 ;
        RECT 1448.150 849.760 1465.030 849.900 ;
        RECT 1448.150 849.700 1448.470 849.760 ;
        RECT 1464.710 849.700 1465.030 849.760 ;
        RECT 1338.670 849.560 1338.990 849.620 ;
        RECT 1393.410 849.560 1393.730 849.620 ;
        RECT 1338.670 849.420 1393.730 849.560 ;
        RECT 1338.670 849.360 1338.990 849.420 ;
        RECT 1393.410 849.360 1393.730 849.420 ;
        RECT 2379.650 849.560 2379.970 849.620 ;
        RECT 2390.690 849.560 2391.010 849.620 ;
        RECT 2379.650 849.420 2391.010 849.560 ;
        RECT 2379.650 849.360 2379.970 849.420 ;
        RECT 2390.690 849.360 2391.010 849.420 ;
        RECT 1630.310 849.220 1630.630 849.280 ;
        RECT 1656.530 849.220 1656.850 849.280 ;
        RECT 1630.310 849.080 1656.850 849.220 ;
        RECT 1630.310 849.020 1630.630 849.080 ;
        RECT 1656.530 849.020 1656.850 849.080 ;
        RECT 2125.270 849.220 2125.590 849.280 ;
        RECT 2172.650 849.220 2172.970 849.280 ;
        RECT 2125.270 849.080 2172.970 849.220 ;
        RECT 2125.270 849.020 2125.590 849.080 ;
        RECT 2172.650 849.020 2172.970 849.080 ;
      LAYER via ;
        RECT 1193.800 851.400 1194.060 851.660 ;
        RECT 1241.640 851.400 1241.900 851.660 ;
        RECT 1448.180 849.700 1448.440 849.960 ;
        RECT 1464.740 849.700 1465.000 849.960 ;
        RECT 1338.700 849.360 1338.960 849.620 ;
        RECT 1393.440 849.360 1393.700 849.620 ;
        RECT 2379.680 849.360 2379.940 849.620 ;
        RECT 2390.720 849.360 2390.980 849.620 ;
        RECT 1630.340 849.020 1630.600 849.280 ;
        RECT 1656.560 849.020 1656.820 849.280 ;
        RECT 2125.300 849.020 2125.560 849.280 ;
        RECT 2172.680 849.020 2172.940 849.280 ;
      LAYER met2 ;
        RECT 1299.590 3214.515 1299.870 3214.885 ;
        RECT 1299.660 3200.000 1299.800 3214.515 ;
        RECT 1299.520 3197.600 1299.800 3200.000 ;
        RECT 2801.030 852.195 2801.310 852.565 ;
        RECT 1193.790 851.515 1194.070 851.885 ;
        RECT 1193.800 851.370 1194.060 851.515 ;
        RECT 1241.640 851.370 1241.900 851.690 ;
        RECT 1296.830 851.515 1297.110 851.885 ;
        RECT 1931.630 851.515 1931.910 851.885 ;
        RECT 2608.290 851.515 2608.570 851.885 ;
        RECT 1241.700 850.525 1241.840 851.370 ;
        RECT 1241.630 850.155 1241.910 850.525 ;
        RECT 1296.900 849.845 1297.040 851.515 ;
        RECT 1779.830 850.835 1780.110 851.205 ;
        RECT 1835.030 850.835 1835.310 851.205 ;
        RECT 1464.730 850.155 1465.010 850.525 ;
        RECT 1490.950 850.155 1491.230 850.525 ;
        RECT 1587.550 850.155 1587.830 850.525 ;
        RECT 1656.550 850.155 1656.830 850.525 ;
        RECT 1690.130 850.155 1690.410 850.525 ;
        RECT 1464.800 849.990 1464.940 850.155 ;
        RECT 1448.180 849.845 1448.440 849.990 ;
        RECT 1296.830 849.475 1297.110 849.845 ;
        RECT 1338.690 849.475 1338.970 849.845 ;
        RECT 1338.700 849.330 1338.960 849.475 ;
        RECT 1393.440 849.330 1393.700 849.650 ;
        RECT 1417.350 849.475 1417.630 849.845 ;
        RECT 1448.170 849.475 1448.450 849.845 ;
        RECT 1464.740 849.670 1465.000 849.990 ;
        RECT 1491.020 849.845 1491.160 850.155 ;
        RECT 1490.950 849.475 1491.230 849.845 ;
        RECT 1393.500 849.165 1393.640 849.330 ;
        RECT 1393.430 848.795 1393.710 849.165 ;
        RECT 1417.420 847.805 1417.560 849.475 ;
        RECT 1587.620 849.165 1587.760 850.155 ;
        RECT 1656.620 849.310 1656.760 850.155 ;
        RECT 1630.340 849.165 1630.600 849.310 ;
        RECT 1587.550 848.795 1587.830 849.165 ;
        RECT 1630.330 848.795 1630.610 849.165 ;
        RECT 1656.560 848.990 1656.820 849.310 ;
        RECT 1690.200 848.485 1690.340 850.155 ;
        RECT 1690.130 848.115 1690.410 848.485 ;
        RECT 1779.900 847.805 1780.040 850.835 ;
        RECT 1835.100 849.165 1835.240 850.835 ;
        RECT 1859.410 850.155 1859.690 850.525 ;
        RECT 1859.480 849.165 1859.620 850.155 ;
        RECT 1931.700 849.845 1931.840 851.515 ;
        RECT 2172.670 850.155 2172.950 850.525 ;
        RECT 1931.630 849.475 1931.910 849.845 ;
        RECT 2090.330 849.475 2090.610 849.845 ;
        RECT 1835.030 848.795 1835.310 849.165 ;
        RECT 1859.410 848.795 1859.690 849.165 ;
        RECT 2090.400 847.805 2090.540 849.475 ;
        RECT 2172.740 849.310 2172.880 850.155 ;
        RECT 2379.670 849.475 2379.950 849.845 ;
        RECT 2390.710 849.475 2390.990 849.845 ;
        RECT 2379.680 849.330 2379.940 849.475 ;
        RECT 2390.720 849.330 2390.980 849.475 ;
        RECT 2125.300 849.165 2125.560 849.310 ;
        RECT 2125.290 848.795 2125.570 849.165 ;
        RECT 2172.680 848.990 2172.940 849.310 ;
        RECT 2608.360 849.165 2608.500 851.515 ;
        RECT 2704.430 850.835 2704.710 851.205 ;
        RECT 2704.500 849.845 2704.640 850.835 ;
        RECT 2801.100 850.525 2801.240 852.195 ;
        RECT 2801.030 850.155 2801.310 850.525 ;
        RECT 2704.430 849.475 2704.710 849.845 ;
        RECT 2863.130 849.475 2863.410 849.845 ;
        RECT 2608.290 848.795 2608.570 849.165 ;
        RECT 2863.200 849.050 2863.340 849.475 ;
        RECT 2863.590 849.050 2863.870 849.165 ;
        RECT 2863.200 848.910 2863.870 849.050 ;
        RECT 2863.590 848.795 2863.870 848.910 ;
        RECT 1417.350 847.435 1417.630 847.805 ;
        RECT 1779.830 847.435 1780.110 847.805 ;
        RECT 2090.330 847.435 2090.610 847.805 ;
      LAYER via2 ;
        RECT 1299.590 3214.560 1299.870 3214.840 ;
        RECT 2801.030 852.240 2801.310 852.520 ;
        RECT 1193.790 851.560 1194.070 851.840 ;
        RECT 1296.830 851.560 1297.110 851.840 ;
        RECT 1931.630 851.560 1931.910 851.840 ;
        RECT 2608.290 851.560 2608.570 851.840 ;
        RECT 1241.630 850.200 1241.910 850.480 ;
        RECT 1779.830 850.880 1780.110 851.160 ;
        RECT 1835.030 850.880 1835.310 851.160 ;
        RECT 1464.730 850.200 1465.010 850.480 ;
        RECT 1490.950 850.200 1491.230 850.480 ;
        RECT 1587.550 850.200 1587.830 850.480 ;
        RECT 1656.550 850.200 1656.830 850.480 ;
        RECT 1690.130 850.200 1690.410 850.480 ;
        RECT 1296.830 849.520 1297.110 849.800 ;
        RECT 1338.690 849.520 1338.970 849.800 ;
        RECT 1417.350 849.520 1417.630 849.800 ;
        RECT 1448.170 849.520 1448.450 849.800 ;
        RECT 1490.950 849.520 1491.230 849.800 ;
        RECT 1393.430 848.840 1393.710 849.120 ;
        RECT 1587.550 848.840 1587.830 849.120 ;
        RECT 1630.330 848.840 1630.610 849.120 ;
        RECT 1690.130 848.160 1690.410 848.440 ;
        RECT 1859.410 850.200 1859.690 850.480 ;
        RECT 2172.670 850.200 2172.950 850.480 ;
        RECT 1931.630 849.520 1931.910 849.800 ;
        RECT 2090.330 849.520 2090.610 849.800 ;
        RECT 1835.030 848.840 1835.310 849.120 ;
        RECT 1859.410 848.840 1859.690 849.120 ;
        RECT 2379.670 849.520 2379.950 849.800 ;
        RECT 2390.710 849.520 2390.990 849.800 ;
        RECT 2125.290 848.840 2125.570 849.120 ;
        RECT 2704.430 850.880 2704.710 851.160 ;
        RECT 2801.030 850.200 2801.310 850.480 ;
        RECT 2704.430 849.520 2704.710 849.800 ;
        RECT 2863.130 849.520 2863.410 849.800 ;
        RECT 2608.290 848.840 2608.570 849.120 ;
        RECT 2863.590 848.840 2863.870 849.120 ;
        RECT 1417.350 847.480 1417.630 847.760 ;
        RECT 1779.830 847.480 1780.110 847.760 ;
        RECT 2090.330 847.480 2090.610 847.760 ;
      LAYER met3 ;
        RECT 1168.670 3214.850 1169.050 3214.860 ;
        RECT 1299.565 3214.850 1299.895 3214.865 ;
        RECT 1168.670 3214.550 1299.895 3214.850 ;
        RECT 1168.670 3214.540 1169.050 3214.550 ;
        RECT 1299.565 3214.535 1299.895 3214.550 ;
        RECT 2752.910 852.530 2753.290 852.540 ;
        RECT 2801.005 852.530 2801.335 852.545 ;
        RECT 2752.910 852.230 2801.335 852.530 ;
        RECT 2752.910 852.220 2753.290 852.230 ;
        RECT 2801.005 852.215 2801.335 852.230 ;
        RECT 1168.670 851.850 1169.050 851.860 ;
        RECT 1193.765 851.850 1194.095 851.865 ;
        RECT 1168.670 851.550 1194.095 851.850 ;
        RECT 1168.670 851.540 1169.050 851.550 ;
        RECT 1193.765 851.535 1194.095 851.550 ;
        RECT 1243.190 851.850 1243.570 851.860 ;
        RECT 1296.805 851.850 1297.135 851.865 ;
        RECT 1243.190 851.550 1297.135 851.850 ;
        RECT 1243.190 851.540 1243.570 851.550 ;
        RECT 1296.805 851.535 1297.135 851.550 ;
        RECT 1883.510 851.850 1883.890 851.860 ;
        RECT 1931.605 851.850 1931.935 851.865 ;
        RECT 1883.510 851.550 1931.935 851.850 ;
        RECT 1883.510 851.540 1883.890 851.550 ;
        RECT 1931.605 851.535 1931.935 851.550 ;
        RECT 2608.265 851.850 2608.595 851.865 ;
        RECT 2608.265 851.550 2656.650 851.850 ;
        RECT 2608.265 851.535 2608.595 851.550 ;
        RECT 1779.805 851.170 1780.135 851.185 ;
        RECT 1835.005 851.170 1835.335 851.185 ;
        RECT 2656.350 851.170 2656.650 851.550 ;
        RECT 2704.405 851.170 2704.735 851.185 ;
        RECT 2752.910 851.170 2753.290 851.180 ;
        RECT 1558.790 850.870 1586.690 851.170 ;
        RECT 1241.605 850.490 1241.935 850.505 ;
        RECT 1242.270 850.490 1242.650 850.500 ;
        RECT 1241.605 850.190 1242.650 850.490 ;
        RECT 1241.605 850.175 1241.935 850.190 ;
        RECT 1242.270 850.180 1242.650 850.190 ;
        RECT 1464.705 850.490 1465.035 850.505 ;
        RECT 1490.925 850.490 1491.255 850.505 ;
        RECT 1464.705 850.190 1491.255 850.490 ;
        RECT 1464.705 850.175 1465.035 850.190 ;
        RECT 1490.925 850.175 1491.255 850.190 ;
        RECT 1296.805 849.810 1297.135 849.825 ;
        RECT 1338.665 849.810 1338.995 849.825 ;
        RECT 1296.805 849.510 1338.995 849.810 ;
        RECT 1296.805 849.495 1297.135 849.510 ;
        RECT 1338.665 849.495 1338.995 849.510 ;
        RECT 1417.325 849.810 1417.655 849.825 ;
        RECT 1448.145 849.810 1448.475 849.825 ;
        RECT 1417.325 849.510 1448.475 849.810 ;
        RECT 1417.325 849.495 1417.655 849.510 ;
        RECT 1448.145 849.495 1448.475 849.510 ;
        RECT 1490.925 849.810 1491.255 849.825 ;
        RECT 1558.790 849.810 1559.090 850.870 ;
        RECT 1586.390 850.490 1586.690 850.870 ;
        RECT 1779.805 850.870 1835.335 851.170 ;
        RECT 1779.805 850.855 1780.135 850.870 ;
        RECT 1835.005 850.855 1835.335 850.870 ;
        RECT 2282.830 850.870 2318.090 851.170 ;
        RECT 1587.525 850.490 1587.855 850.505 ;
        RECT 1586.390 850.190 1587.855 850.490 ;
        RECT 1587.525 850.175 1587.855 850.190 ;
        RECT 1656.525 850.490 1656.855 850.505 ;
        RECT 1690.105 850.490 1690.435 850.505 ;
        RECT 1656.525 850.190 1690.435 850.490 ;
        RECT 1656.525 850.175 1656.855 850.190 ;
        RECT 1690.105 850.175 1690.435 850.190 ;
        RECT 1859.385 850.490 1859.715 850.505 ;
        RECT 1883.510 850.490 1883.890 850.500 ;
        RECT 2172.645 850.490 2172.975 850.505 ;
        RECT 1859.385 850.190 1883.890 850.490 ;
        RECT 1859.385 850.175 1859.715 850.190 ;
        RECT 1883.510 850.180 1883.890 850.190 ;
        RECT 1946.110 850.190 1994.250 850.490 ;
        RECT 1490.925 849.510 1559.090 849.810 ;
        RECT 1931.605 849.810 1931.935 849.825 ;
        RECT 1946.110 849.810 1946.410 850.190 ;
        RECT 1931.605 849.510 1946.410 849.810 ;
        RECT 1490.925 849.495 1491.255 849.510 ;
        RECT 1931.605 849.495 1931.935 849.510 ;
        RECT 1393.405 849.130 1393.735 849.145 ;
        RECT 1587.525 849.130 1587.855 849.145 ;
        RECT 1630.305 849.130 1630.635 849.145 ;
        RECT 1835.005 849.130 1835.335 849.145 ;
        RECT 1859.385 849.130 1859.715 849.145 ;
        RECT 1393.405 848.830 1394.410 849.130 ;
        RECT 1393.405 848.815 1393.735 848.830 ;
        RECT 1394.110 847.770 1394.410 848.830 ;
        RECT 1587.525 848.830 1630.635 849.130 ;
        RECT 1587.525 848.815 1587.855 848.830 ;
        RECT 1630.305 848.815 1630.635 848.830 ;
        RECT 1691.270 848.830 1732.050 849.130 ;
        RECT 1690.105 848.450 1690.435 848.465 ;
        RECT 1691.270 848.450 1691.570 848.830 ;
        RECT 1690.105 848.150 1691.570 848.450 ;
        RECT 1690.105 848.135 1690.435 848.150 ;
        RECT 1417.325 847.770 1417.655 847.785 ;
        RECT 1394.110 847.470 1417.655 847.770 ;
        RECT 1731.750 847.770 1732.050 848.830 ;
        RECT 1835.005 848.830 1859.715 849.130 ;
        RECT 1993.950 849.130 1994.250 850.190 ;
        RECT 2172.645 850.190 2187.450 850.490 ;
        RECT 2172.645 850.175 2172.975 850.190 ;
        RECT 2090.305 849.810 2090.635 849.825 ;
        RECT 2042.710 849.510 2090.635 849.810 ;
        RECT 2042.710 849.130 2043.010 849.510 ;
        RECT 2090.305 849.495 2090.635 849.510 ;
        RECT 2125.265 849.130 2125.595 849.145 ;
        RECT 1993.950 848.830 2043.010 849.130 ;
        RECT 2124.590 848.830 2125.595 849.130 ;
        RECT 2187.150 849.130 2187.450 850.190 ;
        RECT 2282.830 849.810 2283.130 850.870 ;
        RECT 2235.910 849.510 2283.130 849.810 ;
        RECT 2235.910 849.130 2236.210 849.510 ;
        RECT 2187.150 848.830 2236.210 849.130 ;
        RECT 2317.790 849.130 2318.090 850.870 ;
        RECT 2476.030 850.870 2511.290 851.170 ;
        RECT 2656.350 850.870 2704.735 851.170 ;
        RECT 2379.645 849.810 2379.975 849.825 ;
        RECT 2332.510 849.510 2379.975 849.810 ;
        RECT 2332.510 849.130 2332.810 849.510 ;
        RECT 2379.645 849.495 2379.975 849.510 ;
        RECT 2390.685 849.810 2391.015 849.825 ;
        RECT 2476.030 849.810 2476.330 850.870 ;
        RECT 2390.685 849.510 2414.690 849.810 ;
        RECT 2390.685 849.495 2391.015 849.510 ;
        RECT 2317.790 848.830 2332.810 849.130 ;
        RECT 2414.390 849.130 2414.690 849.510 ;
        RECT 2429.110 849.510 2476.330 849.810 ;
        RECT 2429.110 849.130 2429.410 849.510 ;
        RECT 2414.390 848.830 2429.410 849.130 ;
        RECT 2510.990 849.130 2511.290 850.870 ;
        RECT 2704.405 850.855 2704.735 850.870 ;
        RECT 2718.910 850.870 2753.290 851.170 ;
        RECT 2704.405 849.810 2704.735 849.825 ;
        RECT 2718.910 849.810 2719.210 850.870 ;
        RECT 2752.910 850.860 2753.290 850.870 ;
        RECT 2801.005 850.490 2801.335 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2801.005 850.190 2815.810 850.490 ;
        RECT 2801.005 850.175 2801.335 850.190 ;
        RECT 2525.710 849.510 2607.890 849.810 ;
        RECT 2525.710 849.130 2526.010 849.510 ;
        RECT 2510.990 848.830 2526.010 849.130 ;
        RECT 2607.590 849.130 2607.890 849.510 ;
        RECT 2704.405 849.510 2719.210 849.810 ;
        RECT 2704.405 849.495 2704.735 849.510 ;
        RECT 2608.265 849.130 2608.595 849.145 ;
        RECT 2607.590 848.830 2608.595 849.130 ;
        RECT 2815.510 849.130 2815.810 850.190 ;
        RECT 2916.710 850.190 2924.800 850.490 ;
        RECT 2863.105 849.810 2863.435 849.825 ;
        RECT 2916.710 849.810 2917.010 850.190 ;
        RECT 2849.550 849.510 2863.435 849.810 ;
        RECT 2849.550 849.130 2849.850 849.510 ;
        RECT 2863.105 849.495 2863.435 849.510 ;
        RECT 2884.510 849.510 2917.010 849.810 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT 2815.510 848.830 2849.850 849.130 ;
        RECT 2863.565 849.130 2863.895 849.145 ;
        RECT 2884.510 849.130 2884.810 849.510 ;
        RECT 2863.565 848.830 2884.810 849.130 ;
        RECT 1835.005 848.815 1835.335 848.830 ;
        RECT 1859.385 848.815 1859.715 848.830 ;
        RECT 1779.805 847.770 1780.135 847.785 ;
        RECT 1731.750 847.470 1780.135 847.770 ;
        RECT 1417.325 847.455 1417.655 847.470 ;
        RECT 1779.805 847.455 1780.135 847.470 ;
        RECT 2090.305 847.770 2090.635 847.785 ;
        RECT 2124.590 847.770 2124.890 848.830 ;
        RECT 2125.265 848.815 2125.595 848.830 ;
        RECT 2608.265 848.815 2608.595 848.830 ;
        RECT 2863.565 848.815 2863.895 848.830 ;
        RECT 2090.305 847.470 2124.890 847.770 ;
        RECT 2090.305 847.455 2090.635 847.470 ;
      LAYER via3 ;
        RECT 1168.700 3214.540 1169.020 3214.860 ;
        RECT 2752.940 852.220 2753.260 852.540 ;
        RECT 1168.700 851.540 1169.020 851.860 ;
        RECT 1243.220 851.540 1243.540 851.860 ;
        RECT 1883.540 851.540 1883.860 851.860 ;
        RECT 1242.300 850.180 1242.620 850.500 ;
        RECT 1883.540 850.180 1883.860 850.500 ;
        RECT 2752.940 850.860 2753.260 851.180 ;
      LAYER met4 ;
        RECT 1168.695 3214.535 1169.025 3214.865 ;
        RECT 1168.710 851.865 1169.010 3214.535 ;
        RECT 2752.935 852.215 2753.265 852.545 ;
        RECT 1168.695 851.535 1169.025 851.865 ;
        RECT 1243.215 851.535 1243.545 851.865 ;
        RECT 1883.535 851.535 1883.865 851.865 ;
        RECT 1242.295 850.490 1242.625 850.505 ;
        RECT 1243.230 850.490 1243.530 851.535 ;
        RECT 1883.550 850.505 1883.850 851.535 ;
        RECT 2752.950 851.185 2753.250 852.215 ;
        RECT 2752.935 850.855 2753.265 851.185 ;
        RECT 1242.295 850.190 1243.530 850.490 ;
        RECT 1242.295 850.175 1242.625 850.190 ;
        RECT 1883.535 850.175 1883.865 850.505 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.110 3353.660 1345.430 3353.720 ;
        RECT 2887.490 3353.660 2887.810 3353.720 ;
        RECT 1345.110 3353.520 2887.810 3353.660 ;
        RECT 1345.110 3353.460 1345.430 3353.520 ;
        RECT 2887.490 3353.460 2887.810 3353.520 ;
        RECT 1339.130 3213.240 1339.450 3213.300 ;
        RECT 1345.110 3213.240 1345.430 3213.300 ;
        RECT 1339.130 3213.100 1345.430 3213.240 ;
        RECT 1339.130 3213.040 1339.450 3213.100 ;
        RECT 1345.110 3213.040 1345.430 3213.100 ;
        RECT 2887.490 1089.940 2887.810 1090.000 ;
        RECT 2898.070 1089.940 2898.390 1090.000 ;
        RECT 2887.490 1089.800 2898.390 1089.940 ;
        RECT 2887.490 1089.740 2887.810 1089.800 ;
        RECT 2898.070 1089.740 2898.390 1089.800 ;
      LAYER via ;
        RECT 1345.140 3353.460 1345.400 3353.720 ;
        RECT 2887.520 3353.460 2887.780 3353.720 ;
        RECT 1339.160 3213.040 1339.420 3213.300 ;
        RECT 1345.140 3213.040 1345.400 3213.300 ;
        RECT 2887.520 1089.740 2887.780 1090.000 ;
        RECT 2898.100 1089.740 2898.360 1090.000 ;
      LAYER met2 ;
        RECT 1345.140 3353.430 1345.400 3353.750 ;
        RECT 2887.520 3353.430 2887.780 3353.750 ;
        RECT 1345.200 3213.330 1345.340 3353.430 ;
        RECT 1339.160 3213.010 1339.420 3213.330 ;
        RECT 1345.140 3213.010 1345.400 3213.330 ;
        RECT 1339.220 3200.000 1339.360 3213.010 ;
        RECT 1339.080 3197.600 1339.360 3200.000 ;
        RECT 2887.580 1090.030 2887.720 3353.430 ;
        RECT 2887.520 1089.710 2887.780 1090.030 ;
        RECT 2898.100 1089.710 2898.360 1090.030 ;
        RECT 2898.160 1085.125 2898.300 1089.710 ;
        RECT 2898.090 1084.755 2898.370 1085.125 ;
      LAYER via2 ;
        RECT 2898.090 1084.800 2898.370 1085.080 ;
      LAYER met3 ;
        RECT 2898.065 1085.090 2898.395 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2898.065 1084.790 2924.800 1085.090 ;
        RECT 2898.065 1084.775 2898.395 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1378.690 3206.100 1379.010 3206.160 ;
        RECT 2653.810 3206.100 2654.130 3206.160 ;
        RECT 1378.690 3205.960 2654.130 3206.100 ;
        RECT 1378.690 3205.900 1379.010 3205.960 ;
        RECT 2653.810 3205.900 2654.130 3205.960 ;
        RECT 2653.810 1324.540 2654.130 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2653.810 1324.400 2901.150 1324.540 ;
        RECT 2653.810 1324.340 2654.130 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 1378.720 3205.900 1378.980 3206.160 ;
        RECT 2653.840 3205.900 2654.100 3206.160 ;
        RECT 2653.840 1324.340 2654.100 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 1378.720 3205.870 1378.980 3206.190 ;
        RECT 2653.840 3205.870 2654.100 3206.190 ;
        RECT 1378.780 3200.000 1378.920 3205.870 ;
        RECT 1378.640 3197.600 1378.920 3200.000 ;
        RECT 2653.900 1324.630 2654.040 3205.870 ;
        RECT 2653.840 1324.310 2654.100 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2138.700 3215.480 2139.300 3215.620 ;
        RECT 1418.250 3215.280 1418.570 3215.340 ;
        RECT 2138.700 3215.280 2138.840 3215.480 ;
        RECT 2139.160 3215.340 2139.300 3215.480 ;
        RECT 1418.250 3215.140 2138.840 3215.280 ;
        RECT 1418.250 3215.080 1418.570 3215.140 ;
        RECT 2139.070 3215.080 2139.390 3215.340 ;
        RECT 2139.070 3208.480 2139.390 3208.540 ;
        RECT 2901.750 3208.480 2902.070 3208.540 ;
        RECT 2139.070 3208.340 2902.070 3208.480 ;
        RECT 2139.070 3208.280 2139.390 3208.340 ;
        RECT 2901.750 3208.280 2902.070 3208.340 ;
      LAYER via ;
        RECT 1418.280 3215.080 1418.540 3215.340 ;
        RECT 2139.100 3215.080 2139.360 3215.340 ;
        RECT 2139.100 3208.280 2139.360 3208.540 ;
        RECT 2901.780 3208.280 2902.040 3208.540 ;
      LAYER met2 ;
        RECT 1418.280 3215.050 1418.540 3215.370 ;
        RECT 2139.100 3215.050 2139.360 3215.370 ;
        RECT 1418.340 3200.000 1418.480 3215.050 ;
        RECT 2139.160 3208.570 2139.300 3215.050 ;
        RECT 2139.100 3208.250 2139.360 3208.570 ;
        RECT 2901.780 3208.250 2902.040 3208.570 ;
        RECT 1418.200 3197.600 1418.480 3200.000 ;
        RECT 2901.840 3196.410 2901.980 3208.250 ;
        RECT 2900.920 3196.270 2901.980 3196.410 ;
        RECT 2900.920 1554.325 2901.060 3196.270 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1457.350 3205.080 1457.670 3205.140 ;
        RECT 2900.370 3205.080 2900.690 3205.140 ;
        RECT 1457.350 3204.940 2900.690 3205.080 ;
        RECT 1457.350 3204.880 1457.670 3204.940 ;
        RECT 2900.370 3204.880 2900.690 3204.940 ;
      LAYER via ;
        RECT 1457.380 3204.880 1457.640 3205.140 ;
        RECT 2900.400 3204.880 2900.660 3205.140 ;
      LAYER met2 ;
        RECT 1457.380 3204.850 1457.640 3205.170 ;
        RECT 2900.400 3204.850 2900.660 3205.170 ;
        RECT 1457.440 3200.000 1457.580 3204.850 ;
        RECT 1457.300 3197.600 1457.580 3200.000 ;
        RECT 2900.460 1789.605 2900.600 3204.850 ;
        RECT 2900.390 1789.235 2900.670 1789.605 ;
      LAYER via2 ;
        RECT 2900.390 1789.280 2900.670 1789.560 ;
      LAYER met3 ;
        RECT 2900.365 1789.570 2900.695 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.365 1789.270 2924.800 1789.570 ;
        RECT 2900.365 1789.255 2900.695 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1496.910 3206.780 1497.230 3206.840 ;
        RECT 2659.790 3206.780 2660.110 3206.840 ;
        RECT 1496.910 3206.640 2660.110 3206.780 ;
        RECT 1496.910 3206.580 1497.230 3206.640 ;
        RECT 2659.790 3206.580 2660.110 3206.640 ;
        RECT 2659.790 2028.340 2660.110 2028.400 ;
        RECT 2899.450 2028.340 2899.770 2028.400 ;
        RECT 2659.790 2028.200 2899.770 2028.340 ;
        RECT 2659.790 2028.140 2660.110 2028.200 ;
        RECT 2899.450 2028.140 2899.770 2028.200 ;
      LAYER via ;
        RECT 1496.940 3206.580 1497.200 3206.840 ;
        RECT 2659.820 3206.580 2660.080 3206.840 ;
        RECT 2659.820 2028.140 2660.080 2028.400 ;
        RECT 2899.480 2028.140 2899.740 2028.400 ;
      LAYER met2 ;
        RECT 1496.940 3206.550 1497.200 3206.870 ;
        RECT 2659.820 3206.550 2660.080 3206.870 ;
        RECT 1497.000 3200.000 1497.140 3206.550 ;
        RECT 1496.860 3197.600 1497.140 3200.000 ;
        RECT 2659.880 2028.430 2660.020 3206.550 ;
        RECT 2659.820 2028.110 2660.080 2028.430 ;
        RECT 2899.480 2028.110 2899.740 2028.430 ;
        RECT 2899.540 2024.205 2899.680 2028.110 ;
        RECT 2899.470 2023.835 2899.750 2024.205 ;
      LAYER via2 ;
        RECT 2899.470 2023.880 2899.750 2024.160 ;
      LAYER met3 ;
        RECT 2899.445 2024.170 2899.775 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2899.445 2023.870 2924.800 2024.170 ;
        RECT 2899.445 2023.855 2899.775 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1536.470 3214.940 1536.790 3215.000 ;
        RECT 2366.770 3214.940 2367.090 3215.000 ;
        RECT 1536.470 3214.800 2367.090 3214.940 ;
        RECT 1536.470 3214.740 1536.790 3214.800 ;
        RECT 2366.770 3214.740 2367.090 3214.800 ;
        RECT 2366.770 3204.400 2367.090 3204.460 ;
        RECT 2899.450 3204.400 2899.770 3204.460 ;
        RECT 2366.770 3204.260 2899.770 3204.400 ;
        RECT 2366.770 3204.200 2367.090 3204.260 ;
        RECT 2899.450 3204.200 2899.770 3204.260 ;
      LAYER via ;
        RECT 1536.500 3214.740 1536.760 3215.000 ;
        RECT 2366.800 3214.740 2367.060 3215.000 ;
        RECT 2366.800 3204.200 2367.060 3204.460 ;
        RECT 2899.480 3204.200 2899.740 3204.460 ;
      LAYER met2 ;
        RECT 1536.500 3214.710 1536.760 3215.030 ;
        RECT 2366.800 3214.710 2367.060 3215.030 ;
        RECT 1536.560 3200.000 1536.700 3214.710 ;
        RECT 2366.860 3204.490 2367.000 3214.710 ;
        RECT 2366.800 3204.170 2367.060 3204.490 ;
        RECT 2899.480 3204.170 2899.740 3204.490 ;
        RECT 1536.420 3197.600 1536.700 3200.000 ;
        RECT 2899.540 2258.805 2899.680 3204.170 ;
        RECT 2899.470 2258.435 2899.750 2258.805 ;
      LAYER via2 ;
        RECT 2899.470 2258.480 2899.750 2258.760 ;
      LAYER met3 ;
        RECT 2899.445 2258.770 2899.775 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2899.445 2258.470 2924.800 2258.770 ;
        RECT 2899.445 2258.455 2899.775 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1470.305 1580.065 1470.475 1669.655 ;
        RECT 1470.305 745.365 1470.475 793.475 ;
        RECT 1470.305 607.325 1470.475 696.915 ;
        RECT 1470.765 582.845 1470.935 606.815 ;
        RECT 1470.765 145.265 1470.935 193.035 ;
        RECT 1469.845 89.845 1470.015 137.955 ;
        RECT 1469.845 59.245 1470.015 62.475 ;
      LAYER mcon ;
        RECT 1470.305 1669.485 1470.475 1669.655 ;
        RECT 1470.305 793.305 1470.475 793.475 ;
        RECT 1470.305 696.745 1470.475 696.915 ;
        RECT 1470.765 606.645 1470.935 606.815 ;
        RECT 1470.765 192.865 1470.935 193.035 ;
        RECT 1469.845 137.785 1470.015 137.955 ;
        RECT 1469.845 62.305 1470.015 62.475 ;
      LAYER met1 ;
        RECT 1470.230 1669.640 1470.550 1669.700 ;
        RECT 1470.035 1669.500 1470.550 1669.640 ;
        RECT 1470.230 1669.440 1470.550 1669.500 ;
        RECT 1470.245 1580.220 1470.535 1580.265 ;
        RECT 1470.690 1580.220 1471.010 1580.280 ;
        RECT 1470.245 1580.080 1471.010 1580.220 ;
        RECT 1470.245 1580.035 1470.535 1580.080 ;
        RECT 1470.690 1580.020 1471.010 1580.080 ;
        RECT 1470.690 1559.620 1471.010 1559.880 ;
        RECT 1470.780 1559.200 1470.920 1559.620 ;
        RECT 1470.690 1558.940 1471.010 1559.200 ;
        RECT 1470.690 1365.820 1471.010 1366.080 ;
        RECT 1470.780 1365.400 1470.920 1365.820 ;
        RECT 1470.690 1365.140 1471.010 1365.400 ;
        RECT 1470.690 1269.260 1471.010 1269.520 ;
        RECT 1470.780 1268.840 1470.920 1269.260 ;
        RECT 1470.690 1268.580 1471.010 1268.840 ;
        RECT 1470.690 1172.700 1471.010 1172.960 ;
        RECT 1470.780 1172.280 1470.920 1172.700 ;
        RECT 1470.690 1172.020 1471.010 1172.280 ;
        RECT 1470.690 965.980 1471.010 966.240 ;
        RECT 1470.780 965.840 1470.920 965.980 ;
        RECT 1471.150 965.840 1471.470 965.900 ;
        RECT 1470.780 965.700 1471.470 965.840 ;
        RECT 1471.150 965.640 1471.470 965.700 ;
        RECT 1470.230 917.900 1470.550 917.960 ;
        RECT 1471.150 917.900 1471.470 917.960 ;
        RECT 1470.230 917.760 1471.470 917.900 ;
        RECT 1470.230 917.700 1470.550 917.760 ;
        RECT 1471.150 917.700 1471.470 917.760 ;
        RECT 1470.230 883.360 1470.550 883.620 ;
        RECT 1470.320 882.880 1470.460 883.360 ;
        RECT 1470.690 882.880 1471.010 882.940 ;
        RECT 1470.320 882.740 1471.010 882.880 ;
        RECT 1470.690 882.680 1471.010 882.740 ;
        RECT 1470.690 796.860 1471.010 796.920 ;
        RECT 1471.610 796.860 1471.930 796.920 ;
        RECT 1470.690 796.720 1471.930 796.860 ;
        RECT 1470.690 796.660 1471.010 796.720 ;
        RECT 1471.610 796.660 1471.930 796.720 ;
        RECT 1470.245 793.460 1470.535 793.505 ;
        RECT 1471.610 793.460 1471.930 793.520 ;
        RECT 1470.245 793.320 1471.930 793.460 ;
        RECT 1470.245 793.275 1470.535 793.320 ;
        RECT 1471.610 793.260 1471.930 793.320 ;
        RECT 1470.230 745.520 1470.550 745.580 ;
        RECT 1470.035 745.380 1470.550 745.520 ;
        RECT 1470.230 745.320 1470.550 745.380 ;
        RECT 1470.230 696.900 1470.550 696.960 ;
        RECT 1470.035 696.760 1470.550 696.900 ;
        RECT 1470.230 696.700 1470.550 696.760 ;
        RECT 1470.245 607.480 1470.535 607.525 ;
        RECT 1470.690 607.480 1471.010 607.540 ;
        RECT 1470.245 607.340 1471.010 607.480 ;
        RECT 1470.245 607.295 1470.535 607.340 ;
        RECT 1470.690 607.280 1471.010 607.340 ;
        RECT 1470.690 606.800 1471.010 606.860 ;
        RECT 1470.495 606.660 1471.010 606.800 ;
        RECT 1470.690 606.600 1471.010 606.660 ;
        RECT 1470.690 583.000 1471.010 583.060 ;
        RECT 1470.495 582.860 1471.010 583.000 ;
        RECT 1470.690 582.800 1471.010 582.860 ;
        RECT 1470.690 400.560 1471.010 400.820 ;
        RECT 1470.780 400.140 1470.920 400.560 ;
        RECT 1470.690 399.880 1471.010 400.140 ;
        RECT 1469.770 289.920 1470.090 289.980 ;
        RECT 1470.690 289.920 1471.010 289.980 ;
        RECT 1469.770 289.780 1471.010 289.920 ;
        RECT 1469.770 289.720 1470.090 289.780 ;
        RECT 1470.690 289.720 1471.010 289.780 ;
        RECT 1470.690 193.020 1471.010 193.080 ;
        RECT 1470.495 192.880 1471.010 193.020 ;
        RECT 1470.690 192.820 1471.010 192.880 ;
        RECT 1470.690 145.420 1471.010 145.480 ;
        RECT 1470.495 145.280 1471.010 145.420 ;
        RECT 1470.690 145.220 1471.010 145.280 ;
        RECT 1469.770 144.740 1470.090 144.800 ;
        RECT 1470.690 144.740 1471.010 144.800 ;
        RECT 1469.770 144.600 1471.010 144.740 ;
        RECT 1469.770 144.540 1470.090 144.600 ;
        RECT 1470.690 144.540 1471.010 144.600 ;
        RECT 1469.770 137.940 1470.090 138.000 ;
        RECT 1469.575 137.800 1470.090 137.940 ;
        RECT 1469.770 137.740 1470.090 137.800 ;
        RECT 1469.770 90.000 1470.090 90.060 ;
        RECT 1469.575 89.860 1470.090 90.000 ;
        RECT 1469.770 89.800 1470.090 89.860 ;
        RECT 1469.770 62.460 1470.090 62.520 ;
        RECT 1469.575 62.320 1470.090 62.460 ;
        RECT 1469.770 62.260 1470.090 62.320 ;
        RECT 634.410 59.400 634.730 59.460 ;
        RECT 1469.785 59.400 1470.075 59.445 ;
        RECT 634.410 59.260 1470.075 59.400 ;
        RECT 634.410 59.200 634.730 59.260 ;
        RECT 1469.785 59.215 1470.075 59.260 ;
      LAYER via ;
        RECT 1470.260 1669.440 1470.520 1669.700 ;
        RECT 1470.720 1580.020 1470.980 1580.280 ;
        RECT 1470.720 1559.620 1470.980 1559.880 ;
        RECT 1470.720 1558.940 1470.980 1559.200 ;
        RECT 1470.720 1365.820 1470.980 1366.080 ;
        RECT 1470.720 1365.140 1470.980 1365.400 ;
        RECT 1470.720 1269.260 1470.980 1269.520 ;
        RECT 1470.720 1268.580 1470.980 1268.840 ;
        RECT 1470.720 1172.700 1470.980 1172.960 ;
        RECT 1470.720 1172.020 1470.980 1172.280 ;
        RECT 1470.720 965.980 1470.980 966.240 ;
        RECT 1471.180 965.640 1471.440 965.900 ;
        RECT 1470.260 917.700 1470.520 917.960 ;
        RECT 1471.180 917.700 1471.440 917.960 ;
        RECT 1470.260 883.360 1470.520 883.620 ;
        RECT 1470.720 882.680 1470.980 882.940 ;
        RECT 1470.720 796.660 1470.980 796.920 ;
        RECT 1471.640 796.660 1471.900 796.920 ;
        RECT 1471.640 793.260 1471.900 793.520 ;
        RECT 1470.260 745.320 1470.520 745.580 ;
        RECT 1470.260 696.700 1470.520 696.960 ;
        RECT 1470.720 607.280 1470.980 607.540 ;
        RECT 1470.720 606.600 1470.980 606.860 ;
        RECT 1470.720 582.800 1470.980 583.060 ;
        RECT 1470.720 400.560 1470.980 400.820 ;
        RECT 1470.720 399.880 1470.980 400.140 ;
        RECT 1469.800 289.720 1470.060 289.980 ;
        RECT 1470.720 289.720 1470.980 289.980 ;
        RECT 1470.720 192.820 1470.980 193.080 ;
        RECT 1470.720 145.220 1470.980 145.480 ;
        RECT 1469.800 144.540 1470.060 144.800 ;
        RECT 1470.720 144.540 1470.980 144.800 ;
        RECT 1469.800 137.740 1470.060 138.000 ;
        RECT 1469.800 89.800 1470.060 90.060 ;
        RECT 1469.800 62.260 1470.060 62.520 ;
        RECT 634.440 59.200 634.700 59.460 ;
      LAYER met2 ;
        RECT 1474.320 1700.410 1474.600 1702.400 ;
        RECT 1471.700 1700.270 1474.600 1700.410 ;
        RECT 1471.700 1676.725 1471.840 1700.270 ;
        RECT 1474.320 1700.000 1474.600 1700.270 ;
        RECT 1470.250 1676.355 1470.530 1676.725 ;
        RECT 1471.630 1676.355 1471.910 1676.725 ;
        RECT 1470.320 1669.730 1470.460 1676.355 ;
        RECT 1470.260 1669.410 1470.520 1669.730 ;
        RECT 1470.720 1579.990 1470.980 1580.310 ;
        RECT 1470.780 1559.910 1470.920 1579.990 ;
        RECT 1470.720 1559.590 1470.980 1559.910 ;
        RECT 1470.720 1558.910 1470.980 1559.230 ;
        RECT 1470.780 1366.110 1470.920 1558.910 ;
        RECT 1470.720 1365.790 1470.980 1366.110 ;
        RECT 1470.720 1365.110 1470.980 1365.430 ;
        RECT 1470.780 1269.550 1470.920 1365.110 ;
        RECT 1470.720 1269.230 1470.980 1269.550 ;
        RECT 1470.720 1268.550 1470.980 1268.870 ;
        RECT 1470.780 1172.990 1470.920 1268.550 ;
        RECT 1470.720 1172.670 1470.980 1172.990 ;
        RECT 1470.720 1171.990 1470.980 1172.310 ;
        RECT 1470.780 1076.850 1470.920 1171.990 ;
        RECT 1470.320 1076.710 1470.920 1076.850 ;
        RECT 1470.320 1076.170 1470.460 1076.710 ;
        RECT 1470.320 1076.030 1470.920 1076.170 ;
        RECT 1470.780 1008.285 1470.920 1076.030 ;
        RECT 1470.710 1007.915 1470.990 1008.285 ;
        RECT 1470.710 1007.235 1470.990 1007.605 ;
        RECT 1470.780 966.270 1470.920 1007.235 ;
        RECT 1470.720 965.950 1470.980 966.270 ;
        RECT 1471.180 965.610 1471.440 965.930 ;
        RECT 1471.240 917.990 1471.380 965.610 ;
        RECT 1470.260 917.670 1470.520 917.990 ;
        RECT 1471.180 917.670 1471.440 917.990 ;
        RECT 1470.320 883.650 1470.460 917.670 ;
        RECT 1470.260 883.330 1470.520 883.650 ;
        RECT 1470.720 882.650 1470.980 882.970 ;
        RECT 1470.780 796.950 1470.920 882.650 ;
        RECT 1470.720 796.630 1470.980 796.950 ;
        RECT 1471.640 796.630 1471.900 796.950 ;
        RECT 1471.700 793.550 1471.840 796.630 ;
        RECT 1471.640 793.230 1471.900 793.550 ;
        RECT 1470.260 745.290 1470.520 745.610 ;
        RECT 1470.320 696.990 1470.460 745.290 ;
        RECT 1470.260 696.670 1470.520 696.990 ;
        RECT 1470.720 607.250 1470.980 607.570 ;
        RECT 1470.780 606.890 1470.920 607.250 ;
        RECT 1470.720 606.570 1470.980 606.890 ;
        RECT 1470.720 582.770 1470.980 583.090 ;
        RECT 1470.780 400.850 1470.920 582.770 ;
        RECT 1470.720 400.530 1470.980 400.850 ;
        RECT 1470.720 399.850 1470.980 400.170 ;
        RECT 1470.780 362.170 1470.920 399.850 ;
        RECT 1469.860 362.030 1470.920 362.170 ;
        RECT 1469.860 290.010 1470.000 362.030 ;
        RECT 1469.800 289.690 1470.060 290.010 ;
        RECT 1470.720 289.690 1470.980 290.010 ;
        RECT 1470.780 193.110 1470.920 289.690 ;
        RECT 1470.720 192.790 1470.980 193.110 ;
        RECT 1470.720 145.190 1470.980 145.510 ;
        RECT 1470.780 144.830 1470.920 145.190 ;
        RECT 1469.800 144.510 1470.060 144.830 ;
        RECT 1470.720 144.510 1470.980 144.830 ;
        RECT 1469.860 138.030 1470.000 144.510 ;
        RECT 1469.800 137.710 1470.060 138.030 ;
        RECT 1469.800 89.770 1470.060 90.090 ;
        RECT 1469.860 62.550 1470.000 89.770 ;
        RECT 1469.800 62.230 1470.060 62.550 ;
        RECT 634.440 59.170 634.700 59.490 ;
        RECT 634.500 17.410 634.640 59.170 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
      LAYER via2 ;
        RECT 1470.250 1676.400 1470.530 1676.680 ;
        RECT 1471.630 1676.400 1471.910 1676.680 ;
        RECT 1470.710 1007.960 1470.990 1008.240 ;
        RECT 1470.710 1007.280 1470.990 1007.560 ;
      LAYER met3 ;
        RECT 1470.225 1676.690 1470.555 1676.705 ;
        RECT 1471.605 1676.690 1471.935 1676.705 ;
        RECT 1470.225 1676.390 1471.935 1676.690 ;
        RECT 1470.225 1676.375 1470.555 1676.390 ;
        RECT 1471.605 1676.375 1471.935 1676.390 ;
        RECT 1470.685 1008.250 1471.015 1008.265 ;
        RECT 1470.685 1007.950 1471.690 1008.250 ;
        RECT 1470.685 1007.935 1471.015 1007.950 ;
        RECT 1470.685 1007.570 1471.015 1007.585 ;
        RECT 1471.390 1007.570 1471.690 1007.950 ;
        RECT 1470.685 1007.270 1471.690 1007.570 ;
        RECT 1470.685 1007.255 1471.015 1007.270 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2392.530 1688.000 2392.850 1688.060 ;
        RECT 2415.990 1688.000 2416.310 1688.060 ;
        RECT 2392.530 1687.860 2416.310 1688.000 ;
        RECT 2392.530 1687.800 2392.850 1687.860 ;
        RECT 2415.990 1687.800 2416.310 1687.860 ;
      LAYER via ;
        RECT 2392.560 1687.800 2392.820 1688.060 ;
        RECT 2416.020 1687.800 2416.280 1688.060 ;
      LAYER met2 ;
        RECT 2392.480 1700.000 2392.760 1702.400 ;
        RECT 2392.620 1688.090 2392.760 1700.000 ;
        RECT 2392.560 1687.770 2392.820 1688.090 ;
        RECT 2416.020 1687.770 2416.280 1688.090 ;
        RECT 2416.080 3.130 2416.220 1687.770 ;
        RECT 2416.080 2.990 2417.600 3.130 ;
        RECT 2417.460 2.400 2417.600 2.990 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2401.730 1688.680 2402.050 1688.740 ;
        RECT 2407.710 1688.680 2408.030 1688.740 ;
        RECT 2401.730 1688.540 2408.030 1688.680 ;
        RECT 2401.730 1688.480 2402.050 1688.540 ;
        RECT 2407.710 1688.480 2408.030 1688.540 ;
        RECT 2407.710 16.560 2408.030 16.620 ;
        RECT 2434.850 16.560 2435.170 16.620 ;
        RECT 2407.710 16.420 2435.170 16.560 ;
        RECT 2407.710 16.360 2408.030 16.420 ;
        RECT 2434.850 16.360 2435.170 16.420 ;
      LAYER via ;
        RECT 2401.760 1688.480 2402.020 1688.740 ;
        RECT 2407.740 1688.480 2408.000 1688.740 ;
        RECT 2407.740 16.360 2408.000 16.620 ;
        RECT 2434.880 16.360 2435.140 16.620 ;
      LAYER met2 ;
        RECT 2401.680 1700.000 2401.960 1702.400 ;
        RECT 2401.820 1688.770 2401.960 1700.000 ;
        RECT 2401.760 1688.450 2402.020 1688.770 ;
        RECT 2407.740 1688.450 2408.000 1688.770 ;
        RECT 2407.800 16.650 2407.940 1688.450 ;
        RECT 2407.740 16.330 2408.000 16.650 ;
        RECT 2434.880 16.330 2435.140 16.650 ;
        RECT 2434.940 2.400 2435.080 16.330 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2414.610 19.280 2414.930 19.340 ;
        RECT 2452.790 19.280 2453.110 19.340 ;
        RECT 2414.610 19.140 2453.110 19.280 ;
        RECT 2414.610 19.080 2414.930 19.140 ;
        RECT 2452.790 19.080 2453.110 19.140 ;
      LAYER via ;
        RECT 2414.640 19.080 2414.900 19.340 ;
        RECT 2452.820 19.080 2453.080 19.340 ;
      LAYER met2 ;
        RECT 2410.880 1700.410 2411.160 1702.400 ;
        RECT 2410.880 1700.270 2413.920 1700.410 ;
        RECT 2410.880 1700.000 2411.160 1700.270 ;
        RECT 2413.780 1688.340 2413.920 1700.270 ;
        RECT 2413.780 1688.200 2414.840 1688.340 ;
        RECT 2414.700 19.370 2414.840 1688.200 ;
        RECT 2414.640 19.050 2414.900 19.370 ;
        RECT 2452.820 19.050 2453.080 19.370 ;
        RECT 2452.880 2.400 2453.020 19.050 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2421.510 17.920 2421.830 17.980 ;
        RECT 2470.730 17.920 2471.050 17.980 ;
        RECT 2421.510 17.780 2471.050 17.920 ;
        RECT 2421.510 17.720 2421.830 17.780 ;
        RECT 2470.730 17.720 2471.050 17.780 ;
      LAYER via ;
        RECT 2421.540 17.720 2421.800 17.980 ;
        RECT 2470.760 17.720 2471.020 17.980 ;
      LAYER met2 ;
        RECT 2420.080 1700.410 2420.360 1702.400 ;
        RECT 2420.080 1700.270 2421.740 1700.410 ;
        RECT 2420.080 1700.000 2420.360 1700.270 ;
        RECT 2421.600 18.010 2421.740 1700.270 ;
        RECT 2421.540 17.690 2421.800 18.010 ;
        RECT 2470.760 17.690 2471.020 18.010 ;
        RECT 2470.820 2.400 2470.960 17.690 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2429.330 1688.340 2429.650 1688.400 ;
        RECT 2445.890 1688.340 2446.210 1688.400 ;
        RECT 2429.330 1688.200 2446.210 1688.340 ;
        RECT 2429.330 1688.140 2429.650 1688.200 ;
        RECT 2445.890 1688.140 2446.210 1688.200 ;
        RECT 2445.890 18.940 2446.210 19.000 ;
        RECT 2488.670 18.940 2488.990 19.000 ;
        RECT 2445.890 18.800 2488.990 18.940 ;
        RECT 2445.890 18.740 2446.210 18.800 ;
        RECT 2488.670 18.740 2488.990 18.800 ;
      LAYER via ;
        RECT 2429.360 1688.140 2429.620 1688.400 ;
        RECT 2445.920 1688.140 2446.180 1688.400 ;
        RECT 2445.920 18.740 2446.180 19.000 ;
        RECT 2488.700 18.740 2488.960 19.000 ;
      LAYER met2 ;
        RECT 2429.280 1700.000 2429.560 1702.400 ;
        RECT 2429.420 1688.430 2429.560 1700.000 ;
        RECT 2429.360 1688.110 2429.620 1688.430 ;
        RECT 2445.920 1688.110 2446.180 1688.430 ;
        RECT 2445.980 19.030 2446.120 1688.110 ;
        RECT 2445.920 18.710 2446.180 19.030 ;
        RECT 2488.700 18.710 2488.960 19.030 ;
        RECT 2488.760 2.400 2488.900 18.710 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2438.530 1685.280 2438.850 1685.340 ;
        RECT 2442.210 1685.280 2442.530 1685.340 ;
        RECT 2438.530 1685.140 2442.530 1685.280 ;
        RECT 2438.530 1685.080 2438.850 1685.140 ;
        RECT 2442.210 1685.080 2442.530 1685.140 ;
        RECT 2442.210 17.240 2442.530 17.300 ;
        RECT 2506.150 17.240 2506.470 17.300 ;
        RECT 2442.210 17.100 2506.470 17.240 ;
        RECT 2442.210 17.040 2442.530 17.100 ;
        RECT 2506.150 17.040 2506.470 17.100 ;
      LAYER via ;
        RECT 2438.560 1685.080 2438.820 1685.340 ;
        RECT 2442.240 1685.080 2442.500 1685.340 ;
        RECT 2442.240 17.040 2442.500 17.300 ;
        RECT 2506.180 17.040 2506.440 17.300 ;
      LAYER met2 ;
        RECT 2438.480 1700.000 2438.760 1702.400 ;
        RECT 2438.620 1685.370 2438.760 1700.000 ;
        RECT 2438.560 1685.050 2438.820 1685.370 ;
        RECT 2442.240 1685.050 2442.500 1685.370 ;
        RECT 2442.300 17.330 2442.440 1685.050 ;
        RECT 2442.240 17.010 2442.500 17.330 ;
        RECT 2506.180 17.010 2506.440 17.330 ;
        RECT 2506.240 2.400 2506.380 17.010 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2449.110 16.220 2449.430 16.280 ;
        RECT 2524.090 16.220 2524.410 16.280 ;
        RECT 2449.110 16.080 2524.410 16.220 ;
        RECT 2449.110 16.020 2449.430 16.080 ;
        RECT 2524.090 16.020 2524.410 16.080 ;
      LAYER via ;
        RECT 2449.140 16.020 2449.400 16.280 ;
        RECT 2524.120 16.020 2524.380 16.280 ;
      LAYER met2 ;
        RECT 2447.680 1700.410 2447.960 1702.400 ;
        RECT 2447.680 1700.270 2449.340 1700.410 ;
        RECT 2447.680 1700.000 2447.960 1700.270 ;
        RECT 2449.200 16.310 2449.340 1700.270 ;
        RECT 2449.140 15.990 2449.400 16.310 ;
        RECT 2524.120 15.990 2524.380 16.310 ;
        RECT 2524.180 2.400 2524.320 15.990 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2456.930 1688.340 2457.250 1688.400 ;
        RECT 2462.910 1688.340 2463.230 1688.400 ;
        RECT 2456.930 1688.200 2463.230 1688.340 ;
        RECT 2456.930 1688.140 2457.250 1688.200 ;
        RECT 2462.910 1688.140 2463.230 1688.200 ;
        RECT 2462.910 16.900 2463.230 16.960 ;
        RECT 2542.030 16.900 2542.350 16.960 ;
        RECT 2462.910 16.760 2542.350 16.900 ;
        RECT 2462.910 16.700 2463.230 16.760 ;
        RECT 2542.030 16.700 2542.350 16.760 ;
      LAYER via ;
        RECT 2456.960 1688.140 2457.220 1688.400 ;
        RECT 2462.940 1688.140 2463.200 1688.400 ;
        RECT 2462.940 16.700 2463.200 16.960 ;
        RECT 2542.060 16.700 2542.320 16.960 ;
      LAYER met2 ;
        RECT 2456.880 1700.000 2457.160 1702.400 ;
        RECT 2457.020 1688.430 2457.160 1700.000 ;
        RECT 2456.960 1688.110 2457.220 1688.430 ;
        RECT 2462.940 1688.110 2463.200 1688.430 ;
        RECT 2463.000 16.990 2463.140 1688.110 ;
        RECT 2462.940 16.670 2463.200 16.990 ;
        RECT 2542.060 16.670 2542.320 16.990 ;
        RECT 2542.120 2.400 2542.260 16.670 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2466.130 1688.340 2466.450 1688.400 ;
        RECT 2469.810 1688.340 2470.130 1688.400 ;
        RECT 2466.130 1688.200 2470.130 1688.340 ;
        RECT 2466.130 1688.140 2466.450 1688.200 ;
        RECT 2469.810 1688.140 2470.130 1688.200 ;
        RECT 2469.810 20.640 2470.130 20.700 ;
        RECT 2559.970 20.640 2560.290 20.700 ;
        RECT 2469.810 20.500 2560.290 20.640 ;
        RECT 2469.810 20.440 2470.130 20.500 ;
        RECT 2559.970 20.440 2560.290 20.500 ;
      LAYER via ;
        RECT 2466.160 1688.140 2466.420 1688.400 ;
        RECT 2469.840 1688.140 2470.100 1688.400 ;
        RECT 2469.840 20.440 2470.100 20.700 ;
        RECT 2560.000 20.440 2560.260 20.700 ;
      LAYER met2 ;
        RECT 2466.080 1700.000 2466.360 1702.400 ;
        RECT 2466.220 1688.430 2466.360 1700.000 ;
        RECT 2466.160 1688.110 2466.420 1688.430 ;
        RECT 2469.840 1688.110 2470.100 1688.430 ;
        RECT 2469.900 20.730 2470.040 1688.110 ;
        RECT 2469.840 20.410 2470.100 20.730 ;
        RECT 2560.000 20.410 2560.260 20.730 ;
        RECT 2560.060 2.400 2560.200 20.410 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2475.330 1685.280 2475.650 1685.340 ;
        RECT 2480.390 1685.280 2480.710 1685.340 ;
        RECT 2475.330 1685.140 2480.710 1685.280 ;
        RECT 2475.330 1685.080 2475.650 1685.140 ;
        RECT 2480.390 1685.080 2480.710 1685.140 ;
        RECT 2480.390 19.620 2480.710 19.680 ;
        RECT 2480.390 19.480 2549.160 19.620 ;
        RECT 2480.390 19.420 2480.710 19.480 ;
        RECT 2549.020 19.280 2549.160 19.480 ;
        RECT 2577.910 19.280 2578.230 19.340 ;
        RECT 2549.020 19.140 2578.230 19.280 ;
        RECT 2577.910 19.080 2578.230 19.140 ;
      LAYER via ;
        RECT 2475.360 1685.080 2475.620 1685.340 ;
        RECT 2480.420 1685.080 2480.680 1685.340 ;
        RECT 2480.420 19.420 2480.680 19.680 ;
        RECT 2577.940 19.080 2578.200 19.340 ;
      LAYER met2 ;
        RECT 2475.280 1700.000 2475.560 1702.400 ;
        RECT 2475.420 1685.370 2475.560 1700.000 ;
        RECT 2475.360 1685.050 2475.620 1685.370 ;
        RECT 2480.420 1685.050 2480.680 1685.370 ;
        RECT 2480.480 19.710 2480.620 1685.050 ;
        RECT 2480.420 19.390 2480.680 19.710 ;
        RECT 2577.940 19.050 2578.200 19.370 ;
        RECT 2578.000 2.400 2578.140 19.050 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 813.810 60.080 814.130 60.140 ;
        RECT 1566.830 60.080 1567.150 60.140 ;
        RECT 813.810 59.940 1567.150 60.080 ;
        RECT 813.810 59.880 814.130 59.940 ;
        RECT 1566.830 59.880 1567.150 59.940 ;
      LAYER via ;
        RECT 813.840 59.880 814.100 60.140 ;
        RECT 1566.860 59.880 1567.120 60.140 ;
      LAYER met2 ;
        RECT 1566.320 1700.410 1566.600 1702.400 ;
        RECT 1566.320 1700.270 1567.060 1700.410 ;
        RECT 1566.320 1700.000 1566.600 1700.270 ;
        RECT 1566.920 60.170 1567.060 1700.270 ;
        RECT 813.840 59.850 814.100 60.170 ;
        RECT 1566.860 59.850 1567.120 60.170 ;
        RECT 813.900 16.730 814.040 59.850 ;
        RECT 811.600 16.590 814.040 16.730 ;
        RECT 811.600 2.400 811.740 16.590 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2484.530 1688.340 2484.850 1688.400 ;
        RECT 2494.190 1688.340 2494.510 1688.400 ;
        RECT 2484.530 1688.200 2494.510 1688.340 ;
        RECT 2484.530 1688.140 2484.850 1688.200 ;
        RECT 2494.190 1688.140 2494.510 1688.200 ;
        RECT 2494.190 18.940 2494.510 19.000 ;
        RECT 2595.390 18.940 2595.710 19.000 ;
        RECT 2494.190 18.800 2595.710 18.940 ;
        RECT 2494.190 18.740 2494.510 18.800 ;
        RECT 2595.390 18.740 2595.710 18.800 ;
      LAYER via ;
        RECT 2484.560 1688.140 2484.820 1688.400 ;
        RECT 2494.220 1688.140 2494.480 1688.400 ;
        RECT 2494.220 18.740 2494.480 19.000 ;
        RECT 2595.420 18.740 2595.680 19.000 ;
      LAYER met2 ;
        RECT 2484.480 1700.000 2484.760 1702.400 ;
        RECT 2484.620 1688.430 2484.760 1700.000 ;
        RECT 2484.560 1688.110 2484.820 1688.430 ;
        RECT 2494.220 1688.110 2494.480 1688.430 ;
        RECT 2494.280 19.030 2494.420 1688.110 ;
        RECT 2494.220 18.710 2494.480 19.030 ;
        RECT 2595.420 18.710 2595.680 19.030 ;
        RECT 2595.480 2.400 2595.620 18.710 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2493.730 1690.040 2494.050 1690.100 ;
        RECT 2497.410 1690.040 2497.730 1690.100 ;
        RECT 2493.730 1689.900 2497.730 1690.040 ;
        RECT 2493.730 1689.840 2494.050 1689.900 ;
        RECT 2497.410 1689.840 2497.730 1689.900 ;
        RECT 2497.410 18.600 2497.730 18.660 ;
        RECT 2613.330 18.600 2613.650 18.660 ;
        RECT 2497.410 18.460 2613.650 18.600 ;
        RECT 2497.410 18.400 2497.730 18.460 ;
        RECT 2613.330 18.400 2613.650 18.460 ;
      LAYER via ;
        RECT 2493.760 1689.840 2494.020 1690.100 ;
        RECT 2497.440 1689.840 2497.700 1690.100 ;
        RECT 2497.440 18.400 2497.700 18.660 ;
        RECT 2613.360 18.400 2613.620 18.660 ;
      LAYER met2 ;
        RECT 2493.680 1700.000 2493.960 1702.400 ;
        RECT 2493.820 1690.130 2493.960 1700.000 ;
        RECT 2493.760 1689.810 2494.020 1690.130 ;
        RECT 2497.440 1689.810 2497.700 1690.130 ;
        RECT 2497.500 18.690 2497.640 1689.810 ;
        RECT 2497.440 18.370 2497.700 18.690 ;
        RECT 2613.360 18.370 2613.620 18.690 ;
        RECT 2613.420 2.400 2613.560 18.370 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2504.310 17.580 2504.630 17.640 ;
        RECT 2631.270 17.580 2631.590 17.640 ;
        RECT 2504.310 17.440 2631.590 17.580 ;
        RECT 2504.310 17.380 2504.630 17.440 ;
        RECT 2631.270 17.380 2631.590 17.440 ;
      LAYER via ;
        RECT 2504.340 17.380 2504.600 17.640 ;
        RECT 2631.300 17.380 2631.560 17.640 ;
      LAYER met2 ;
        RECT 2502.880 1700.410 2503.160 1702.400 ;
        RECT 2502.880 1700.270 2504.540 1700.410 ;
        RECT 2502.880 1700.000 2503.160 1700.270 ;
        RECT 2504.400 17.670 2504.540 1700.270 ;
        RECT 2504.340 17.350 2504.600 17.670 ;
        RECT 2631.300 17.350 2631.560 17.670 ;
        RECT 2631.360 2.400 2631.500 17.350 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2512.130 1688.340 2512.450 1688.400 ;
        RECT 2517.650 1688.340 2517.970 1688.400 ;
        RECT 2512.130 1688.200 2517.970 1688.340 ;
        RECT 2512.130 1688.140 2512.450 1688.200 ;
        RECT 2517.650 1688.140 2517.970 1688.200 ;
        RECT 2517.650 24.720 2517.970 24.780 ;
        RECT 2648.290 24.720 2648.610 24.780 ;
        RECT 2517.650 24.580 2648.610 24.720 ;
        RECT 2517.650 24.520 2517.970 24.580 ;
        RECT 2648.290 24.520 2648.610 24.580 ;
      LAYER via ;
        RECT 2512.160 1688.140 2512.420 1688.400 ;
        RECT 2517.680 1688.140 2517.940 1688.400 ;
        RECT 2517.680 24.520 2517.940 24.780 ;
        RECT 2648.320 24.520 2648.580 24.780 ;
      LAYER met2 ;
        RECT 2512.080 1700.000 2512.360 1702.400 ;
        RECT 2512.220 1688.430 2512.360 1700.000 ;
        RECT 2512.160 1688.110 2512.420 1688.430 ;
        RECT 2517.680 1688.110 2517.940 1688.430 ;
        RECT 2517.740 24.810 2517.880 1688.110 ;
        RECT 2517.680 24.490 2517.940 24.810 ;
        RECT 2648.320 24.490 2648.580 24.810 ;
        RECT 2648.380 16.730 2648.520 24.490 ;
        RECT 2648.380 16.590 2649.440 16.730 ;
        RECT 2649.300 2.400 2649.440 16.590 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2521.330 1688.680 2521.650 1688.740 ;
        RECT 2525.010 1688.680 2525.330 1688.740 ;
        RECT 2521.330 1688.540 2525.330 1688.680 ;
        RECT 2521.330 1688.480 2521.650 1688.540 ;
        RECT 2525.010 1688.480 2525.330 1688.540 ;
        RECT 2525.010 14.520 2525.330 14.580 ;
        RECT 2667.150 14.520 2667.470 14.580 ;
        RECT 2525.010 14.380 2667.470 14.520 ;
        RECT 2525.010 14.320 2525.330 14.380 ;
        RECT 2667.150 14.320 2667.470 14.380 ;
      LAYER via ;
        RECT 2521.360 1688.480 2521.620 1688.740 ;
        RECT 2525.040 1688.480 2525.300 1688.740 ;
        RECT 2525.040 14.320 2525.300 14.580 ;
        RECT 2667.180 14.320 2667.440 14.580 ;
      LAYER met2 ;
        RECT 2521.280 1700.000 2521.560 1702.400 ;
        RECT 2521.420 1688.770 2521.560 1700.000 ;
        RECT 2521.360 1688.450 2521.620 1688.770 ;
        RECT 2525.040 1688.450 2525.300 1688.770 ;
        RECT 2525.100 14.610 2525.240 1688.450 ;
        RECT 2525.040 14.290 2525.300 14.610 ;
        RECT 2667.180 14.290 2667.440 14.610 ;
        RECT 2667.240 2.400 2667.380 14.290 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2531.450 24.040 2531.770 24.100 ;
        RECT 2684.630 24.040 2684.950 24.100 ;
        RECT 2531.450 23.900 2684.950 24.040 ;
        RECT 2531.450 23.840 2531.770 23.900 ;
        RECT 2684.630 23.840 2684.950 23.900 ;
      LAYER via ;
        RECT 2531.480 23.840 2531.740 24.100 ;
        RECT 2684.660 23.840 2684.920 24.100 ;
      LAYER met2 ;
        RECT 2530.480 1700.410 2530.760 1702.400 ;
        RECT 2530.480 1700.270 2531.680 1700.410 ;
        RECT 2530.480 1700.000 2530.760 1700.270 ;
        RECT 2531.540 24.130 2531.680 1700.270 ;
        RECT 2531.480 23.810 2531.740 24.130 ;
        RECT 2684.660 23.810 2684.920 24.130 ;
        RECT 2684.720 2.400 2684.860 23.810 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2539.730 1688.680 2540.050 1688.740 ;
        RECT 2545.710 1688.680 2546.030 1688.740 ;
        RECT 2539.730 1688.540 2546.030 1688.680 ;
        RECT 2539.730 1688.480 2540.050 1688.540 ;
        RECT 2545.710 1688.480 2546.030 1688.540 ;
        RECT 2545.710 24.380 2546.030 24.440 ;
        RECT 2702.570 24.380 2702.890 24.440 ;
        RECT 2545.710 24.240 2702.890 24.380 ;
        RECT 2545.710 24.180 2546.030 24.240 ;
        RECT 2702.570 24.180 2702.890 24.240 ;
      LAYER via ;
        RECT 2539.760 1688.480 2540.020 1688.740 ;
        RECT 2545.740 1688.480 2546.000 1688.740 ;
        RECT 2545.740 24.180 2546.000 24.440 ;
        RECT 2702.600 24.180 2702.860 24.440 ;
      LAYER met2 ;
        RECT 2539.680 1700.000 2539.960 1702.400 ;
        RECT 2539.820 1688.770 2539.960 1700.000 ;
        RECT 2539.760 1688.450 2540.020 1688.770 ;
        RECT 2545.740 1688.450 2546.000 1688.770 ;
        RECT 2545.800 24.470 2545.940 1688.450 ;
        RECT 2545.740 24.150 2546.000 24.470 ;
        RECT 2702.600 24.150 2702.860 24.470 ;
        RECT 2702.660 2.400 2702.800 24.150 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2548.930 1685.280 2549.250 1685.340 ;
        RECT 2701.650 1685.280 2701.970 1685.340 ;
        RECT 2548.930 1685.140 2701.970 1685.280 ;
        RECT 2548.930 1685.080 2549.250 1685.140 ;
        RECT 2701.650 1685.080 2701.970 1685.140 ;
        RECT 2701.650 15.880 2701.970 15.940 ;
        RECT 2720.510 15.880 2720.830 15.940 ;
        RECT 2701.650 15.740 2720.830 15.880 ;
        RECT 2701.650 15.680 2701.970 15.740 ;
        RECT 2720.510 15.680 2720.830 15.740 ;
      LAYER via ;
        RECT 2548.960 1685.080 2549.220 1685.340 ;
        RECT 2701.680 1685.080 2701.940 1685.340 ;
        RECT 2701.680 15.680 2701.940 15.940 ;
        RECT 2720.540 15.680 2720.800 15.940 ;
      LAYER met2 ;
        RECT 2548.880 1700.000 2549.160 1702.400 ;
        RECT 2549.020 1685.370 2549.160 1700.000 ;
        RECT 2548.960 1685.050 2549.220 1685.370 ;
        RECT 2701.680 1685.050 2701.940 1685.370 ;
        RECT 2701.740 15.970 2701.880 1685.050 ;
        RECT 2701.680 15.650 2701.940 15.970 ;
        RECT 2720.540 15.650 2720.800 15.970 ;
        RECT 2720.600 2.400 2720.740 15.650 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2700.805 14.705 2700.975 16.235 ;
      LAYER mcon ;
        RECT 2700.805 16.065 2700.975 16.235 ;
      LAYER met1 ;
        RECT 2559.050 16.220 2559.370 16.280 ;
        RECT 2700.745 16.220 2701.035 16.265 ;
        RECT 2559.050 16.080 2701.035 16.220 ;
        RECT 2559.050 16.020 2559.370 16.080 ;
        RECT 2700.745 16.035 2701.035 16.080 ;
        RECT 2700.745 14.860 2701.035 14.905 ;
        RECT 2738.450 14.860 2738.770 14.920 ;
        RECT 2700.745 14.720 2738.770 14.860 ;
        RECT 2700.745 14.675 2701.035 14.720 ;
        RECT 2738.450 14.660 2738.770 14.720 ;
      LAYER via ;
        RECT 2559.080 16.020 2559.340 16.280 ;
        RECT 2738.480 14.660 2738.740 14.920 ;
      LAYER met2 ;
        RECT 2558.080 1700.410 2558.360 1702.400 ;
        RECT 2558.080 1700.270 2559.280 1700.410 ;
        RECT 2558.080 1700.000 2558.360 1700.270 ;
        RECT 2559.140 16.310 2559.280 1700.270 ;
        RECT 2559.080 15.990 2559.340 16.310 ;
        RECT 2738.480 14.630 2738.740 14.950 ;
        RECT 2738.540 2.400 2738.680 14.630 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2618.005 1684.105 2618.175 1687.675 ;
      LAYER mcon ;
        RECT 2618.005 1687.505 2618.175 1687.675 ;
      LAYER met1 ;
        RECT 2569.170 1687.660 2569.490 1687.720 ;
        RECT 2617.945 1687.660 2618.235 1687.705 ;
        RECT 2569.170 1687.520 2618.235 1687.660 ;
        RECT 2569.170 1687.460 2569.490 1687.520 ;
        RECT 2617.945 1687.475 2618.235 1687.520 ;
        RECT 2617.945 1684.260 2618.235 1684.305 ;
        RECT 2714.990 1684.260 2715.310 1684.320 ;
        RECT 2617.945 1684.120 2715.310 1684.260 ;
        RECT 2617.945 1684.075 2618.235 1684.120 ;
        RECT 2714.990 1684.060 2715.310 1684.120 ;
        RECT 2755.930 14.860 2756.250 14.920 ;
        RECT 2739.000 14.720 2756.250 14.860 ;
        RECT 2714.990 14.180 2715.310 14.240 ;
        RECT 2739.000 14.180 2739.140 14.720 ;
        RECT 2755.930 14.660 2756.250 14.720 ;
        RECT 2714.990 14.040 2739.140 14.180 ;
        RECT 2714.990 13.980 2715.310 14.040 ;
      LAYER via ;
        RECT 2569.200 1687.460 2569.460 1687.720 ;
        RECT 2715.020 1684.060 2715.280 1684.320 ;
        RECT 2715.020 13.980 2715.280 14.240 ;
        RECT 2755.960 14.660 2756.220 14.920 ;
      LAYER met2 ;
        RECT 2567.280 1700.410 2567.560 1702.400 ;
        RECT 2567.280 1700.270 2569.400 1700.410 ;
        RECT 2567.280 1700.000 2567.560 1700.270 ;
        RECT 2569.260 1687.750 2569.400 1700.270 ;
        RECT 2569.200 1687.430 2569.460 1687.750 ;
        RECT 2715.020 1684.030 2715.280 1684.350 ;
        RECT 2715.080 14.270 2715.220 1684.030 ;
        RECT 2755.960 14.630 2756.220 14.950 ;
        RECT 2715.020 13.950 2715.280 14.270 ;
        RECT 2756.020 2.400 2756.160 14.630 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.510 60.420 834.830 60.480 ;
        RECT 1573.730 60.420 1574.050 60.480 ;
        RECT 834.510 60.280 1574.050 60.420 ;
        RECT 834.510 60.220 834.830 60.280 ;
        RECT 1573.730 60.220 1574.050 60.280 ;
      LAYER via ;
        RECT 834.540 60.220 834.800 60.480 ;
        RECT 1573.760 60.220 1574.020 60.480 ;
      LAYER met2 ;
        RECT 1575.520 1700.410 1575.800 1702.400 ;
        RECT 1573.820 1700.270 1575.800 1700.410 ;
        RECT 1573.820 60.510 1573.960 1700.270 ;
        RECT 1575.520 1700.000 1575.800 1700.270 ;
        RECT 834.540 60.190 834.800 60.510 ;
        RECT 1573.760 60.190 1574.020 60.510 ;
        RECT 834.600 16.730 834.740 60.190 ;
        RECT 829.540 16.590 834.740 16.730 ;
        RECT 829.540 2.400 829.680 16.590 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2618.465 1684.785 2618.635 1685.975 ;
      LAYER mcon ;
        RECT 2618.465 1685.805 2618.635 1685.975 ;
      LAYER met1 ;
        RECT 2576.530 1685.960 2576.850 1686.020 ;
        RECT 2618.405 1685.960 2618.695 1686.005 ;
        RECT 2576.530 1685.820 2618.695 1685.960 ;
        RECT 2576.530 1685.760 2576.850 1685.820 ;
        RECT 2618.405 1685.775 2618.695 1685.820 ;
        RECT 2618.405 1684.940 2618.695 1684.985 ;
        RECT 2728.790 1684.940 2729.110 1685.000 ;
        RECT 2618.405 1684.800 2729.110 1684.940 ;
        RECT 2618.405 1684.755 2618.695 1684.800 ;
        RECT 2728.790 1684.740 2729.110 1684.800 ;
        RECT 2728.790 15.540 2729.110 15.600 ;
        RECT 2773.870 15.540 2774.190 15.600 ;
        RECT 2728.790 15.400 2774.190 15.540 ;
        RECT 2728.790 15.340 2729.110 15.400 ;
        RECT 2773.870 15.340 2774.190 15.400 ;
      LAYER via ;
        RECT 2576.560 1685.760 2576.820 1686.020 ;
        RECT 2728.820 1684.740 2729.080 1685.000 ;
        RECT 2728.820 15.340 2729.080 15.600 ;
        RECT 2773.900 15.340 2774.160 15.600 ;
      LAYER met2 ;
        RECT 2576.480 1700.000 2576.760 1702.400 ;
        RECT 2576.620 1686.050 2576.760 1700.000 ;
        RECT 2576.560 1685.730 2576.820 1686.050 ;
        RECT 2728.820 1684.710 2729.080 1685.030 ;
        RECT 2728.880 15.630 2729.020 1684.710 ;
        RECT 2728.820 15.310 2729.080 15.630 ;
        RECT 2773.900 15.310 2774.160 15.630 ;
        RECT 2773.960 2.400 2774.100 15.310 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2585.730 1686.640 2586.050 1686.700 ;
        RECT 2749.490 1686.640 2749.810 1686.700 ;
        RECT 2585.730 1686.500 2749.810 1686.640 ;
        RECT 2585.730 1686.440 2586.050 1686.500 ;
        RECT 2749.490 1686.440 2749.810 1686.500 ;
        RECT 2791.810 16.220 2792.130 16.280 ;
        RECT 2774.420 16.080 2792.130 16.220 ;
        RECT 2749.490 15.200 2749.810 15.260 ;
        RECT 2774.420 15.200 2774.560 16.080 ;
        RECT 2791.810 16.020 2792.130 16.080 ;
        RECT 2749.490 15.060 2774.560 15.200 ;
        RECT 2749.490 15.000 2749.810 15.060 ;
      LAYER via ;
        RECT 2585.760 1686.440 2586.020 1686.700 ;
        RECT 2749.520 1686.440 2749.780 1686.700 ;
        RECT 2749.520 15.000 2749.780 15.260 ;
        RECT 2791.840 16.020 2792.100 16.280 ;
      LAYER met2 ;
        RECT 2585.680 1700.000 2585.960 1702.400 ;
        RECT 2585.820 1686.730 2585.960 1700.000 ;
        RECT 2585.760 1686.410 2586.020 1686.730 ;
        RECT 2749.520 1686.410 2749.780 1686.730 ;
        RECT 2749.580 15.290 2749.720 1686.410 ;
        RECT 2791.840 15.990 2792.100 16.310 ;
        RECT 2749.520 14.970 2749.780 15.290 ;
        RECT 2791.900 2.400 2792.040 15.990 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2594.930 1688.000 2595.250 1688.060 ;
        RECT 2600.450 1688.000 2600.770 1688.060 ;
        RECT 2594.930 1687.860 2600.770 1688.000 ;
        RECT 2594.930 1687.800 2595.250 1687.860 ;
        RECT 2600.450 1687.800 2600.770 1687.860 ;
        RECT 2600.450 20.300 2600.770 20.360 ;
        RECT 2809.750 20.300 2810.070 20.360 ;
        RECT 2600.450 20.160 2810.070 20.300 ;
        RECT 2600.450 20.100 2600.770 20.160 ;
        RECT 2809.750 20.100 2810.070 20.160 ;
      LAYER via ;
        RECT 2594.960 1687.800 2595.220 1688.060 ;
        RECT 2600.480 1687.800 2600.740 1688.060 ;
        RECT 2600.480 20.100 2600.740 20.360 ;
        RECT 2809.780 20.100 2810.040 20.360 ;
      LAYER met2 ;
        RECT 2594.880 1700.000 2595.160 1702.400 ;
        RECT 2595.020 1688.090 2595.160 1700.000 ;
        RECT 2594.960 1687.770 2595.220 1688.090 ;
        RECT 2600.480 1687.770 2600.740 1688.090 ;
        RECT 2600.540 20.390 2600.680 1687.770 ;
        RECT 2600.480 20.070 2600.740 20.390 ;
        RECT 2809.780 20.070 2810.040 20.390 ;
        RECT 2809.840 2.400 2809.980 20.070 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2604.130 1689.360 2604.450 1689.420 ;
        RECT 2783.990 1689.360 2784.310 1689.420 ;
        RECT 2604.130 1689.220 2784.310 1689.360 ;
        RECT 2604.130 1689.160 2604.450 1689.220 ;
        RECT 2783.990 1689.160 2784.310 1689.220 ;
        RECT 2783.990 16.560 2784.310 16.620 ;
        RECT 2827.690 16.560 2828.010 16.620 ;
        RECT 2783.990 16.420 2828.010 16.560 ;
        RECT 2783.990 16.360 2784.310 16.420 ;
        RECT 2827.690 16.360 2828.010 16.420 ;
      LAYER via ;
        RECT 2604.160 1689.160 2604.420 1689.420 ;
        RECT 2784.020 1689.160 2784.280 1689.420 ;
        RECT 2784.020 16.360 2784.280 16.620 ;
        RECT 2827.720 16.360 2827.980 16.620 ;
      LAYER met2 ;
        RECT 2604.080 1700.000 2604.360 1702.400 ;
        RECT 2604.220 1689.450 2604.360 1700.000 ;
        RECT 2604.160 1689.130 2604.420 1689.450 ;
        RECT 2784.020 1689.130 2784.280 1689.450 ;
        RECT 2784.080 16.650 2784.220 1689.130 ;
        RECT 2784.020 16.330 2784.280 16.650 ;
        RECT 2827.720 16.330 2827.980 16.650 ;
        RECT 2827.780 2.400 2827.920 16.330 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2614.710 18.940 2615.030 19.000 ;
        RECT 2845.170 18.940 2845.490 19.000 ;
        RECT 2614.710 18.800 2845.490 18.940 ;
        RECT 2614.710 18.740 2615.030 18.800 ;
        RECT 2845.170 18.740 2845.490 18.800 ;
      LAYER via ;
        RECT 2614.740 18.740 2615.000 19.000 ;
        RECT 2845.200 18.740 2845.460 19.000 ;
      LAYER met2 ;
        RECT 2613.280 1700.410 2613.560 1702.400 ;
        RECT 2613.280 1700.270 2614.940 1700.410 ;
        RECT 2613.280 1700.000 2613.560 1700.270 ;
        RECT 2614.800 19.030 2614.940 1700.270 ;
        RECT 2614.740 18.710 2615.000 19.030 ;
        RECT 2845.200 18.710 2845.460 19.030 ;
        RECT 2845.260 2.400 2845.400 18.710 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2622.530 1683.920 2622.850 1683.980 ;
        RECT 2628.050 1683.920 2628.370 1683.980 ;
        RECT 2622.530 1683.780 2628.370 1683.920 ;
        RECT 2622.530 1683.720 2622.850 1683.780 ;
        RECT 2628.050 1683.720 2628.370 1683.780 ;
        RECT 2628.050 19.280 2628.370 19.340 ;
        RECT 2863.110 19.280 2863.430 19.340 ;
        RECT 2628.050 19.140 2863.430 19.280 ;
        RECT 2628.050 19.080 2628.370 19.140 ;
        RECT 2863.110 19.080 2863.430 19.140 ;
      LAYER via ;
        RECT 2622.560 1683.720 2622.820 1683.980 ;
        RECT 2628.080 1683.720 2628.340 1683.980 ;
        RECT 2628.080 19.080 2628.340 19.340 ;
        RECT 2863.140 19.080 2863.400 19.340 ;
      LAYER met2 ;
        RECT 2622.480 1700.000 2622.760 1702.400 ;
        RECT 2622.620 1684.010 2622.760 1700.000 ;
        RECT 2622.560 1683.690 2622.820 1684.010 ;
        RECT 2628.080 1683.690 2628.340 1684.010 ;
        RECT 2628.140 19.370 2628.280 1683.690 ;
        RECT 2628.080 19.050 2628.340 19.370 ;
        RECT 2863.140 19.050 2863.400 19.370 ;
        RECT 2863.200 2.400 2863.340 19.050 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2643.305 1685.805 2649.455 1685.975 ;
      LAYER mcon ;
        RECT 2649.285 1685.805 2649.455 1685.975 ;
      LAYER met1 ;
        RECT 2634.030 1685.960 2634.350 1686.020 ;
        RECT 2643.245 1685.960 2643.535 1686.005 ;
        RECT 2634.030 1685.820 2643.535 1685.960 ;
        RECT 2634.030 1685.760 2634.350 1685.820 ;
        RECT 2643.245 1685.775 2643.535 1685.820 ;
        RECT 2649.225 1685.960 2649.515 1686.005 ;
        RECT 2790.890 1685.960 2791.210 1686.020 ;
        RECT 2649.225 1685.820 2791.210 1685.960 ;
        RECT 2649.225 1685.775 2649.515 1685.820 ;
        RECT 2790.890 1685.760 2791.210 1685.820 ;
        RECT 2790.890 16.900 2791.210 16.960 ;
        RECT 2790.890 16.760 2845.860 16.900 ;
        RECT 2790.890 16.700 2791.210 16.760 ;
        RECT 2845.720 16.220 2845.860 16.760 ;
        RECT 2881.050 16.220 2881.370 16.280 ;
        RECT 2845.720 16.080 2881.370 16.220 ;
        RECT 2881.050 16.020 2881.370 16.080 ;
      LAYER via ;
        RECT 2634.060 1685.760 2634.320 1686.020 ;
        RECT 2790.920 1685.760 2791.180 1686.020 ;
        RECT 2790.920 16.700 2791.180 16.960 ;
        RECT 2881.080 16.020 2881.340 16.280 ;
      LAYER met2 ;
        RECT 2631.680 1700.410 2631.960 1702.400 ;
        RECT 2631.680 1700.270 2634.260 1700.410 ;
        RECT 2631.680 1700.000 2631.960 1700.270 ;
        RECT 2634.120 1686.050 2634.260 1700.270 ;
        RECT 2634.060 1685.730 2634.320 1686.050 ;
        RECT 2790.920 1685.730 2791.180 1686.050 ;
        RECT 2790.980 16.990 2791.120 1685.730 ;
        RECT 2790.920 16.670 2791.180 16.990 ;
        RECT 2881.080 15.990 2881.340 16.310 ;
        RECT 2881.140 2.400 2881.280 15.990 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2825.390 19.960 2825.710 20.020 ;
        RECT 2898.990 19.960 2899.310 20.020 ;
        RECT 2825.390 19.820 2899.310 19.960 ;
        RECT 2825.390 19.760 2825.710 19.820 ;
        RECT 2898.990 19.760 2899.310 19.820 ;
      LAYER via ;
        RECT 2825.420 19.760 2825.680 20.020 ;
        RECT 2899.020 19.760 2899.280 20.020 ;
      LAYER met2 ;
        RECT 2640.880 1700.000 2641.160 1702.400 ;
        RECT 2641.020 1686.925 2641.160 1700.000 ;
        RECT 2640.950 1686.555 2641.230 1686.925 ;
        RECT 2825.410 1686.555 2825.690 1686.925 ;
        RECT 2825.480 20.050 2825.620 1686.555 ;
        RECT 2825.420 19.730 2825.680 20.050 ;
        RECT 2899.020 19.730 2899.280 20.050 ;
        RECT 2899.080 2.400 2899.220 19.730 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 2640.950 1686.600 2641.230 1686.880 ;
        RECT 2825.410 1686.600 2825.690 1686.880 ;
      LAYER met3 ;
        RECT 2640.925 1686.890 2641.255 1686.905 ;
        RECT 2825.385 1686.890 2825.715 1686.905 ;
        RECT 2640.925 1686.590 2825.715 1686.890 ;
        RECT 2640.925 1686.575 2641.255 1686.590 ;
        RECT 2825.385 1686.575 2825.715 1686.590 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1580.170 1689.700 1580.490 1689.760 ;
        RECT 1583.390 1689.700 1583.710 1689.760 ;
        RECT 1580.170 1689.560 1583.710 1689.700 ;
        RECT 1580.170 1689.500 1580.490 1689.560 ;
        RECT 1583.390 1689.500 1583.710 1689.560 ;
        RECT 848.310 60.760 848.630 60.820 ;
        RECT 1580.170 60.760 1580.490 60.820 ;
        RECT 848.310 60.620 1580.490 60.760 ;
        RECT 848.310 60.560 848.630 60.620 ;
        RECT 1580.170 60.560 1580.490 60.620 ;
      LAYER via ;
        RECT 1580.200 1689.500 1580.460 1689.760 ;
        RECT 1583.420 1689.500 1583.680 1689.760 ;
        RECT 848.340 60.560 848.600 60.820 ;
        RECT 1580.200 60.560 1580.460 60.820 ;
      LAYER met2 ;
        RECT 1584.720 1700.410 1585.000 1702.400 ;
        RECT 1583.480 1700.270 1585.000 1700.410 ;
        RECT 1583.480 1689.790 1583.620 1700.270 ;
        RECT 1584.720 1700.000 1585.000 1700.270 ;
        RECT 1580.200 1689.470 1580.460 1689.790 ;
        RECT 1583.420 1689.470 1583.680 1689.790 ;
        RECT 1580.260 60.850 1580.400 1689.470 ;
        RECT 848.340 60.530 848.600 60.850 ;
        RECT 1580.200 60.530 1580.460 60.850 ;
        RECT 848.400 16.730 848.540 60.530 ;
        RECT 847.020 16.590 848.540 16.730 ;
        RECT 847.020 2.400 847.160 16.590 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1587.990 1689.700 1588.310 1689.760 ;
        RECT 1591.670 1689.700 1591.990 1689.760 ;
        RECT 1587.990 1689.560 1591.990 1689.700 ;
        RECT 1587.990 1689.500 1588.310 1689.560 ;
        RECT 1591.670 1689.500 1591.990 1689.560 ;
        RECT 869.010 61.100 869.330 61.160 ;
        RECT 1587.990 61.100 1588.310 61.160 ;
        RECT 869.010 60.960 1588.310 61.100 ;
        RECT 869.010 60.900 869.330 60.960 ;
        RECT 1587.990 60.900 1588.310 60.960 ;
        RECT 864.870 2.960 865.190 3.020 ;
        RECT 869.010 2.960 869.330 3.020 ;
        RECT 864.870 2.820 869.330 2.960 ;
        RECT 864.870 2.760 865.190 2.820 ;
        RECT 869.010 2.760 869.330 2.820 ;
      LAYER via ;
        RECT 1588.020 1689.500 1588.280 1689.760 ;
        RECT 1591.700 1689.500 1591.960 1689.760 ;
        RECT 869.040 60.900 869.300 61.160 ;
        RECT 1588.020 60.900 1588.280 61.160 ;
        RECT 864.900 2.760 865.160 3.020 ;
        RECT 869.040 2.760 869.300 3.020 ;
      LAYER met2 ;
        RECT 1593.460 1700.410 1593.740 1702.400 ;
        RECT 1591.760 1700.270 1593.740 1700.410 ;
        RECT 1591.760 1689.790 1591.900 1700.270 ;
        RECT 1593.460 1700.000 1593.740 1700.270 ;
        RECT 1588.020 1689.470 1588.280 1689.790 ;
        RECT 1591.700 1689.470 1591.960 1689.790 ;
        RECT 1588.080 61.190 1588.220 1689.470 ;
        RECT 869.040 60.870 869.300 61.190 ;
        RECT 1588.020 60.870 1588.280 61.190 ;
        RECT 869.100 3.050 869.240 60.870 ;
        RECT 864.900 2.730 865.160 3.050 ;
        RECT 869.040 2.730 869.300 3.050 ;
        RECT 864.960 2.400 865.100 2.730 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 61.440 883.130 61.500 ;
        RECT 1601.330 61.440 1601.650 61.500 ;
        RECT 882.810 61.300 1601.650 61.440 ;
        RECT 882.810 61.240 883.130 61.300 ;
        RECT 1601.330 61.240 1601.650 61.300 ;
      LAYER via ;
        RECT 882.840 61.240 883.100 61.500 ;
        RECT 1601.360 61.240 1601.620 61.500 ;
      LAYER met2 ;
        RECT 1602.660 1700.410 1602.940 1702.400 ;
        RECT 1601.420 1700.270 1602.940 1700.410 ;
        RECT 1601.420 61.530 1601.560 1700.270 ;
        RECT 1602.660 1700.000 1602.940 1700.270 ;
        RECT 882.840 61.210 883.100 61.530 ;
        RECT 1601.360 61.210 1601.620 61.530 ;
        RECT 882.900 2.400 883.040 61.210 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1608.765 717.825 1608.935 765.935 ;
        RECT 1608.765 614.125 1608.935 662.235 ;
        RECT 1608.305 89.845 1608.475 137.955 ;
      LAYER mcon ;
        RECT 1608.765 765.765 1608.935 765.935 ;
        RECT 1608.765 662.065 1608.935 662.235 ;
        RECT 1608.305 137.785 1608.475 137.955 ;
      LAYER met1 ;
        RECT 1608.690 931.840 1609.010 931.900 ;
        RECT 1608.320 931.700 1609.010 931.840 ;
        RECT 1608.320 931.560 1608.460 931.700 ;
        RECT 1608.690 931.640 1609.010 931.700 ;
        RECT 1608.230 931.300 1608.550 931.560 ;
        RECT 1608.230 883.360 1608.550 883.620 ;
        RECT 1608.320 882.880 1608.460 883.360 ;
        RECT 1608.690 882.880 1609.010 882.940 ;
        RECT 1608.320 882.740 1609.010 882.880 ;
        RECT 1608.690 882.680 1609.010 882.740 ;
        RECT 1608.690 765.920 1609.010 765.980 ;
        RECT 1608.495 765.780 1609.010 765.920 ;
        RECT 1608.690 765.720 1609.010 765.780 ;
        RECT 1608.690 717.980 1609.010 718.040 ;
        RECT 1608.495 717.840 1609.010 717.980 ;
        RECT 1608.690 717.780 1609.010 717.840 ;
        RECT 1608.690 662.220 1609.010 662.280 ;
        RECT 1608.495 662.080 1609.010 662.220 ;
        RECT 1608.690 662.020 1609.010 662.080 ;
        RECT 1608.690 614.280 1609.010 614.340 ;
        RECT 1608.495 614.140 1609.010 614.280 ;
        RECT 1608.690 614.080 1609.010 614.140 ;
        RECT 1608.690 593.680 1609.010 593.940 ;
        RECT 1608.780 593.260 1608.920 593.680 ;
        RECT 1608.690 593.000 1609.010 593.260 ;
        RECT 1608.690 497.120 1609.010 497.380 ;
        RECT 1608.780 496.700 1608.920 497.120 ;
        RECT 1608.690 496.440 1609.010 496.700 ;
        RECT 1608.230 137.940 1608.550 138.000 ;
        RECT 1608.035 137.800 1608.550 137.940 ;
        RECT 1608.230 137.740 1608.550 137.800 ;
        RECT 1608.245 90.000 1608.535 90.045 ;
        RECT 1608.690 90.000 1609.010 90.060 ;
        RECT 1608.245 89.860 1609.010 90.000 ;
        RECT 1608.245 89.815 1608.535 89.860 ;
        RECT 1608.690 89.800 1609.010 89.860 ;
        RECT 903.510 61.780 903.830 61.840 ;
        RECT 1608.690 61.780 1609.010 61.840 ;
        RECT 903.510 61.640 1609.010 61.780 ;
        RECT 903.510 61.580 903.830 61.640 ;
        RECT 1608.690 61.580 1609.010 61.640 ;
        RECT 900.750 2.960 901.070 3.020 ;
        RECT 903.510 2.960 903.830 3.020 ;
        RECT 900.750 2.820 903.830 2.960 ;
        RECT 900.750 2.760 901.070 2.820 ;
        RECT 903.510 2.760 903.830 2.820 ;
      LAYER via ;
        RECT 1608.720 931.640 1608.980 931.900 ;
        RECT 1608.260 931.300 1608.520 931.560 ;
        RECT 1608.260 883.360 1608.520 883.620 ;
        RECT 1608.720 882.680 1608.980 882.940 ;
        RECT 1608.720 765.720 1608.980 765.980 ;
        RECT 1608.720 717.780 1608.980 718.040 ;
        RECT 1608.720 662.020 1608.980 662.280 ;
        RECT 1608.720 614.080 1608.980 614.340 ;
        RECT 1608.720 593.680 1608.980 593.940 ;
        RECT 1608.720 593.000 1608.980 593.260 ;
        RECT 1608.720 497.120 1608.980 497.380 ;
        RECT 1608.720 496.440 1608.980 496.700 ;
        RECT 1608.260 137.740 1608.520 138.000 ;
        RECT 1608.720 89.800 1608.980 90.060 ;
        RECT 903.540 61.580 903.800 61.840 ;
        RECT 1608.720 61.580 1608.980 61.840 ;
        RECT 900.780 2.760 901.040 3.020 ;
        RECT 903.540 2.760 903.800 3.020 ;
      LAYER met2 ;
        RECT 1611.860 1700.410 1612.140 1702.400 ;
        RECT 1610.620 1700.270 1612.140 1700.410 ;
        RECT 1610.620 1656.210 1610.760 1700.270 ;
        RECT 1611.860 1700.000 1612.140 1700.270 ;
        RECT 1608.780 1656.070 1610.760 1656.210 ;
        RECT 1608.780 980.290 1608.920 1656.070 ;
        RECT 1608.320 980.150 1608.920 980.290 ;
        RECT 1608.320 979.610 1608.460 980.150 ;
        RECT 1608.320 979.470 1608.920 979.610 ;
        RECT 1608.780 931.930 1608.920 979.470 ;
        RECT 1608.720 931.610 1608.980 931.930 ;
        RECT 1608.260 931.270 1608.520 931.590 ;
        RECT 1608.320 883.650 1608.460 931.270 ;
        RECT 1608.260 883.330 1608.520 883.650 ;
        RECT 1608.720 882.650 1608.980 882.970 ;
        RECT 1608.780 787.170 1608.920 882.650 ;
        RECT 1608.320 787.030 1608.920 787.170 ;
        RECT 1608.320 786.490 1608.460 787.030 ;
        RECT 1608.320 786.350 1608.920 786.490 ;
        RECT 1608.780 766.010 1608.920 786.350 ;
        RECT 1608.720 765.690 1608.980 766.010 ;
        RECT 1608.720 717.750 1608.980 718.070 ;
        RECT 1608.780 663.410 1608.920 717.750 ;
        RECT 1608.320 663.270 1608.920 663.410 ;
        RECT 1608.320 662.730 1608.460 663.270 ;
        RECT 1608.320 662.590 1608.920 662.730 ;
        RECT 1608.780 662.310 1608.920 662.590 ;
        RECT 1608.720 661.990 1608.980 662.310 ;
        RECT 1608.720 614.050 1608.980 614.370 ;
        RECT 1608.780 593.970 1608.920 614.050 ;
        RECT 1608.720 593.650 1608.980 593.970 ;
        RECT 1608.720 592.970 1608.980 593.290 ;
        RECT 1608.780 497.410 1608.920 592.970 ;
        RECT 1608.720 497.090 1608.980 497.410 ;
        RECT 1608.720 496.410 1608.980 496.730 ;
        RECT 1608.780 362.170 1608.920 496.410 ;
        RECT 1608.320 362.030 1608.920 362.170 ;
        RECT 1608.320 290.770 1608.460 362.030 ;
        RECT 1608.320 290.630 1608.920 290.770 ;
        RECT 1608.780 289.410 1608.920 290.630 ;
        RECT 1608.320 289.270 1608.920 289.410 ;
        RECT 1608.320 138.030 1608.460 289.270 ;
        RECT 1608.260 137.710 1608.520 138.030 ;
        RECT 1608.720 89.770 1608.980 90.090 ;
        RECT 1608.780 61.870 1608.920 89.770 ;
        RECT 903.540 61.550 903.800 61.870 ;
        RECT 1608.720 61.550 1608.980 61.870 ;
        RECT 903.600 3.050 903.740 61.550 ;
        RECT 900.780 2.730 901.040 3.050 ;
        RECT 903.540 2.730 903.800 3.050 ;
        RECT 900.840 2.400 900.980 2.730 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1615.590 1678.140 1615.910 1678.200 ;
        RECT 1619.270 1678.140 1619.590 1678.200 ;
        RECT 1615.590 1678.000 1619.590 1678.140 ;
        RECT 1615.590 1677.940 1615.910 1678.000 ;
        RECT 1619.270 1677.940 1619.590 1678.000 ;
        RECT 924.210 62.120 924.530 62.180 ;
        RECT 1615.590 62.120 1615.910 62.180 ;
        RECT 924.210 61.980 1615.910 62.120 ;
        RECT 924.210 61.920 924.530 61.980 ;
        RECT 1615.590 61.920 1615.910 61.980 ;
      LAYER via ;
        RECT 1615.620 1677.940 1615.880 1678.200 ;
        RECT 1619.300 1677.940 1619.560 1678.200 ;
        RECT 924.240 61.920 924.500 62.180 ;
        RECT 1615.620 61.920 1615.880 62.180 ;
      LAYER met2 ;
        RECT 1621.060 1700.410 1621.340 1702.400 ;
        RECT 1619.360 1700.270 1621.340 1700.410 ;
        RECT 1619.360 1678.230 1619.500 1700.270 ;
        RECT 1621.060 1700.000 1621.340 1700.270 ;
        RECT 1615.620 1677.910 1615.880 1678.230 ;
        RECT 1619.300 1677.910 1619.560 1678.230 ;
        RECT 1615.680 62.210 1615.820 1677.910 ;
        RECT 924.240 61.890 924.500 62.210 ;
        RECT 1615.620 61.890 1615.880 62.210 ;
        RECT 924.300 29.650 924.440 61.890 ;
        RECT 918.780 29.510 924.440 29.650 ;
        RECT 918.780 2.400 918.920 29.510 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 938.010 58.380 938.330 58.440 ;
        RECT 1628.930 58.380 1629.250 58.440 ;
        RECT 938.010 58.240 1629.250 58.380 ;
        RECT 938.010 58.180 938.330 58.240 ;
        RECT 1628.930 58.180 1629.250 58.240 ;
      LAYER via ;
        RECT 938.040 58.180 938.300 58.440 ;
        RECT 1628.960 58.180 1629.220 58.440 ;
      LAYER met2 ;
        RECT 1630.260 1700.410 1630.540 1702.400 ;
        RECT 1629.020 1700.270 1630.540 1700.410 ;
        RECT 1629.020 58.470 1629.160 1700.270 ;
        RECT 1630.260 1700.000 1630.540 1700.270 ;
        RECT 938.040 58.150 938.300 58.470 ;
        RECT 1628.960 58.150 1629.220 58.470 ;
        RECT 938.100 17.410 938.240 58.150 ;
        RECT 936.260 17.270 938.240 17.410 ;
        RECT 936.260 2.400 936.400 17.270 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1636.365 1545.725 1636.535 1593.835 ;
        RECT 1636.365 1360.765 1636.535 1400.715 ;
        RECT 1636.365 1256.045 1636.535 1304.155 ;
        RECT 1635.905 662.405 1636.075 676.515 ;
        RECT 1635.905 524.365 1636.075 572.475 ;
        RECT 1636.365 427.805 1636.535 475.915 ;
        RECT 1635.905 331.245 1636.075 379.355 ;
      LAYER mcon ;
        RECT 1636.365 1593.665 1636.535 1593.835 ;
        RECT 1636.365 1400.545 1636.535 1400.715 ;
        RECT 1636.365 1303.985 1636.535 1304.155 ;
        RECT 1635.905 676.345 1636.075 676.515 ;
        RECT 1635.905 572.305 1636.075 572.475 ;
        RECT 1636.365 475.745 1636.535 475.915 ;
        RECT 1635.905 379.185 1636.075 379.355 ;
      LAYER met1 ;
        RECT 1636.290 1593.820 1636.610 1593.880 ;
        RECT 1636.095 1593.680 1636.610 1593.820 ;
        RECT 1636.290 1593.620 1636.610 1593.680 ;
        RECT 1636.290 1545.880 1636.610 1545.940 ;
        RECT 1636.095 1545.740 1636.610 1545.880 ;
        RECT 1636.290 1545.680 1636.610 1545.740 ;
        RECT 1636.290 1463.060 1636.610 1463.320 ;
        RECT 1636.380 1462.640 1636.520 1463.060 ;
        RECT 1636.290 1462.380 1636.610 1462.640 ;
        RECT 1636.290 1400.700 1636.610 1400.760 ;
        RECT 1636.095 1400.560 1636.610 1400.700 ;
        RECT 1636.290 1400.500 1636.610 1400.560 ;
        RECT 1636.290 1360.920 1636.610 1360.980 ;
        RECT 1636.095 1360.780 1636.610 1360.920 ;
        RECT 1636.290 1360.720 1636.610 1360.780 ;
        RECT 1636.290 1304.140 1636.610 1304.200 ;
        RECT 1636.095 1304.000 1636.610 1304.140 ;
        RECT 1636.290 1303.940 1636.610 1304.000 ;
        RECT 1636.290 1256.200 1636.610 1256.260 ;
        RECT 1636.095 1256.060 1636.610 1256.200 ;
        RECT 1636.290 1256.000 1636.610 1256.060 ;
        RECT 1636.750 1173.240 1637.070 1173.300 ;
        RECT 1636.380 1173.100 1637.070 1173.240 ;
        RECT 1636.380 1172.960 1636.520 1173.100 ;
        RECT 1636.750 1173.040 1637.070 1173.100 ;
        RECT 1636.290 1172.700 1636.610 1172.960 ;
        RECT 1636.750 1076.680 1637.070 1076.740 ;
        RECT 1636.380 1076.540 1637.070 1076.680 ;
        RECT 1636.380 1076.400 1636.520 1076.540 ;
        RECT 1636.750 1076.480 1637.070 1076.540 ;
        RECT 1636.290 1076.140 1636.610 1076.400 ;
        RECT 1636.750 966.320 1637.070 966.580 ;
        RECT 1636.840 965.900 1636.980 966.320 ;
        RECT 1636.750 965.640 1637.070 965.900 ;
        RECT 1635.830 940.680 1636.150 940.740 ;
        RECT 1636.750 940.680 1637.070 940.740 ;
        RECT 1635.830 940.540 1637.070 940.680 ;
        RECT 1635.830 940.480 1636.150 940.540 ;
        RECT 1636.750 940.480 1637.070 940.540 ;
        RECT 1635.830 883.360 1636.150 883.620 ;
        RECT 1635.920 882.880 1636.060 883.360 ;
        RECT 1636.290 882.880 1636.610 882.940 ;
        RECT 1635.920 882.740 1636.610 882.880 ;
        RECT 1636.290 882.680 1636.610 882.740 ;
        RECT 1636.290 738.380 1636.610 738.440 ;
        RECT 1635.920 738.240 1636.610 738.380 ;
        RECT 1635.920 738.100 1636.060 738.240 ;
        RECT 1636.290 738.180 1636.610 738.240 ;
        RECT 1635.830 737.840 1636.150 738.100 ;
        RECT 1635.830 676.500 1636.150 676.560 ;
        RECT 1635.635 676.360 1636.150 676.500 ;
        RECT 1635.830 676.300 1636.150 676.360 ;
        RECT 1635.830 662.560 1636.150 662.620 ;
        RECT 1635.635 662.420 1636.150 662.560 ;
        RECT 1635.830 662.360 1636.150 662.420 ;
        RECT 1635.830 572.460 1636.150 572.520 ;
        RECT 1635.635 572.320 1636.150 572.460 ;
        RECT 1635.830 572.260 1636.150 572.320 ;
        RECT 1635.845 524.520 1636.135 524.565 ;
        RECT 1636.290 524.520 1636.610 524.580 ;
        RECT 1635.845 524.380 1636.610 524.520 ;
        RECT 1635.845 524.335 1636.135 524.380 ;
        RECT 1636.290 524.320 1636.610 524.380 ;
        RECT 1636.290 497.460 1636.610 497.720 ;
        RECT 1636.380 496.700 1636.520 497.460 ;
        RECT 1636.290 496.440 1636.610 496.700 ;
        RECT 1636.290 475.900 1636.610 475.960 ;
        RECT 1636.095 475.760 1636.610 475.900 ;
        RECT 1636.290 475.700 1636.610 475.760 ;
        RECT 1636.290 427.960 1636.610 428.020 ;
        RECT 1636.095 427.820 1636.610 427.960 ;
        RECT 1636.290 427.760 1636.610 427.820 ;
        RECT 1636.290 386.820 1636.610 386.880 ;
        RECT 1635.920 386.680 1636.610 386.820 ;
        RECT 1635.920 386.200 1636.060 386.680 ;
        RECT 1636.290 386.620 1636.610 386.680 ;
        RECT 1635.830 385.940 1636.150 386.200 ;
        RECT 1635.830 379.340 1636.150 379.400 ;
        RECT 1635.635 379.200 1636.150 379.340 ;
        RECT 1635.830 379.140 1636.150 379.200 ;
        RECT 1635.845 331.400 1636.135 331.445 ;
        RECT 1636.290 331.400 1636.610 331.460 ;
        RECT 1635.845 331.260 1636.610 331.400 ;
        RECT 1635.845 331.215 1636.135 331.260 ;
        RECT 1636.290 331.200 1636.610 331.260 ;
        RECT 1636.290 241.980 1636.610 242.040 ;
        RECT 1635.920 241.840 1636.610 241.980 ;
        RECT 1635.920 241.700 1636.060 241.840 ;
        RECT 1636.290 241.780 1636.610 241.840 ;
        RECT 1635.830 241.440 1636.150 241.700 ;
        RECT 1635.830 138.280 1636.150 138.340 ;
        RECT 1636.290 138.280 1636.610 138.340 ;
        RECT 1635.830 138.140 1636.610 138.280 ;
        RECT 1635.830 138.080 1636.150 138.140 ;
        RECT 1636.290 138.080 1636.610 138.140 ;
        RECT 958.710 58.040 959.030 58.100 ;
        RECT 1636.290 58.040 1636.610 58.100 ;
        RECT 958.710 57.900 1636.610 58.040 ;
        RECT 958.710 57.840 959.030 57.900 ;
        RECT 1636.290 57.840 1636.610 57.900 ;
      LAYER via ;
        RECT 1636.320 1593.620 1636.580 1593.880 ;
        RECT 1636.320 1545.680 1636.580 1545.940 ;
        RECT 1636.320 1463.060 1636.580 1463.320 ;
        RECT 1636.320 1462.380 1636.580 1462.640 ;
        RECT 1636.320 1400.500 1636.580 1400.760 ;
        RECT 1636.320 1360.720 1636.580 1360.980 ;
        RECT 1636.320 1303.940 1636.580 1304.200 ;
        RECT 1636.320 1256.000 1636.580 1256.260 ;
        RECT 1636.780 1173.040 1637.040 1173.300 ;
        RECT 1636.320 1172.700 1636.580 1172.960 ;
        RECT 1636.780 1076.480 1637.040 1076.740 ;
        RECT 1636.320 1076.140 1636.580 1076.400 ;
        RECT 1636.780 966.320 1637.040 966.580 ;
        RECT 1636.780 965.640 1637.040 965.900 ;
        RECT 1635.860 940.480 1636.120 940.740 ;
        RECT 1636.780 940.480 1637.040 940.740 ;
        RECT 1635.860 883.360 1636.120 883.620 ;
        RECT 1636.320 882.680 1636.580 882.940 ;
        RECT 1636.320 738.180 1636.580 738.440 ;
        RECT 1635.860 737.840 1636.120 738.100 ;
        RECT 1635.860 676.300 1636.120 676.560 ;
        RECT 1635.860 662.360 1636.120 662.620 ;
        RECT 1635.860 572.260 1636.120 572.520 ;
        RECT 1636.320 524.320 1636.580 524.580 ;
        RECT 1636.320 497.460 1636.580 497.720 ;
        RECT 1636.320 496.440 1636.580 496.700 ;
        RECT 1636.320 475.700 1636.580 475.960 ;
        RECT 1636.320 427.760 1636.580 428.020 ;
        RECT 1636.320 386.620 1636.580 386.880 ;
        RECT 1635.860 385.940 1636.120 386.200 ;
        RECT 1635.860 379.140 1636.120 379.400 ;
        RECT 1636.320 331.200 1636.580 331.460 ;
        RECT 1636.320 241.780 1636.580 242.040 ;
        RECT 1635.860 241.440 1636.120 241.700 ;
        RECT 1635.860 138.080 1636.120 138.340 ;
        RECT 1636.320 138.080 1636.580 138.340 ;
        RECT 958.740 57.840 959.000 58.100 ;
        RECT 1636.320 57.840 1636.580 58.100 ;
      LAYER met2 ;
        RECT 1639.460 1700.410 1639.740 1702.400 ;
        RECT 1637.300 1700.270 1639.740 1700.410 ;
        RECT 1637.300 1643.405 1637.440 1700.270 ;
        RECT 1639.460 1700.000 1639.740 1700.270 ;
        RECT 1637.230 1643.035 1637.510 1643.405 ;
        RECT 1635.850 1642.355 1636.130 1642.725 ;
        RECT 1635.920 1606.570 1636.060 1642.355 ;
        RECT 1635.920 1606.430 1636.520 1606.570 ;
        RECT 1636.380 1593.910 1636.520 1606.430 ;
        RECT 1636.320 1593.590 1636.580 1593.910 ;
        RECT 1636.320 1545.650 1636.580 1545.970 ;
        RECT 1636.380 1463.350 1636.520 1545.650 ;
        RECT 1636.320 1463.030 1636.580 1463.350 ;
        RECT 1636.320 1462.350 1636.580 1462.670 ;
        RECT 1636.380 1400.790 1636.520 1462.350 ;
        RECT 1636.320 1400.470 1636.580 1400.790 ;
        RECT 1636.320 1360.690 1636.580 1361.010 ;
        RECT 1636.380 1304.230 1636.520 1360.690 ;
        RECT 1636.320 1303.910 1636.580 1304.230 ;
        RECT 1636.320 1255.970 1636.580 1256.290 ;
        RECT 1636.380 1207.410 1636.520 1255.970 ;
        RECT 1636.380 1207.270 1636.980 1207.410 ;
        RECT 1636.840 1173.330 1636.980 1207.270 ;
        RECT 1636.780 1173.010 1637.040 1173.330 ;
        RECT 1636.320 1172.670 1636.580 1172.990 ;
        RECT 1636.380 1110.850 1636.520 1172.670 ;
        RECT 1636.380 1110.710 1636.980 1110.850 ;
        RECT 1636.840 1076.770 1636.980 1110.710 ;
        RECT 1636.780 1076.450 1637.040 1076.770 ;
        RECT 1636.320 1076.110 1636.580 1076.430 ;
        RECT 1636.380 983.010 1636.520 1076.110 ;
        RECT 1636.380 982.870 1636.980 983.010 ;
        RECT 1636.840 966.610 1636.980 982.870 ;
        RECT 1636.780 966.290 1637.040 966.610 ;
        RECT 1636.780 965.610 1637.040 965.930 ;
        RECT 1636.840 940.770 1636.980 965.610 ;
        RECT 1635.860 940.450 1636.120 940.770 ;
        RECT 1636.780 940.450 1637.040 940.770 ;
        RECT 1635.920 883.650 1636.060 940.450 ;
        RECT 1635.860 883.330 1636.120 883.650 ;
        RECT 1636.320 882.650 1636.580 882.970 ;
        RECT 1636.380 787.170 1636.520 882.650 ;
        RECT 1635.920 787.030 1636.520 787.170 ;
        RECT 1635.920 786.490 1636.060 787.030 ;
        RECT 1635.920 786.350 1636.520 786.490 ;
        RECT 1636.380 738.470 1636.520 786.350 ;
        RECT 1636.320 738.150 1636.580 738.470 ;
        RECT 1635.860 737.810 1636.120 738.130 ;
        RECT 1635.920 676.590 1636.060 737.810 ;
        RECT 1635.860 676.270 1636.120 676.590 ;
        RECT 1635.860 662.330 1636.120 662.650 ;
        RECT 1635.920 621.365 1636.060 662.330 ;
        RECT 1635.850 620.995 1636.130 621.365 ;
        RECT 1635.850 619.635 1636.130 620.005 ;
        RECT 1635.920 572.550 1636.060 619.635 ;
        RECT 1635.860 572.230 1636.120 572.550 ;
        RECT 1636.320 524.290 1636.580 524.610 ;
        RECT 1636.380 497.750 1636.520 524.290 ;
        RECT 1636.320 497.430 1636.580 497.750 ;
        RECT 1636.320 496.410 1636.580 496.730 ;
        RECT 1636.380 475.990 1636.520 496.410 ;
        RECT 1636.320 475.670 1636.580 475.990 ;
        RECT 1636.320 427.730 1636.580 428.050 ;
        RECT 1636.380 386.910 1636.520 427.730 ;
        RECT 1636.320 386.590 1636.580 386.910 ;
        RECT 1635.860 385.910 1636.120 386.230 ;
        RECT 1635.920 379.430 1636.060 385.910 ;
        RECT 1635.860 379.110 1636.120 379.430 ;
        RECT 1636.320 331.170 1636.580 331.490 ;
        RECT 1636.380 242.070 1636.520 331.170 ;
        RECT 1636.320 241.750 1636.580 242.070 ;
        RECT 1635.860 241.410 1636.120 241.730 ;
        RECT 1635.920 138.370 1636.060 241.410 ;
        RECT 1635.860 138.050 1636.120 138.370 ;
        RECT 1636.320 138.050 1636.580 138.370 ;
        RECT 1636.380 58.130 1636.520 138.050 ;
        RECT 958.740 57.810 959.000 58.130 ;
        RECT 1636.320 57.810 1636.580 58.130 ;
        RECT 958.800 17.410 958.940 57.810 ;
        RECT 954.200 17.270 958.940 17.410 ;
        RECT 954.200 2.400 954.340 17.270 ;
        RECT 953.990 -4.800 954.550 2.400 ;
      LAYER via2 ;
        RECT 1637.230 1643.080 1637.510 1643.360 ;
        RECT 1635.850 1642.400 1636.130 1642.680 ;
        RECT 1635.850 621.040 1636.130 621.320 ;
        RECT 1635.850 619.680 1636.130 619.960 ;
      LAYER met3 ;
        RECT 1637.205 1643.370 1637.535 1643.385 ;
        RECT 1635.150 1643.070 1637.535 1643.370 ;
        RECT 1635.150 1642.690 1635.450 1643.070 ;
        RECT 1637.205 1643.055 1637.535 1643.070 ;
        RECT 1635.825 1642.690 1636.155 1642.705 ;
        RECT 1635.150 1642.390 1636.155 1642.690 ;
        RECT 1635.825 1642.375 1636.155 1642.390 ;
        RECT 1635.825 621.330 1636.155 621.345 ;
        RECT 1635.825 621.030 1637.290 621.330 ;
        RECT 1635.825 621.015 1636.155 621.030 ;
        RECT 1635.825 619.970 1636.155 619.985 ;
        RECT 1636.990 619.970 1637.290 621.030 ;
        RECT 1635.825 619.670 1637.290 619.970 ;
        RECT 1635.825 619.655 1636.155 619.670 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1643.190 1678.140 1643.510 1678.200 ;
        RECT 1646.870 1678.140 1647.190 1678.200 ;
        RECT 1643.190 1678.000 1647.190 1678.140 ;
        RECT 1643.190 1677.940 1643.510 1678.000 ;
        RECT 1646.870 1677.940 1647.190 1678.000 ;
        RECT 972.510 57.700 972.830 57.760 ;
        RECT 1643.190 57.700 1643.510 57.760 ;
        RECT 972.510 57.560 1643.510 57.700 ;
        RECT 972.510 57.500 972.830 57.560 ;
        RECT 1643.190 57.500 1643.510 57.560 ;
      LAYER via ;
        RECT 1643.220 1677.940 1643.480 1678.200 ;
        RECT 1646.900 1677.940 1647.160 1678.200 ;
        RECT 972.540 57.500 972.800 57.760 ;
        RECT 1643.220 57.500 1643.480 57.760 ;
      LAYER met2 ;
        RECT 1648.660 1700.410 1648.940 1702.400 ;
        RECT 1646.960 1700.270 1648.940 1700.410 ;
        RECT 1646.960 1678.230 1647.100 1700.270 ;
        RECT 1648.660 1700.000 1648.940 1700.270 ;
        RECT 1643.220 1677.910 1643.480 1678.230 ;
        RECT 1646.900 1677.910 1647.160 1678.230 ;
        RECT 1643.280 57.790 1643.420 1677.910 ;
        RECT 972.540 57.470 972.800 57.790 ;
        RECT 1643.220 57.470 1643.480 57.790 ;
        RECT 972.600 17.410 972.740 57.470 ;
        RECT 972.140 17.270 972.740 17.410 ;
        RECT 972.140 2.400 972.280 17.270 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 26.760 651.290 26.820 ;
        RECT 1483.570 26.760 1483.890 26.820 ;
        RECT 650.970 26.620 1483.890 26.760 ;
        RECT 650.970 26.560 651.290 26.620 ;
        RECT 1483.570 26.560 1483.890 26.620 ;
      LAYER via ;
        RECT 651.000 26.560 651.260 26.820 ;
        RECT 1483.600 26.560 1483.860 26.820 ;
      LAYER met2 ;
        RECT 1483.520 1700.000 1483.800 1702.400 ;
        RECT 1483.660 26.850 1483.800 1700.000 ;
        RECT 651.000 26.530 651.260 26.850 ;
        RECT 1483.600 26.530 1483.860 26.850 ;
        RECT 651.060 2.400 651.200 26.530 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1656.070 966.320 1656.390 966.580 ;
        RECT 1656.160 965.900 1656.300 966.320 ;
        RECT 1656.070 965.640 1656.390 965.900 ;
        RECT 993.210 57.360 993.530 57.420 ;
        RECT 1656.070 57.360 1656.390 57.420 ;
        RECT 993.210 57.220 1656.390 57.360 ;
        RECT 993.210 57.160 993.530 57.220 ;
        RECT 1656.070 57.160 1656.390 57.220 ;
      LAYER via ;
        RECT 1656.100 966.320 1656.360 966.580 ;
        RECT 1656.100 965.640 1656.360 965.900 ;
        RECT 993.240 57.160 993.500 57.420 ;
        RECT 1656.100 57.160 1656.360 57.420 ;
      LAYER met2 ;
        RECT 1657.860 1700.410 1658.140 1702.400 ;
        RECT 1656.160 1700.270 1658.140 1700.410 ;
        RECT 1656.160 966.610 1656.300 1700.270 ;
        RECT 1657.860 1700.000 1658.140 1700.270 ;
        RECT 1656.100 966.290 1656.360 966.610 ;
        RECT 1656.100 965.610 1656.360 965.930 ;
        RECT 1656.160 57.450 1656.300 965.610 ;
        RECT 993.240 57.130 993.500 57.450 ;
        RECT 1656.100 57.130 1656.360 57.450 ;
        RECT 993.300 17.410 993.440 57.130 ;
        RECT 990.080 17.270 993.440 17.410 ;
        RECT 990.080 2.400 990.220 17.270 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1663.965 1545.725 1664.135 1593.835 ;
        RECT 1664.425 275.825 1664.595 317.475 ;
        RECT 1663.505 179.605 1663.675 227.715 ;
      LAYER mcon ;
        RECT 1663.965 1593.665 1664.135 1593.835 ;
        RECT 1664.425 317.305 1664.595 317.475 ;
        RECT 1663.505 227.545 1663.675 227.715 ;
      LAYER met1 ;
        RECT 1663.430 1642.440 1663.750 1642.500 ;
        RECT 1664.810 1642.440 1665.130 1642.500 ;
        RECT 1663.430 1642.300 1665.130 1642.440 ;
        RECT 1663.430 1642.240 1663.750 1642.300 ;
        RECT 1664.810 1642.240 1665.130 1642.300 ;
        RECT 1663.890 1593.820 1664.210 1593.880 ;
        RECT 1663.695 1593.680 1664.210 1593.820 ;
        RECT 1663.890 1593.620 1664.210 1593.680 ;
        RECT 1663.890 1545.880 1664.210 1545.940 ;
        RECT 1663.695 1545.740 1664.210 1545.880 ;
        RECT 1663.890 1545.680 1664.210 1545.740 ;
        RECT 1663.890 1463.060 1664.210 1463.320 ;
        RECT 1663.980 1462.640 1664.120 1463.060 ;
        RECT 1663.890 1462.380 1664.210 1462.640 ;
        RECT 1663.890 1366.500 1664.210 1366.760 ;
        RECT 1663.980 1366.080 1664.120 1366.500 ;
        RECT 1663.890 1365.820 1664.210 1366.080 ;
        RECT 1663.890 324.260 1664.210 324.320 ;
        RECT 1664.350 324.260 1664.670 324.320 ;
        RECT 1663.890 324.120 1664.670 324.260 ;
        RECT 1663.890 324.060 1664.210 324.120 ;
        RECT 1664.350 324.060 1664.670 324.120 ;
        RECT 1664.350 317.460 1664.670 317.520 ;
        RECT 1664.155 317.320 1664.670 317.460 ;
        RECT 1664.350 317.260 1664.670 317.320 ;
        RECT 1664.350 275.980 1664.670 276.040 ;
        RECT 1664.155 275.840 1664.670 275.980 ;
        RECT 1664.350 275.780 1664.670 275.840 ;
        RECT 1664.350 234.640 1664.670 234.900 ;
        RECT 1664.440 234.220 1664.580 234.640 ;
        RECT 1664.350 233.960 1664.670 234.220 ;
        RECT 1663.445 227.700 1663.735 227.745 ;
        RECT 1664.350 227.700 1664.670 227.760 ;
        RECT 1663.445 227.560 1664.670 227.700 ;
        RECT 1663.445 227.515 1663.735 227.560 ;
        RECT 1664.350 227.500 1664.670 227.560 ;
        RECT 1663.430 179.760 1663.750 179.820 ;
        RECT 1663.235 179.620 1663.750 179.760 ;
        RECT 1663.430 179.560 1663.750 179.620 ;
        RECT 1007.470 57.020 1007.790 57.080 ;
        RECT 1663.890 57.020 1664.210 57.080 ;
        RECT 1007.470 56.880 1664.210 57.020 ;
        RECT 1007.470 56.820 1007.790 56.880 ;
        RECT 1663.890 56.820 1664.210 56.880 ;
      LAYER via ;
        RECT 1663.460 1642.240 1663.720 1642.500 ;
        RECT 1664.840 1642.240 1665.100 1642.500 ;
        RECT 1663.920 1593.620 1664.180 1593.880 ;
        RECT 1663.920 1545.680 1664.180 1545.940 ;
        RECT 1663.920 1463.060 1664.180 1463.320 ;
        RECT 1663.920 1462.380 1664.180 1462.640 ;
        RECT 1663.920 1366.500 1664.180 1366.760 ;
        RECT 1663.920 1365.820 1664.180 1366.080 ;
        RECT 1663.920 324.060 1664.180 324.320 ;
        RECT 1664.380 324.060 1664.640 324.320 ;
        RECT 1664.380 317.260 1664.640 317.520 ;
        RECT 1664.380 275.780 1664.640 276.040 ;
        RECT 1664.380 234.640 1664.640 234.900 ;
        RECT 1664.380 233.960 1664.640 234.220 ;
        RECT 1664.380 227.500 1664.640 227.760 ;
        RECT 1663.460 179.560 1663.720 179.820 ;
        RECT 1007.500 56.820 1007.760 57.080 ;
        RECT 1663.920 56.820 1664.180 57.080 ;
      LAYER met2 ;
        RECT 1667.060 1700.410 1667.340 1702.400 ;
        RECT 1665.820 1700.270 1667.340 1700.410 ;
        RECT 1665.820 1690.380 1665.960 1700.270 ;
        RECT 1667.060 1700.000 1667.340 1700.270 ;
        RECT 1664.900 1690.240 1665.960 1690.380 ;
        RECT 1664.900 1642.530 1665.040 1690.240 ;
        RECT 1663.460 1642.210 1663.720 1642.530 ;
        RECT 1664.840 1642.210 1665.100 1642.530 ;
        RECT 1663.520 1642.045 1663.660 1642.210 ;
        RECT 1663.450 1641.675 1663.730 1642.045 ;
        RECT 1663.910 1594.075 1664.190 1594.445 ;
        RECT 1663.980 1593.910 1664.120 1594.075 ;
        RECT 1663.920 1593.590 1664.180 1593.910 ;
        RECT 1663.920 1545.650 1664.180 1545.970 ;
        RECT 1663.980 1463.350 1664.120 1545.650 ;
        RECT 1663.920 1463.030 1664.180 1463.350 ;
        RECT 1663.920 1462.350 1664.180 1462.670 ;
        RECT 1663.980 1366.790 1664.120 1462.350 ;
        RECT 1663.920 1366.470 1664.180 1366.790 ;
        RECT 1663.920 1365.790 1664.180 1366.110 ;
        RECT 1663.980 787.170 1664.120 1365.790 ;
        RECT 1663.520 787.030 1664.120 787.170 ;
        RECT 1663.520 786.490 1663.660 787.030 ;
        RECT 1663.520 786.350 1664.120 786.490 ;
        RECT 1663.980 594.050 1664.120 786.350 ;
        RECT 1663.520 593.910 1664.120 594.050 ;
        RECT 1663.520 593.370 1663.660 593.910 ;
        RECT 1663.520 593.230 1664.120 593.370 ;
        RECT 1663.980 324.350 1664.120 593.230 ;
        RECT 1663.920 324.030 1664.180 324.350 ;
        RECT 1664.380 324.030 1664.640 324.350 ;
        RECT 1664.440 317.550 1664.580 324.030 ;
        RECT 1664.380 317.230 1664.640 317.550 ;
        RECT 1664.380 275.750 1664.640 276.070 ;
        RECT 1664.440 234.930 1664.580 275.750 ;
        RECT 1664.380 234.610 1664.640 234.930 ;
        RECT 1664.380 233.930 1664.640 234.250 ;
        RECT 1664.440 227.790 1664.580 233.930 ;
        RECT 1664.380 227.470 1664.640 227.790 ;
        RECT 1663.460 179.530 1663.720 179.850 ;
        RECT 1663.520 150.690 1663.660 179.530 ;
        RECT 1663.520 150.550 1664.120 150.690 ;
        RECT 1663.980 57.110 1664.120 150.550 ;
        RECT 1007.500 56.790 1007.760 57.110 ;
        RECT 1663.920 56.790 1664.180 57.110 ;
        RECT 1007.560 2.400 1007.700 56.790 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
      LAYER via2 ;
        RECT 1663.450 1641.720 1663.730 1642.000 ;
        RECT 1663.910 1594.120 1664.190 1594.400 ;
      LAYER met3 ;
        RECT 1663.425 1642.020 1663.755 1642.025 ;
        RECT 1663.425 1642.010 1664.010 1642.020 ;
        RECT 1663.200 1641.710 1664.010 1642.010 ;
        RECT 1663.425 1641.700 1664.010 1641.710 ;
        RECT 1663.425 1641.695 1663.755 1641.700 ;
        RECT 1663.630 1595.090 1664.010 1595.100 ;
        RECT 1663.630 1594.790 1664.890 1595.090 ;
        RECT 1663.630 1594.780 1664.010 1594.790 ;
        RECT 1663.885 1594.410 1664.215 1594.425 ;
        RECT 1664.590 1594.410 1664.890 1594.790 ;
        RECT 1663.885 1594.110 1664.890 1594.410 ;
        RECT 1663.885 1594.095 1664.215 1594.110 ;
      LAYER via3 ;
        RECT 1663.660 1641.700 1663.980 1642.020 ;
        RECT 1663.660 1594.780 1663.980 1595.100 ;
      LAYER met4 ;
        RECT 1663.655 1641.695 1663.985 1642.025 ;
        RECT 1663.670 1595.105 1663.970 1641.695 ;
        RECT 1663.655 1594.775 1663.985 1595.105 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1672.245 1538.925 1672.415 1545.895 ;
        RECT 1671.325 1413.805 1671.495 1490.475 ;
        RECT 1671.785 1352.945 1671.955 1400.715 ;
        RECT 1671.785 1256.385 1671.955 1304.155 ;
        RECT 1671.785 1220.685 1671.955 1255.875 ;
        RECT 1672.245 917.745 1672.415 932.195 ;
        RECT 1671.785 848.725 1671.955 879.495 ;
        RECT 1671.785 675.665 1671.955 724.455 ;
        RECT 1671.785 565.845 1671.955 572.815 ;
        RECT 1671.785 469.285 1671.955 517.395 ;
        RECT 1671.785 386.325 1671.955 434.435 ;
        RECT 1671.785 241.485 1671.955 278.375 ;
        RECT 1671.785 131.325 1671.955 179.435 ;
      LAYER mcon ;
        RECT 1672.245 1545.725 1672.415 1545.895 ;
        RECT 1671.325 1490.305 1671.495 1490.475 ;
        RECT 1671.785 1400.545 1671.955 1400.715 ;
        RECT 1671.785 1303.985 1671.955 1304.155 ;
        RECT 1671.785 1255.705 1671.955 1255.875 ;
        RECT 1672.245 932.025 1672.415 932.195 ;
        RECT 1671.785 879.325 1671.955 879.495 ;
        RECT 1671.785 724.285 1671.955 724.455 ;
        RECT 1671.785 572.645 1671.955 572.815 ;
        RECT 1671.785 517.225 1671.955 517.395 ;
        RECT 1671.785 434.265 1671.955 434.435 ;
        RECT 1671.785 278.205 1671.955 278.375 ;
        RECT 1671.785 179.265 1671.955 179.435 ;
      LAYER met1 ;
        RECT 1672.170 1642.440 1672.490 1642.500 ;
        RECT 1674.010 1642.440 1674.330 1642.500 ;
        RECT 1672.170 1642.300 1674.330 1642.440 ;
        RECT 1672.170 1642.240 1672.490 1642.300 ;
        RECT 1674.010 1642.240 1674.330 1642.300 ;
        RECT 1672.170 1545.880 1672.490 1545.940 ;
        RECT 1671.975 1545.740 1672.490 1545.880 ;
        RECT 1672.170 1545.680 1672.490 1545.740 ;
        RECT 1672.170 1539.080 1672.490 1539.140 ;
        RECT 1671.975 1538.940 1672.490 1539.080 ;
        RECT 1672.170 1538.880 1672.490 1538.940 ;
        RECT 1671.250 1497.260 1671.570 1497.320 ;
        RECT 1672.170 1497.260 1672.490 1497.320 ;
        RECT 1671.250 1497.120 1672.490 1497.260 ;
        RECT 1671.250 1497.060 1671.570 1497.120 ;
        RECT 1672.170 1497.060 1672.490 1497.120 ;
        RECT 1671.250 1490.460 1671.570 1490.520 ;
        RECT 1671.055 1490.320 1671.570 1490.460 ;
        RECT 1671.250 1490.260 1671.570 1490.320 ;
        RECT 1671.265 1413.960 1671.555 1414.005 ;
        RECT 1672.170 1413.960 1672.490 1414.020 ;
        RECT 1671.265 1413.820 1672.490 1413.960 ;
        RECT 1671.265 1413.775 1671.555 1413.820 ;
        RECT 1672.170 1413.760 1672.490 1413.820 ;
        RECT 1671.725 1400.700 1672.015 1400.745 ;
        RECT 1672.170 1400.700 1672.490 1400.760 ;
        RECT 1671.725 1400.560 1672.490 1400.700 ;
        RECT 1671.725 1400.515 1672.015 1400.560 ;
        RECT 1672.170 1400.500 1672.490 1400.560 ;
        RECT 1671.710 1353.100 1672.030 1353.160 ;
        RECT 1671.515 1352.960 1672.030 1353.100 ;
        RECT 1671.710 1352.900 1672.030 1352.960 ;
        RECT 1671.710 1317.880 1672.030 1318.140 ;
        RECT 1671.800 1317.400 1671.940 1317.880 ;
        RECT 1672.170 1317.400 1672.490 1317.460 ;
        RECT 1671.800 1317.260 1672.490 1317.400 ;
        RECT 1672.170 1317.200 1672.490 1317.260 ;
        RECT 1671.725 1304.140 1672.015 1304.185 ;
        RECT 1672.170 1304.140 1672.490 1304.200 ;
        RECT 1671.725 1304.000 1672.490 1304.140 ;
        RECT 1671.725 1303.955 1672.015 1304.000 ;
        RECT 1672.170 1303.940 1672.490 1304.000 ;
        RECT 1671.710 1256.540 1672.030 1256.600 ;
        RECT 1671.515 1256.400 1672.030 1256.540 ;
        RECT 1671.710 1256.340 1672.030 1256.400 ;
        RECT 1671.710 1255.860 1672.030 1255.920 ;
        RECT 1671.515 1255.720 1672.030 1255.860 ;
        RECT 1671.710 1255.660 1672.030 1255.720 ;
        RECT 1671.710 1220.840 1672.030 1220.900 ;
        RECT 1671.515 1220.700 1672.030 1220.840 ;
        RECT 1671.710 1220.640 1672.030 1220.700 ;
        RECT 1671.710 1159.980 1672.030 1160.040 ;
        RECT 1671.710 1159.840 1672.400 1159.980 ;
        RECT 1671.710 1159.780 1672.030 1159.840 ;
        RECT 1672.260 1159.360 1672.400 1159.840 ;
        RECT 1672.170 1159.100 1672.490 1159.360 ;
        RECT 1671.710 1063.420 1672.030 1063.480 ;
        RECT 1671.710 1063.280 1672.400 1063.420 ;
        RECT 1671.710 1063.220 1672.030 1063.280 ;
        RECT 1672.260 1062.800 1672.400 1063.280 ;
        RECT 1672.170 1062.540 1672.490 1062.800 ;
        RECT 1671.710 966.860 1672.030 966.920 ;
        RECT 1671.710 966.720 1672.400 966.860 ;
        RECT 1671.710 966.660 1672.030 966.720 ;
        RECT 1672.260 966.240 1672.400 966.720 ;
        RECT 1672.170 965.980 1672.490 966.240 ;
        RECT 1672.170 932.180 1672.490 932.240 ;
        RECT 1671.975 932.040 1672.490 932.180 ;
        RECT 1672.170 931.980 1672.490 932.040 ;
        RECT 1672.170 917.900 1672.490 917.960 ;
        RECT 1671.975 917.760 1672.490 917.900 ;
        RECT 1672.170 917.700 1672.490 917.760 ;
        RECT 1671.710 879.480 1672.030 879.540 ;
        RECT 1671.515 879.340 1672.030 879.480 ;
        RECT 1671.710 879.280 1672.030 879.340 ;
        RECT 1671.725 848.880 1672.015 848.925 ;
        RECT 1672.630 848.880 1672.950 848.940 ;
        RECT 1671.725 848.740 1672.950 848.880 ;
        RECT 1671.725 848.695 1672.015 848.740 ;
        RECT 1672.630 848.680 1672.950 848.740 ;
        RECT 1671.710 807.400 1672.030 807.460 ;
        RECT 1672.630 807.400 1672.950 807.460 ;
        RECT 1671.710 807.260 1672.950 807.400 ;
        RECT 1671.710 807.200 1672.030 807.260 ;
        RECT 1672.630 807.200 1672.950 807.260 ;
        RECT 1671.710 738.520 1672.030 738.780 ;
        RECT 1671.800 738.100 1671.940 738.520 ;
        RECT 1671.710 737.840 1672.030 738.100 ;
        RECT 1671.725 724.440 1672.015 724.485 ;
        RECT 1672.170 724.440 1672.490 724.500 ;
        RECT 1671.725 724.300 1672.490 724.440 ;
        RECT 1671.725 724.255 1672.015 724.300 ;
        RECT 1672.170 724.240 1672.490 724.300 ;
        RECT 1671.725 675.820 1672.015 675.865 ;
        RECT 1672.170 675.820 1672.490 675.880 ;
        RECT 1671.725 675.680 1672.490 675.820 ;
        RECT 1671.725 675.635 1672.015 675.680 ;
        RECT 1672.170 675.620 1672.490 675.680 ;
        RECT 1671.725 572.800 1672.015 572.845 ;
        RECT 1672.170 572.800 1672.490 572.860 ;
        RECT 1671.725 572.660 1672.490 572.800 ;
        RECT 1671.725 572.615 1672.015 572.660 ;
        RECT 1672.170 572.600 1672.490 572.660 ;
        RECT 1671.710 566.000 1672.030 566.060 ;
        RECT 1671.515 565.860 1672.030 566.000 ;
        RECT 1671.710 565.800 1672.030 565.860 ;
        RECT 1671.710 524.520 1672.030 524.580 ;
        RECT 1672.170 524.520 1672.490 524.580 ;
        RECT 1671.710 524.380 1672.490 524.520 ;
        RECT 1671.710 524.320 1672.030 524.380 ;
        RECT 1672.170 524.320 1672.490 524.380 ;
        RECT 1671.725 517.380 1672.015 517.425 ;
        RECT 1672.170 517.380 1672.490 517.440 ;
        RECT 1671.725 517.240 1672.490 517.380 ;
        RECT 1671.725 517.195 1672.015 517.240 ;
        RECT 1672.170 517.180 1672.490 517.240 ;
        RECT 1671.710 469.440 1672.030 469.500 ;
        RECT 1671.515 469.300 1672.030 469.440 ;
        RECT 1671.710 469.240 1672.030 469.300 ;
        RECT 1671.710 434.420 1672.030 434.480 ;
        RECT 1671.515 434.280 1672.030 434.420 ;
        RECT 1671.710 434.220 1672.030 434.280 ;
        RECT 1671.710 386.480 1672.030 386.540 ;
        RECT 1671.515 386.340 1672.030 386.480 ;
        RECT 1671.710 386.280 1672.030 386.340 ;
        RECT 1671.710 278.360 1672.030 278.420 ;
        RECT 1671.515 278.220 1672.030 278.360 ;
        RECT 1671.710 278.160 1672.030 278.220 ;
        RECT 1671.725 241.640 1672.015 241.685 ;
        RECT 1672.170 241.640 1672.490 241.700 ;
        RECT 1671.725 241.500 1672.490 241.640 ;
        RECT 1671.725 241.455 1672.015 241.500 ;
        RECT 1672.170 241.440 1672.490 241.500 ;
        RECT 1672.170 186.900 1672.490 186.960 ;
        RECT 1671.800 186.760 1672.490 186.900 ;
        RECT 1671.800 186.620 1671.940 186.760 ;
        RECT 1672.170 186.700 1672.490 186.760 ;
        RECT 1671.710 186.360 1672.030 186.620 ;
        RECT 1671.710 179.420 1672.030 179.480 ;
        RECT 1671.515 179.280 1672.030 179.420 ;
        RECT 1671.710 179.220 1672.030 179.280 ;
        RECT 1671.725 131.480 1672.015 131.525 ;
        RECT 1672.630 131.480 1672.950 131.540 ;
        RECT 1671.725 131.340 1672.950 131.480 ;
        RECT 1671.725 131.295 1672.015 131.340 ;
        RECT 1672.630 131.280 1672.950 131.340 ;
        RECT 1671.710 130.800 1672.030 130.860 ;
        RECT 1672.630 130.800 1672.950 130.860 ;
        RECT 1671.710 130.660 1672.950 130.800 ;
        RECT 1671.710 130.600 1672.030 130.660 ;
        RECT 1672.630 130.600 1672.950 130.660 ;
        RECT 1027.710 56.680 1028.030 56.740 ;
        RECT 1672.170 56.680 1672.490 56.740 ;
        RECT 1027.710 56.540 1672.490 56.680 ;
        RECT 1027.710 56.480 1028.030 56.540 ;
        RECT 1672.170 56.480 1672.490 56.540 ;
        RECT 1025.410 2.960 1025.730 3.020 ;
        RECT 1027.710 2.960 1028.030 3.020 ;
        RECT 1025.410 2.820 1028.030 2.960 ;
        RECT 1025.410 2.760 1025.730 2.820 ;
        RECT 1027.710 2.760 1028.030 2.820 ;
      LAYER via ;
        RECT 1672.200 1642.240 1672.460 1642.500 ;
        RECT 1674.040 1642.240 1674.300 1642.500 ;
        RECT 1672.200 1545.680 1672.460 1545.940 ;
        RECT 1672.200 1538.880 1672.460 1539.140 ;
        RECT 1671.280 1497.060 1671.540 1497.320 ;
        RECT 1672.200 1497.060 1672.460 1497.320 ;
        RECT 1671.280 1490.260 1671.540 1490.520 ;
        RECT 1672.200 1413.760 1672.460 1414.020 ;
        RECT 1672.200 1400.500 1672.460 1400.760 ;
        RECT 1671.740 1352.900 1672.000 1353.160 ;
        RECT 1671.740 1317.880 1672.000 1318.140 ;
        RECT 1672.200 1317.200 1672.460 1317.460 ;
        RECT 1672.200 1303.940 1672.460 1304.200 ;
        RECT 1671.740 1256.340 1672.000 1256.600 ;
        RECT 1671.740 1255.660 1672.000 1255.920 ;
        RECT 1671.740 1220.640 1672.000 1220.900 ;
        RECT 1671.740 1159.780 1672.000 1160.040 ;
        RECT 1672.200 1159.100 1672.460 1159.360 ;
        RECT 1671.740 1063.220 1672.000 1063.480 ;
        RECT 1672.200 1062.540 1672.460 1062.800 ;
        RECT 1671.740 966.660 1672.000 966.920 ;
        RECT 1672.200 965.980 1672.460 966.240 ;
        RECT 1672.200 931.980 1672.460 932.240 ;
        RECT 1672.200 917.700 1672.460 917.960 ;
        RECT 1671.740 879.280 1672.000 879.540 ;
        RECT 1672.660 848.680 1672.920 848.940 ;
        RECT 1671.740 807.200 1672.000 807.460 ;
        RECT 1672.660 807.200 1672.920 807.460 ;
        RECT 1671.740 738.520 1672.000 738.780 ;
        RECT 1671.740 737.840 1672.000 738.100 ;
        RECT 1672.200 724.240 1672.460 724.500 ;
        RECT 1672.200 675.620 1672.460 675.880 ;
        RECT 1672.200 572.600 1672.460 572.860 ;
        RECT 1671.740 565.800 1672.000 566.060 ;
        RECT 1671.740 524.320 1672.000 524.580 ;
        RECT 1672.200 524.320 1672.460 524.580 ;
        RECT 1672.200 517.180 1672.460 517.440 ;
        RECT 1671.740 469.240 1672.000 469.500 ;
        RECT 1671.740 434.220 1672.000 434.480 ;
        RECT 1671.740 386.280 1672.000 386.540 ;
        RECT 1671.740 278.160 1672.000 278.420 ;
        RECT 1672.200 241.440 1672.460 241.700 ;
        RECT 1672.200 186.700 1672.460 186.960 ;
        RECT 1671.740 186.360 1672.000 186.620 ;
        RECT 1671.740 179.220 1672.000 179.480 ;
        RECT 1672.660 131.280 1672.920 131.540 ;
        RECT 1671.740 130.600 1672.000 130.860 ;
        RECT 1672.660 130.600 1672.920 130.860 ;
        RECT 1027.740 56.480 1028.000 56.740 ;
        RECT 1672.200 56.480 1672.460 56.740 ;
        RECT 1025.440 2.760 1025.700 3.020 ;
        RECT 1027.740 2.760 1028.000 3.020 ;
      LAYER met2 ;
        RECT 1676.260 1701.090 1676.540 1702.400 ;
        RECT 1674.100 1700.950 1676.540 1701.090 ;
        RECT 1674.100 1642.530 1674.240 1700.950 ;
        RECT 1676.260 1700.000 1676.540 1700.950 ;
        RECT 1672.200 1642.210 1672.460 1642.530 ;
        RECT 1674.040 1642.210 1674.300 1642.530 ;
        RECT 1672.260 1545.970 1672.400 1642.210 ;
        RECT 1672.200 1545.650 1672.460 1545.970 ;
        RECT 1672.200 1538.850 1672.460 1539.170 ;
        RECT 1672.260 1497.350 1672.400 1538.850 ;
        RECT 1671.280 1497.030 1671.540 1497.350 ;
        RECT 1672.200 1497.030 1672.460 1497.350 ;
        RECT 1671.340 1490.550 1671.480 1497.030 ;
        RECT 1671.280 1490.230 1671.540 1490.550 ;
        RECT 1672.200 1413.730 1672.460 1414.050 ;
        RECT 1672.260 1400.790 1672.400 1413.730 ;
        RECT 1672.200 1400.470 1672.460 1400.790 ;
        RECT 1671.740 1352.870 1672.000 1353.190 ;
        RECT 1671.800 1318.170 1671.940 1352.870 ;
        RECT 1671.740 1317.850 1672.000 1318.170 ;
        RECT 1672.200 1317.170 1672.460 1317.490 ;
        RECT 1672.260 1304.230 1672.400 1317.170 ;
        RECT 1672.200 1303.910 1672.460 1304.230 ;
        RECT 1671.740 1256.310 1672.000 1256.630 ;
        RECT 1671.800 1255.950 1671.940 1256.310 ;
        RECT 1671.740 1255.630 1672.000 1255.950 ;
        RECT 1671.740 1220.610 1672.000 1220.930 ;
        RECT 1671.800 1160.070 1671.940 1220.610 ;
        RECT 1671.740 1159.750 1672.000 1160.070 ;
        RECT 1672.200 1159.070 1672.460 1159.390 ;
        RECT 1672.260 1134.650 1672.400 1159.070 ;
        RECT 1671.800 1134.510 1672.400 1134.650 ;
        RECT 1671.800 1063.510 1671.940 1134.510 ;
        RECT 1671.740 1063.190 1672.000 1063.510 ;
        RECT 1672.200 1062.510 1672.460 1062.830 ;
        RECT 1672.260 1038.090 1672.400 1062.510 ;
        RECT 1671.800 1037.950 1672.400 1038.090 ;
        RECT 1671.800 966.950 1671.940 1037.950 ;
        RECT 1671.740 966.630 1672.000 966.950 ;
        RECT 1672.200 965.950 1672.460 966.270 ;
        RECT 1672.260 932.270 1672.400 965.950 ;
        RECT 1672.200 931.950 1672.460 932.270 ;
        RECT 1672.260 917.990 1672.400 918.145 ;
        RECT 1672.200 917.730 1672.460 917.990 ;
        RECT 1671.800 917.670 1672.460 917.730 ;
        RECT 1671.800 917.590 1672.400 917.670 ;
        RECT 1671.800 879.570 1671.940 917.590 ;
        RECT 1671.740 879.250 1672.000 879.570 ;
        RECT 1672.660 848.650 1672.920 848.970 ;
        RECT 1672.720 807.490 1672.860 848.650 ;
        RECT 1671.740 807.170 1672.000 807.490 ;
        RECT 1672.660 807.170 1672.920 807.490 ;
        RECT 1671.800 806.890 1671.940 807.170 ;
        RECT 1671.340 806.750 1671.940 806.890 ;
        RECT 1671.340 787.170 1671.480 806.750 ;
        RECT 1671.340 787.030 1672.400 787.170 ;
        RECT 1672.260 783.770 1672.400 787.030 ;
        RECT 1671.800 783.630 1672.400 783.770 ;
        RECT 1671.800 738.810 1671.940 783.630 ;
        RECT 1671.740 738.490 1672.000 738.810 ;
        RECT 1671.740 737.810 1672.000 738.130 ;
        RECT 1671.800 724.610 1671.940 737.810 ;
        RECT 1671.800 724.530 1672.400 724.610 ;
        RECT 1671.800 724.470 1672.460 724.530 ;
        RECT 1672.200 724.210 1672.460 724.470 ;
        RECT 1672.200 675.590 1672.460 675.910 ;
        RECT 1672.260 572.890 1672.400 675.590 ;
        RECT 1672.200 572.570 1672.460 572.890 ;
        RECT 1671.740 565.770 1672.000 566.090 ;
        RECT 1671.800 524.610 1671.940 565.770 ;
        RECT 1671.740 524.290 1672.000 524.610 ;
        RECT 1672.200 524.290 1672.460 524.610 ;
        RECT 1672.260 517.470 1672.400 524.290 ;
        RECT 1672.200 517.150 1672.460 517.470 ;
        RECT 1671.740 469.210 1672.000 469.530 ;
        RECT 1671.800 434.510 1671.940 469.210 ;
        RECT 1671.740 434.190 1672.000 434.510 ;
        RECT 1671.740 386.250 1672.000 386.570 ;
        RECT 1671.800 278.450 1671.940 386.250 ;
        RECT 1671.740 278.130 1672.000 278.450 ;
        RECT 1672.200 241.410 1672.460 241.730 ;
        RECT 1672.260 186.990 1672.400 241.410 ;
        RECT 1672.200 186.670 1672.460 186.990 ;
        RECT 1671.740 186.330 1672.000 186.650 ;
        RECT 1671.800 179.510 1671.940 186.330 ;
        RECT 1671.740 179.190 1672.000 179.510 ;
        RECT 1672.660 131.250 1672.920 131.570 ;
        RECT 1672.720 130.890 1672.860 131.250 ;
        RECT 1671.740 130.570 1672.000 130.890 ;
        RECT 1672.660 130.570 1672.920 130.890 ;
        RECT 1671.800 106.490 1671.940 130.570 ;
        RECT 1671.800 106.350 1672.400 106.490 ;
        RECT 1672.260 56.770 1672.400 106.350 ;
        RECT 1027.740 56.450 1028.000 56.770 ;
        RECT 1672.200 56.450 1672.460 56.770 ;
        RECT 1027.800 3.050 1027.940 56.450 ;
        RECT 1025.440 2.730 1025.700 3.050 ;
        RECT 1027.740 2.730 1028.000 3.050 ;
        RECT 1025.500 2.400 1025.640 2.730 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1418.250 1686.300 1418.570 1686.360 ;
        RECT 1685.510 1686.300 1685.830 1686.360 ;
        RECT 1418.250 1686.160 1685.830 1686.300 ;
        RECT 1418.250 1686.100 1418.570 1686.160 ;
        RECT 1685.510 1686.100 1685.830 1686.160 ;
        RECT 1043.350 22.680 1043.670 22.740 ;
        RECT 1417.790 22.680 1418.110 22.740 ;
        RECT 1043.350 22.540 1418.110 22.680 ;
        RECT 1043.350 22.480 1043.670 22.540 ;
        RECT 1417.790 22.480 1418.110 22.540 ;
      LAYER via ;
        RECT 1418.280 1686.100 1418.540 1686.360 ;
        RECT 1685.540 1686.100 1685.800 1686.360 ;
        RECT 1043.380 22.480 1043.640 22.740 ;
        RECT 1417.820 22.480 1418.080 22.740 ;
      LAYER met2 ;
        RECT 1685.460 1700.000 1685.740 1702.400 ;
        RECT 1685.600 1686.390 1685.740 1700.000 ;
        RECT 1418.280 1686.070 1418.540 1686.390 ;
        RECT 1685.540 1686.070 1685.800 1686.390 ;
        RECT 1418.340 39.850 1418.480 1686.070 ;
        RECT 1417.880 39.710 1418.480 39.850 ;
        RECT 1417.880 22.770 1418.020 39.710 ;
        RECT 1043.380 22.450 1043.640 22.770 ;
        RECT 1417.820 22.450 1418.080 22.770 ;
        RECT 1043.440 2.400 1043.580 22.450 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1424.690 1686.640 1425.010 1686.700 ;
        RECT 1694.710 1686.640 1695.030 1686.700 ;
        RECT 1424.690 1686.500 1695.030 1686.640 ;
        RECT 1424.690 1686.440 1425.010 1686.500 ;
        RECT 1694.710 1686.440 1695.030 1686.500 ;
        RECT 1061.290 22.340 1061.610 22.400 ;
        RECT 1424.690 22.340 1425.010 22.400 ;
        RECT 1061.290 22.200 1425.010 22.340 ;
        RECT 1061.290 22.140 1061.610 22.200 ;
        RECT 1424.690 22.140 1425.010 22.200 ;
      LAYER via ;
        RECT 1424.720 1686.440 1424.980 1686.700 ;
        RECT 1694.740 1686.440 1695.000 1686.700 ;
        RECT 1061.320 22.140 1061.580 22.400 ;
        RECT 1424.720 22.140 1424.980 22.400 ;
      LAYER met2 ;
        RECT 1694.660 1700.000 1694.940 1702.400 ;
        RECT 1694.800 1686.730 1694.940 1700.000 ;
        RECT 1424.720 1686.410 1424.980 1686.730 ;
        RECT 1694.740 1686.410 1695.000 1686.730 ;
        RECT 1424.780 22.430 1424.920 1686.410 ;
        RECT 1061.320 22.110 1061.580 22.430 ;
        RECT 1424.720 22.110 1424.980 22.430 ;
        RECT 1061.380 2.400 1061.520 22.110 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.470 1678.140 1697.790 1678.200 ;
        RECT 1702.070 1678.140 1702.390 1678.200 ;
        RECT 1697.470 1678.000 1702.390 1678.140 ;
        RECT 1697.470 1677.940 1697.790 1678.000 ;
        RECT 1702.070 1677.940 1702.390 1678.000 ;
        RECT 1079.230 23.700 1079.550 23.760 ;
        RECT 1697.470 23.700 1697.790 23.760 ;
        RECT 1079.230 23.560 1697.790 23.700 ;
        RECT 1079.230 23.500 1079.550 23.560 ;
        RECT 1697.470 23.500 1697.790 23.560 ;
      LAYER via ;
        RECT 1697.500 1677.940 1697.760 1678.200 ;
        RECT 1702.100 1677.940 1702.360 1678.200 ;
        RECT 1079.260 23.500 1079.520 23.760 ;
        RECT 1697.500 23.500 1697.760 23.760 ;
      LAYER met2 ;
        RECT 1703.860 1700.410 1704.140 1702.400 ;
        RECT 1702.160 1700.270 1704.140 1700.410 ;
        RECT 1702.160 1678.230 1702.300 1700.270 ;
        RECT 1703.860 1700.000 1704.140 1700.270 ;
        RECT 1697.500 1677.910 1697.760 1678.230 ;
        RECT 1702.100 1677.910 1702.360 1678.230 ;
        RECT 1697.560 23.790 1697.700 1677.910 ;
        RECT 1079.260 23.470 1079.520 23.790 ;
        RECT 1697.500 23.470 1697.760 23.790 ;
        RECT 1079.320 2.400 1079.460 23.470 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1713.060 1700.410 1713.340 1702.400 ;
        RECT 1711.360 1700.270 1713.340 1700.410 ;
        RECT 1711.360 24.325 1711.500 1700.270 ;
        RECT 1713.060 1700.000 1713.340 1700.270 ;
        RECT 1096.730 23.955 1097.010 24.325 ;
        RECT 1711.290 23.955 1711.570 24.325 ;
        RECT 1096.800 2.400 1096.940 23.955 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
      LAYER via2 ;
        RECT 1096.730 24.000 1097.010 24.280 ;
        RECT 1711.290 24.000 1711.570 24.280 ;
      LAYER met3 ;
        RECT 1096.705 24.290 1097.035 24.305 ;
        RECT 1711.265 24.290 1711.595 24.305 ;
        RECT 1096.705 23.990 1711.595 24.290 ;
        RECT 1096.705 23.975 1097.035 23.990 ;
        RECT 1711.265 23.975 1711.595 23.990 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1718.170 1657.740 1718.490 1657.800 ;
        RECT 1720.470 1657.740 1720.790 1657.800 ;
        RECT 1718.170 1657.600 1720.790 1657.740 ;
        RECT 1718.170 1657.540 1718.490 1657.600 ;
        RECT 1720.470 1657.540 1720.790 1657.600 ;
        RECT 1114.650 23.360 1114.970 23.420 ;
        RECT 1718.170 23.360 1718.490 23.420 ;
        RECT 1114.650 23.220 1718.490 23.360 ;
        RECT 1114.650 23.160 1114.970 23.220 ;
        RECT 1718.170 23.160 1718.490 23.220 ;
      LAYER via ;
        RECT 1718.200 1657.540 1718.460 1657.800 ;
        RECT 1720.500 1657.540 1720.760 1657.800 ;
        RECT 1114.680 23.160 1114.940 23.420 ;
        RECT 1718.200 23.160 1718.460 23.420 ;
      LAYER met2 ;
        RECT 1722.260 1700.410 1722.540 1702.400 ;
        RECT 1720.560 1700.270 1722.540 1700.410 ;
        RECT 1720.560 1657.830 1720.700 1700.270 ;
        RECT 1722.260 1700.000 1722.540 1700.270 ;
        RECT 1718.200 1657.510 1718.460 1657.830 ;
        RECT 1720.500 1657.510 1720.760 1657.830 ;
        RECT 1718.260 23.450 1718.400 1657.510 ;
        RECT 1114.680 23.130 1114.940 23.450 ;
        RECT 1718.200 23.130 1718.460 23.450 ;
        RECT 1114.740 2.400 1114.880 23.130 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1725.070 1678.140 1725.390 1678.200 ;
        RECT 1729.670 1678.140 1729.990 1678.200 ;
        RECT 1725.070 1678.000 1729.990 1678.140 ;
        RECT 1725.070 1677.940 1725.390 1678.000 ;
        RECT 1729.670 1677.940 1729.990 1678.000 ;
        RECT 1132.590 23.020 1132.910 23.080 ;
        RECT 1725.070 23.020 1725.390 23.080 ;
        RECT 1132.590 22.880 1725.390 23.020 ;
        RECT 1132.590 22.820 1132.910 22.880 ;
        RECT 1725.070 22.820 1725.390 22.880 ;
      LAYER via ;
        RECT 1725.100 1677.940 1725.360 1678.200 ;
        RECT 1729.700 1677.940 1729.960 1678.200 ;
        RECT 1132.620 22.820 1132.880 23.080 ;
        RECT 1725.100 22.820 1725.360 23.080 ;
      LAYER met2 ;
        RECT 1731.460 1700.410 1731.740 1702.400 ;
        RECT 1729.760 1700.270 1731.740 1700.410 ;
        RECT 1729.760 1678.230 1729.900 1700.270 ;
        RECT 1731.460 1700.000 1731.740 1700.270 ;
        RECT 1725.100 1677.910 1725.360 1678.230 ;
        RECT 1729.700 1677.910 1729.960 1678.230 ;
        RECT 1725.160 23.110 1725.300 1677.910 ;
        RECT 1132.620 22.790 1132.880 23.110 ;
        RECT 1725.100 22.790 1725.360 23.110 ;
        RECT 1132.680 2.400 1132.820 22.790 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1150.530 24.380 1150.850 24.440 ;
        RECT 1738.870 24.380 1739.190 24.440 ;
        RECT 1150.530 24.240 1739.190 24.380 ;
        RECT 1150.530 24.180 1150.850 24.240 ;
        RECT 1738.870 24.180 1739.190 24.240 ;
      LAYER via ;
        RECT 1150.560 24.180 1150.820 24.440 ;
        RECT 1738.900 24.180 1739.160 24.440 ;
      LAYER met2 ;
        RECT 1740.660 1700.410 1740.940 1702.400 ;
        RECT 1738.960 1700.270 1740.940 1700.410 ;
        RECT 1738.960 24.470 1739.100 1700.270 ;
        RECT 1740.660 1700.000 1740.940 1700.270 ;
        RECT 1150.560 24.150 1150.820 24.470 ;
        RECT 1738.900 24.150 1739.160 24.470 ;
        RECT 1150.620 2.400 1150.760 24.150 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 27.100 669.230 27.160 ;
        RECT 1490.470 27.100 1490.790 27.160 ;
        RECT 668.910 26.960 1490.790 27.100 ;
        RECT 668.910 26.900 669.230 26.960 ;
        RECT 1490.470 26.900 1490.790 26.960 ;
      LAYER via ;
        RECT 668.940 26.900 669.200 27.160 ;
        RECT 1490.500 26.900 1490.760 27.160 ;
      LAYER met2 ;
        RECT 1492.720 1700.410 1493.000 1702.400 ;
        RECT 1490.560 1700.270 1493.000 1700.410 ;
        RECT 1490.560 27.190 1490.700 1700.270 ;
        RECT 1492.720 1700.000 1493.000 1700.270 ;
        RECT 668.940 26.870 669.200 27.190 ;
        RECT 1490.500 26.870 1490.760 27.190 ;
        RECT 669.000 2.400 669.140 26.870 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1745.770 1659.100 1746.090 1659.160 ;
        RECT 1748.070 1659.100 1748.390 1659.160 ;
        RECT 1745.770 1658.960 1748.390 1659.100 ;
        RECT 1745.770 1658.900 1746.090 1658.960 ;
        RECT 1748.070 1658.900 1748.390 1658.960 ;
        RECT 1168.470 24.040 1168.790 24.100 ;
        RECT 1745.770 24.040 1746.090 24.100 ;
        RECT 1168.470 23.900 1746.090 24.040 ;
        RECT 1168.470 23.840 1168.790 23.900 ;
        RECT 1745.770 23.840 1746.090 23.900 ;
      LAYER via ;
        RECT 1745.800 1658.900 1746.060 1659.160 ;
        RECT 1748.100 1658.900 1748.360 1659.160 ;
        RECT 1168.500 23.840 1168.760 24.100 ;
        RECT 1745.800 23.840 1746.060 24.100 ;
      LAYER met2 ;
        RECT 1749.860 1700.410 1750.140 1702.400 ;
        RECT 1748.160 1700.270 1750.140 1700.410 ;
        RECT 1748.160 1659.190 1748.300 1700.270 ;
        RECT 1749.860 1700.000 1750.140 1700.270 ;
        RECT 1745.800 1658.870 1746.060 1659.190 ;
        RECT 1748.100 1658.870 1748.360 1659.190 ;
        RECT 1745.860 24.130 1746.000 1658.870 ;
        RECT 1168.500 23.810 1168.760 24.130 ;
        RECT 1745.800 23.810 1746.060 24.130 ;
        RECT 1168.560 2.400 1168.700 23.810 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1752.670 1678.140 1752.990 1678.200 ;
        RECT 1757.270 1678.140 1757.590 1678.200 ;
        RECT 1752.670 1678.000 1757.590 1678.140 ;
        RECT 1752.670 1677.940 1752.990 1678.000 ;
        RECT 1757.270 1677.940 1757.590 1678.000 ;
        RECT 1185.950 24.720 1186.270 24.780 ;
        RECT 1752.670 24.720 1752.990 24.780 ;
        RECT 1185.950 24.580 1752.990 24.720 ;
        RECT 1185.950 24.520 1186.270 24.580 ;
        RECT 1752.670 24.520 1752.990 24.580 ;
      LAYER via ;
        RECT 1752.700 1677.940 1752.960 1678.200 ;
        RECT 1757.300 1677.940 1757.560 1678.200 ;
        RECT 1185.980 24.520 1186.240 24.780 ;
        RECT 1752.700 24.520 1752.960 24.780 ;
      LAYER met2 ;
        RECT 1759.060 1700.410 1759.340 1702.400 ;
        RECT 1757.360 1700.270 1759.340 1700.410 ;
        RECT 1757.360 1678.230 1757.500 1700.270 ;
        RECT 1759.060 1700.000 1759.340 1700.270 ;
        RECT 1752.700 1677.910 1752.960 1678.230 ;
        RECT 1757.300 1677.910 1757.560 1678.230 ;
        RECT 1752.760 24.810 1752.900 1677.910 ;
        RECT 1185.980 24.490 1186.240 24.810 ;
        RECT 1752.700 24.490 1752.960 24.810 ;
        RECT 1186.040 2.400 1186.180 24.490 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 25.060 1204.210 25.120 ;
        RECT 1766.470 25.060 1766.790 25.120 ;
        RECT 1203.890 24.920 1766.790 25.060 ;
        RECT 1203.890 24.860 1204.210 24.920 ;
        RECT 1766.470 24.860 1766.790 24.920 ;
      LAYER via ;
        RECT 1203.920 24.860 1204.180 25.120 ;
        RECT 1766.500 24.860 1766.760 25.120 ;
      LAYER met2 ;
        RECT 1768.260 1700.410 1768.540 1702.400 ;
        RECT 1766.560 1700.270 1768.540 1700.410 ;
        RECT 1766.560 25.150 1766.700 1700.270 ;
        RECT 1768.260 1700.000 1768.540 1700.270 ;
        RECT 1203.920 24.830 1204.180 25.150 ;
        RECT 1766.500 24.830 1766.760 25.150 ;
        RECT 1203.980 2.400 1204.120 24.830 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1773.370 1678.140 1773.690 1678.200 ;
        RECT 1775.670 1678.140 1775.990 1678.200 ;
        RECT 1773.370 1678.000 1775.990 1678.140 ;
        RECT 1773.370 1677.940 1773.690 1678.000 ;
        RECT 1775.670 1677.940 1775.990 1678.000 ;
        RECT 1221.830 25.400 1222.150 25.460 ;
        RECT 1773.370 25.400 1773.690 25.460 ;
        RECT 1221.830 25.260 1773.690 25.400 ;
        RECT 1221.830 25.200 1222.150 25.260 ;
        RECT 1773.370 25.200 1773.690 25.260 ;
      LAYER via ;
        RECT 1773.400 1677.940 1773.660 1678.200 ;
        RECT 1775.700 1677.940 1775.960 1678.200 ;
        RECT 1221.860 25.200 1222.120 25.460 ;
        RECT 1773.400 25.200 1773.660 25.460 ;
      LAYER met2 ;
        RECT 1777.460 1700.410 1777.740 1702.400 ;
        RECT 1775.760 1700.270 1777.740 1700.410 ;
        RECT 1775.760 1678.230 1775.900 1700.270 ;
        RECT 1777.460 1700.000 1777.740 1700.270 ;
        RECT 1773.400 1677.910 1773.660 1678.230 ;
        RECT 1775.700 1677.910 1775.960 1678.230 ;
        RECT 1773.460 25.490 1773.600 1677.910 ;
        RECT 1221.860 25.170 1222.120 25.490 ;
        RECT 1773.400 25.170 1773.660 25.490 ;
        RECT 1221.920 2.400 1222.060 25.170 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1782.645 1628.345 1782.815 1683.595 ;
        RECT 1782.645 1490.645 1782.815 1579.895 ;
        RECT 1782.185 1255.365 1782.355 1270.155 ;
        RECT 1782.185 1145.885 1782.355 1173.595 ;
        RECT 1782.185 1124.465 1782.355 1145.375 ;
        RECT 1782.185 1013.965 1782.355 1055.615 ;
        RECT 1782.185 766.105 1782.355 814.215 ;
        RECT 1782.185 524.705 1782.355 572.475 ;
        RECT 1782.185 476.085 1782.355 524.195 ;
        RECT 1782.185 289.765 1782.355 337.875 ;
      LAYER mcon ;
        RECT 1782.645 1683.425 1782.815 1683.595 ;
        RECT 1782.645 1579.725 1782.815 1579.895 ;
        RECT 1782.185 1269.985 1782.355 1270.155 ;
        RECT 1782.185 1173.425 1782.355 1173.595 ;
        RECT 1782.185 1145.205 1782.355 1145.375 ;
        RECT 1782.185 1055.445 1782.355 1055.615 ;
        RECT 1782.185 814.045 1782.355 814.215 ;
        RECT 1782.185 572.305 1782.355 572.475 ;
        RECT 1782.185 524.025 1782.355 524.195 ;
        RECT 1782.185 337.705 1782.355 337.875 ;
      LAYER met1 ;
        RECT 1782.585 1683.580 1782.875 1683.625 ;
        RECT 1783.950 1683.580 1784.270 1683.640 ;
        RECT 1782.585 1683.440 1784.270 1683.580 ;
        RECT 1782.585 1683.395 1782.875 1683.440 ;
        RECT 1783.950 1683.380 1784.270 1683.440 ;
        RECT 1782.570 1628.500 1782.890 1628.560 ;
        RECT 1782.375 1628.360 1782.890 1628.500 ;
        RECT 1782.570 1628.300 1782.890 1628.360 ;
        RECT 1782.570 1579.880 1782.890 1579.940 ;
        RECT 1782.375 1579.740 1782.890 1579.880 ;
        RECT 1782.570 1579.680 1782.890 1579.740 ;
        RECT 1782.585 1490.800 1782.875 1490.845 ;
        RECT 1783.030 1490.800 1783.350 1490.860 ;
        RECT 1782.585 1490.660 1783.350 1490.800 ;
        RECT 1782.585 1490.615 1782.875 1490.660 ;
        RECT 1783.030 1490.600 1783.350 1490.660 ;
        RECT 1782.110 1448.780 1782.430 1449.040 ;
        RECT 1782.200 1448.640 1782.340 1448.780 ;
        RECT 1782.570 1448.640 1782.890 1448.700 ;
        RECT 1782.200 1448.500 1782.890 1448.640 ;
        RECT 1782.570 1448.440 1782.890 1448.500 ;
        RECT 1782.110 1400.700 1782.430 1400.760 ;
        RECT 1782.570 1400.700 1782.890 1400.760 ;
        RECT 1782.110 1400.560 1782.890 1400.700 ;
        RECT 1782.110 1400.500 1782.430 1400.560 ;
        RECT 1782.570 1400.500 1782.890 1400.560 ;
        RECT 1782.110 1366.500 1782.430 1366.760 ;
        RECT 1782.200 1366.080 1782.340 1366.500 ;
        RECT 1782.110 1365.820 1782.430 1366.080 ;
        RECT 1782.570 1304.480 1782.890 1304.540 ;
        RECT 1782.200 1304.340 1782.890 1304.480 ;
        RECT 1782.200 1303.860 1782.340 1304.340 ;
        RECT 1782.570 1304.280 1782.890 1304.340 ;
        RECT 1782.110 1303.600 1782.430 1303.860 ;
        RECT 1782.110 1270.140 1782.430 1270.200 ;
        RECT 1781.915 1270.000 1782.430 1270.140 ;
        RECT 1782.110 1269.940 1782.430 1270.000 ;
        RECT 1782.110 1255.520 1782.430 1255.580 ;
        RECT 1781.915 1255.380 1782.430 1255.520 ;
        RECT 1782.110 1255.320 1782.430 1255.380 ;
        RECT 1782.110 1221.320 1782.430 1221.580 ;
        RECT 1782.200 1220.840 1782.340 1221.320 ;
        RECT 1782.570 1220.840 1782.890 1220.900 ;
        RECT 1782.200 1220.700 1782.890 1220.840 ;
        RECT 1782.570 1220.640 1782.890 1220.700 ;
        RECT 1782.125 1173.580 1782.415 1173.625 ;
        RECT 1782.570 1173.580 1782.890 1173.640 ;
        RECT 1782.125 1173.440 1782.890 1173.580 ;
        RECT 1782.125 1173.395 1782.415 1173.440 ;
        RECT 1782.570 1173.380 1782.890 1173.440 ;
        RECT 1782.110 1146.040 1782.430 1146.100 ;
        RECT 1781.915 1145.900 1782.430 1146.040 ;
        RECT 1782.110 1145.840 1782.430 1145.900 ;
        RECT 1782.110 1145.360 1782.430 1145.420 ;
        RECT 1781.915 1145.220 1782.430 1145.360 ;
        RECT 1782.110 1145.160 1782.430 1145.220 ;
        RECT 1782.110 1124.620 1782.430 1124.680 ;
        RECT 1781.915 1124.480 1782.430 1124.620 ;
        RECT 1782.110 1124.420 1782.430 1124.480 ;
        RECT 1782.570 1063.080 1782.890 1063.140 ;
        RECT 1782.200 1062.940 1782.890 1063.080 ;
        RECT 1782.200 1062.800 1782.340 1062.940 ;
        RECT 1782.570 1062.880 1782.890 1062.940 ;
        RECT 1782.110 1062.540 1782.430 1062.800 ;
        RECT 1782.110 1055.600 1782.430 1055.660 ;
        RECT 1781.915 1055.460 1782.430 1055.600 ;
        RECT 1782.110 1055.400 1782.430 1055.460 ;
        RECT 1782.110 1014.120 1782.430 1014.180 ;
        RECT 1781.915 1013.980 1782.430 1014.120 ;
        RECT 1782.110 1013.920 1782.430 1013.980 ;
        RECT 1782.570 966.520 1782.890 966.580 ;
        RECT 1782.200 966.380 1782.890 966.520 ;
        RECT 1782.200 966.240 1782.340 966.380 ;
        RECT 1782.570 966.320 1782.890 966.380 ;
        RECT 1782.110 965.980 1782.430 966.240 ;
        RECT 1782.110 869.620 1782.430 869.680 ;
        RECT 1783.030 869.620 1783.350 869.680 ;
        RECT 1782.110 869.480 1783.350 869.620 ;
        RECT 1782.110 869.420 1782.430 869.480 ;
        RECT 1783.030 869.420 1783.350 869.480 ;
        RECT 1782.110 821.000 1782.430 821.060 ;
        RECT 1782.570 821.000 1782.890 821.060 ;
        RECT 1782.110 820.860 1782.890 821.000 ;
        RECT 1782.110 820.800 1782.430 820.860 ;
        RECT 1782.570 820.800 1782.890 820.860 ;
        RECT 1782.110 814.200 1782.430 814.260 ;
        RECT 1781.915 814.060 1782.430 814.200 ;
        RECT 1782.110 814.000 1782.430 814.060 ;
        RECT 1782.110 766.260 1782.430 766.320 ;
        RECT 1781.915 766.120 1782.430 766.260 ;
        RECT 1782.110 766.060 1782.430 766.120 ;
        RECT 1782.110 738.380 1782.430 738.440 ;
        RECT 1782.110 738.240 1782.800 738.380 ;
        RECT 1782.110 738.180 1782.430 738.240 ;
        RECT 1782.660 737.420 1782.800 738.240 ;
        RECT 1782.570 737.160 1782.890 737.420 ;
        RECT 1782.570 724.440 1782.890 724.500 ;
        RECT 1783.030 724.440 1783.350 724.500 ;
        RECT 1782.570 724.300 1783.350 724.440 ;
        RECT 1782.570 724.240 1782.890 724.300 ;
        RECT 1783.030 724.240 1783.350 724.300 ;
        RECT 1782.110 675.960 1782.430 676.220 ;
        RECT 1782.200 675.820 1782.340 675.960 ;
        RECT 1782.570 675.820 1782.890 675.880 ;
        RECT 1782.200 675.680 1782.890 675.820 ;
        RECT 1782.570 675.620 1782.890 675.680 ;
        RECT 1782.110 621.080 1782.430 621.140 ;
        RECT 1782.570 621.080 1782.890 621.140 ;
        RECT 1782.110 620.940 1782.890 621.080 ;
        RECT 1782.110 620.880 1782.430 620.940 ;
        RECT 1782.570 620.880 1782.890 620.940 ;
        RECT 1782.110 579.600 1782.430 579.660 ;
        RECT 1783.030 579.600 1783.350 579.660 ;
        RECT 1782.110 579.460 1783.350 579.600 ;
        RECT 1782.110 579.400 1782.430 579.460 ;
        RECT 1783.030 579.400 1783.350 579.460 ;
        RECT 1782.125 572.460 1782.415 572.505 ;
        RECT 1783.030 572.460 1783.350 572.520 ;
        RECT 1782.125 572.320 1783.350 572.460 ;
        RECT 1782.125 572.275 1782.415 572.320 ;
        RECT 1783.030 572.260 1783.350 572.320 ;
        RECT 1782.110 524.860 1782.430 524.920 ;
        RECT 1781.915 524.720 1782.430 524.860 ;
        RECT 1782.110 524.660 1782.430 524.720 ;
        RECT 1782.110 524.180 1782.430 524.240 ;
        RECT 1781.915 524.040 1782.430 524.180 ;
        RECT 1782.110 523.980 1782.430 524.040 ;
        RECT 1782.125 476.240 1782.415 476.285 ;
        RECT 1783.030 476.240 1783.350 476.300 ;
        RECT 1782.125 476.100 1783.350 476.240 ;
        RECT 1782.125 476.055 1782.415 476.100 ;
        RECT 1783.030 476.040 1783.350 476.100 ;
        RECT 1782.110 427.960 1782.430 428.020 ;
        RECT 1783.030 427.960 1783.350 428.020 ;
        RECT 1782.110 427.820 1783.350 427.960 ;
        RECT 1782.110 427.760 1782.430 427.820 ;
        RECT 1783.030 427.760 1783.350 427.820 ;
        RECT 1782.125 337.860 1782.415 337.905 ;
        RECT 1782.570 337.860 1782.890 337.920 ;
        RECT 1782.125 337.720 1782.890 337.860 ;
        RECT 1782.125 337.675 1782.415 337.720 ;
        RECT 1782.570 337.660 1782.890 337.720 ;
        RECT 1782.110 289.920 1782.430 289.980 ;
        RECT 1781.915 289.780 1782.430 289.920 ;
        RECT 1782.110 289.720 1782.430 289.780 ;
        RECT 1782.110 144.740 1782.430 144.800 ;
        RECT 1782.570 144.740 1782.890 144.800 ;
        RECT 1782.110 144.600 1782.890 144.740 ;
        RECT 1782.110 144.540 1782.430 144.600 ;
        RECT 1782.570 144.540 1782.890 144.600 ;
        RECT 1239.770 25.740 1240.090 25.800 ;
        RECT 1782.110 25.740 1782.430 25.800 ;
        RECT 1239.770 25.600 1782.430 25.740 ;
        RECT 1239.770 25.540 1240.090 25.600 ;
        RECT 1782.110 25.540 1782.430 25.600 ;
      LAYER via ;
        RECT 1783.980 1683.380 1784.240 1683.640 ;
        RECT 1782.600 1628.300 1782.860 1628.560 ;
        RECT 1782.600 1579.680 1782.860 1579.940 ;
        RECT 1783.060 1490.600 1783.320 1490.860 ;
        RECT 1782.140 1448.780 1782.400 1449.040 ;
        RECT 1782.600 1448.440 1782.860 1448.700 ;
        RECT 1782.140 1400.500 1782.400 1400.760 ;
        RECT 1782.600 1400.500 1782.860 1400.760 ;
        RECT 1782.140 1366.500 1782.400 1366.760 ;
        RECT 1782.140 1365.820 1782.400 1366.080 ;
        RECT 1782.600 1304.280 1782.860 1304.540 ;
        RECT 1782.140 1303.600 1782.400 1303.860 ;
        RECT 1782.140 1269.940 1782.400 1270.200 ;
        RECT 1782.140 1255.320 1782.400 1255.580 ;
        RECT 1782.140 1221.320 1782.400 1221.580 ;
        RECT 1782.600 1220.640 1782.860 1220.900 ;
        RECT 1782.600 1173.380 1782.860 1173.640 ;
        RECT 1782.140 1145.840 1782.400 1146.100 ;
        RECT 1782.140 1145.160 1782.400 1145.420 ;
        RECT 1782.140 1124.420 1782.400 1124.680 ;
        RECT 1782.600 1062.880 1782.860 1063.140 ;
        RECT 1782.140 1062.540 1782.400 1062.800 ;
        RECT 1782.140 1055.400 1782.400 1055.660 ;
        RECT 1782.140 1013.920 1782.400 1014.180 ;
        RECT 1782.600 966.320 1782.860 966.580 ;
        RECT 1782.140 965.980 1782.400 966.240 ;
        RECT 1782.140 869.420 1782.400 869.680 ;
        RECT 1783.060 869.420 1783.320 869.680 ;
        RECT 1782.140 820.800 1782.400 821.060 ;
        RECT 1782.600 820.800 1782.860 821.060 ;
        RECT 1782.140 814.000 1782.400 814.260 ;
        RECT 1782.140 766.060 1782.400 766.320 ;
        RECT 1782.140 738.180 1782.400 738.440 ;
        RECT 1782.600 737.160 1782.860 737.420 ;
        RECT 1782.600 724.240 1782.860 724.500 ;
        RECT 1783.060 724.240 1783.320 724.500 ;
        RECT 1782.140 675.960 1782.400 676.220 ;
        RECT 1782.600 675.620 1782.860 675.880 ;
        RECT 1782.140 620.880 1782.400 621.140 ;
        RECT 1782.600 620.880 1782.860 621.140 ;
        RECT 1782.140 579.400 1782.400 579.660 ;
        RECT 1783.060 579.400 1783.320 579.660 ;
        RECT 1783.060 572.260 1783.320 572.520 ;
        RECT 1782.140 524.660 1782.400 524.920 ;
        RECT 1782.140 523.980 1782.400 524.240 ;
        RECT 1783.060 476.040 1783.320 476.300 ;
        RECT 1782.140 427.760 1782.400 428.020 ;
        RECT 1783.060 427.760 1783.320 428.020 ;
        RECT 1782.600 337.660 1782.860 337.920 ;
        RECT 1782.140 289.720 1782.400 289.980 ;
        RECT 1782.140 144.540 1782.400 144.800 ;
        RECT 1782.600 144.540 1782.860 144.800 ;
        RECT 1239.800 25.540 1240.060 25.800 ;
        RECT 1782.140 25.540 1782.400 25.800 ;
      LAYER met2 ;
        RECT 1786.660 1701.090 1786.940 1702.400 ;
        RECT 1784.040 1700.950 1786.940 1701.090 ;
        RECT 1784.040 1683.670 1784.180 1700.950 ;
        RECT 1786.660 1700.000 1786.940 1700.950 ;
        RECT 1783.980 1683.350 1784.240 1683.670 ;
        RECT 1782.600 1628.270 1782.860 1628.590 ;
        RECT 1782.660 1579.970 1782.800 1628.270 ;
        RECT 1782.600 1579.650 1782.860 1579.970 ;
        RECT 1783.060 1490.570 1783.320 1490.890 ;
        RECT 1783.120 1449.490 1783.260 1490.570 ;
        RECT 1782.200 1449.350 1783.260 1449.490 ;
        RECT 1782.200 1449.070 1782.340 1449.350 ;
        RECT 1782.140 1448.750 1782.400 1449.070 ;
        RECT 1782.600 1448.410 1782.860 1448.730 ;
        RECT 1782.660 1400.790 1782.800 1448.410 ;
        RECT 1782.140 1400.470 1782.400 1400.790 ;
        RECT 1782.600 1400.470 1782.860 1400.790 ;
        RECT 1782.200 1366.790 1782.340 1400.470 ;
        RECT 1782.140 1366.470 1782.400 1366.790 ;
        RECT 1782.140 1365.790 1782.400 1366.110 ;
        RECT 1782.200 1345.450 1782.340 1365.790 ;
        RECT 1782.200 1345.310 1782.800 1345.450 ;
        RECT 1782.660 1304.570 1782.800 1345.310 ;
        RECT 1782.600 1304.250 1782.860 1304.570 ;
        RECT 1782.140 1303.570 1782.400 1303.890 ;
        RECT 1782.200 1270.230 1782.340 1303.570 ;
        RECT 1782.140 1269.910 1782.400 1270.230 ;
        RECT 1782.140 1255.290 1782.400 1255.610 ;
        RECT 1782.200 1221.610 1782.340 1255.290 ;
        RECT 1782.140 1221.290 1782.400 1221.610 ;
        RECT 1782.600 1220.610 1782.860 1220.930 ;
        RECT 1782.660 1173.670 1782.800 1220.610 ;
        RECT 1782.600 1173.350 1782.860 1173.670 ;
        RECT 1782.140 1145.810 1782.400 1146.130 ;
        RECT 1782.200 1145.450 1782.340 1145.810 ;
        RECT 1782.140 1145.130 1782.400 1145.450 ;
        RECT 1782.140 1124.390 1782.400 1124.710 ;
        RECT 1782.200 1097.250 1782.340 1124.390 ;
        RECT 1782.200 1097.110 1782.800 1097.250 ;
        RECT 1782.660 1063.170 1782.800 1097.110 ;
        RECT 1782.600 1062.850 1782.860 1063.170 ;
        RECT 1782.140 1062.510 1782.400 1062.830 ;
        RECT 1782.200 1055.690 1782.340 1062.510 ;
        RECT 1782.140 1055.370 1782.400 1055.690 ;
        RECT 1782.140 1013.890 1782.400 1014.210 ;
        RECT 1782.200 1007.490 1782.340 1013.890 ;
        RECT 1782.200 1007.350 1782.800 1007.490 ;
        RECT 1782.660 966.610 1782.800 1007.350 ;
        RECT 1782.600 966.290 1782.860 966.610 ;
        RECT 1782.140 966.010 1782.400 966.270 ;
        RECT 1782.140 965.950 1782.800 966.010 ;
        RECT 1782.200 965.870 1782.800 965.950 ;
        RECT 1782.660 965.330 1782.800 965.870 ;
        RECT 1782.660 965.190 1783.260 965.330 ;
        RECT 1783.120 869.710 1783.260 965.190 ;
        RECT 1782.140 869.565 1782.400 869.710 ;
        RECT 1782.130 869.195 1782.410 869.565 ;
        RECT 1783.060 869.390 1783.320 869.710 ;
        RECT 1782.590 868.515 1782.870 868.885 ;
        RECT 1782.660 821.090 1782.800 868.515 ;
        RECT 1782.140 820.770 1782.400 821.090 ;
        RECT 1782.600 820.770 1782.860 821.090 ;
        RECT 1782.200 814.290 1782.340 820.770 ;
        RECT 1782.140 813.970 1782.400 814.290 ;
        RECT 1782.140 766.030 1782.400 766.350 ;
        RECT 1782.200 738.470 1782.340 766.030 ;
        RECT 1782.140 738.150 1782.400 738.470 ;
        RECT 1782.600 737.130 1782.860 737.450 ;
        RECT 1782.660 724.530 1782.800 737.130 ;
        RECT 1782.600 724.210 1782.860 724.530 ;
        RECT 1783.060 724.210 1783.320 724.530 ;
        RECT 1783.120 676.445 1783.260 724.210 ;
        RECT 1782.130 676.075 1782.410 676.445 ;
        RECT 1783.050 676.075 1783.330 676.445 ;
        RECT 1782.140 675.930 1782.400 676.075 ;
        RECT 1782.600 675.590 1782.860 675.910 ;
        RECT 1782.660 621.170 1782.800 675.590 ;
        RECT 1782.140 620.850 1782.400 621.170 ;
        RECT 1782.600 620.850 1782.860 621.170 ;
        RECT 1782.200 579.690 1782.340 620.850 ;
        RECT 1782.140 579.370 1782.400 579.690 ;
        RECT 1783.060 579.370 1783.320 579.690 ;
        RECT 1783.120 572.550 1783.260 579.370 ;
        RECT 1783.060 572.230 1783.320 572.550 ;
        RECT 1782.140 524.630 1782.400 524.950 ;
        RECT 1782.200 524.270 1782.340 524.630 ;
        RECT 1782.140 523.950 1782.400 524.270 ;
        RECT 1783.060 476.010 1783.320 476.330 ;
        RECT 1783.120 428.050 1783.260 476.010 ;
        RECT 1782.140 427.730 1782.400 428.050 ;
        RECT 1783.060 427.730 1783.320 428.050 ;
        RECT 1782.200 362.850 1782.340 427.730 ;
        RECT 1782.200 362.710 1783.260 362.850 ;
        RECT 1783.120 351.290 1783.260 362.710 ;
        RECT 1782.660 351.150 1783.260 351.290 ;
        RECT 1782.660 337.950 1782.800 351.150 ;
        RECT 1782.600 337.630 1782.860 337.950 ;
        RECT 1782.140 289.690 1782.400 290.010 ;
        RECT 1782.200 289.410 1782.340 289.690 ;
        RECT 1782.200 289.270 1782.800 289.410 ;
        RECT 1782.660 207.810 1782.800 289.270 ;
        RECT 1782.660 207.670 1783.260 207.810 ;
        RECT 1783.120 196.930 1783.260 207.670 ;
        RECT 1782.660 196.790 1783.260 196.930 ;
        RECT 1782.660 144.830 1782.800 196.790 ;
        RECT 1782.140 144.510 1782.400 144.830 ;
        RECT 1782.600 144.510 1782.860 144.830 ;
        RECT 1782.200 25.830 1782.340 144.510 ;
        RECT 1239.800 25.510 1240.060 25.830 ;
        RECT 1782.140 25.510 1782.400 25.830 ;
        RECT 1239.860 2.400 1240.000 25.510 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
      LAYER via2 ;
        RECT 1782.130 869.240 1782.410 869.520 ;
        RECT 1782.590 868.560 1782.870 868.840 ;
        RECT 1782.130 676.120 1782.410 676.400 ;
        RECT 1783.050 676.120 1783.330 676.400 ;
      LAYER met3 ;
        RECT 1782.105 869.530 1782.435 869.545 ;
        RECT 1782.105 869.215 1782.650 869.530 ;
        RECT 1782.350 868.865 1782.650 869.215 ;
        RECT 1782.350 868.550 1782.895 868.865 ;
        RECT 1782.565 868.535 1782.895 868.550 ;
        RECT 1782.105 676.410 1782.435 676.425 ;
        RECT 1783.025 676.410 1783.355 676.425 ;
        RECT 1782.105 676.110 1783.355 676.410 ;
        RECT 1782.105 676.095 1782.435 676.110 ;
        RECT 1783.025 676.095 1783.355 676.110 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1257.250 26.080 1257.570 26.140 ;
        RECT 1794.070 26.080 1794.390 26.140 ;
        RECT 1257.250 25.940 1794.390 26.080 ;
        RECT 1257.250 25.880 1257.570 25.940 ;
        RECT 1794.070 25.880 1794.390 25.940 ;
      LAYER via ;
        RECT 1257.280 25.880 1257.540 26.140 ;
        RECT 1794.100 25.880 1794.360 26.140 ;
      LAYER met2 ;
        RECT 1795.860 1700.410 1796.140 1702.400 ;
        RECT 1794.160 1700.270 1796.140 1700.410 ;
        RECT 1794.160 26.170 1794.300 1700.270 ;
        RECT 1795.860 1700.000 1796.140 1700.270 ;
        RECT 1257.280 25.850 1257.540 26.170 ;
        RECT 1794.100 25.850 1794.360 26.170 ;
        RECT 1257.340 2.400 1257.480 25.850 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.970 1678.140 1801.290 1678.200 ;
        RECT 1803.270 1678.140 1803.590 1678.200 ;
        RECT 1800.970 1678.000 1803.590 1678.140 ;
        RECT 1800.970 1677.940 1801.290 1678.000 ;
        RECT 1803.270 1677.940 1803.590 1678.000 ;
        RECT 1626.630 29.480 1626.950 29.540 ;
        RECT 1800.970 29.480 1801.290 29.540 ;
        RECT 1626.630 29.340 1801.290 29.480 ;
        RECT 1626.630 29.280 1626.950 29.340 ;
        RECT 1800.970 29.280 1801.290 29.340 ;
        RECT 1275.190 19.280 1275.510 19.340 ;
        RECT 1275.190 19.140 1583.620 19.280 ;
        RECT 1275.190 19.080 1275.510 19.140 ;
        RECT 1583.480 18.600 1583.620 19.140 ;
        RECT 1626.630 18.600 1626.950 18.660 ;
        RECT 1583.480 18.460 1626.950 18.600 ;
        RECT 1626.630 18.400 1626.950 18.460 ;
      LAYER via ;
        RECT 1801.000 1677.940 1801.260 1678.200 ;
        RECT 1803.300 1677.940 1803.560 1678.200 ;
        RECT 1626.660 29.280 1626.920 29.540 ;
        RECT 1801.000 29.280 1801.260 29.540 ;
        RECT 1275.220 19.080 1275.480 19.340 ;
        RECT 1626.660 18.400 1626.920 18.660 ;
      LAYER met2 ;
        RECT 1805.060 1700.410 1805.340 1702.400 ;
        RECT 1803.360 1700.270 1805.340 1700.410 ;
        RECT 1803.360 1678.230 1803.500 1700.270 ;
        RECT 1805.060 1700.000 1805.340 1700.270 ;
        RECT 1801.000 1677.910 1801.260 1678.230 ;
        RECT 1803.300 1677.910 1803.560 1678.230 ;
        RECT 1801.060 29.570 1801.200 1677.910 ;
        RECT 1626.660 29.250 1626.920 29.570 ;
        RECT 1801.000 29.250 1801.260 29.570 ;
        RECT 1275.220 19.050 1275.480 19.370 ;
        RECT 1275.280 2.400 1275.420 19.050 ;
        RECT 1626.720 18.690 1626.860 29.250 ;
        RECT 1626.660 18.370 1626.920 18.690 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1808.330 1678.140 1808.650 1678.200 ;
        RECT 1812.470 1678.140 1812.790 1678.200 ;
        RECT 1808.330 1678.000 1812.790 1678.140 ;
        RECT 1808.330 1677.940 1808.650 1678.000 ;
        RECT 1812.470 1677.940 1812.790 1678.000 ;
        RECT 1808.330 46.480 1808.650 46.540 ;
        RECT 1626.720 46.340 1808.650 46.480 ;
        RECT 1612.830 45.800 1613.150 45.860 ;
        RECT 1626.720 45.800 1626.860 46.340 ;
        RECT 1808.330 46.280 1808.650 46.340 ;
        RECT 1612.830 45.660 1626.860 45.800 ;
        RECT 1612.830 45.600 1613.150 45.660 ;
        RECT 1293.130 19.620 1293.450 19.680 ;
        RECT 1612.830 19.620 1613.150 19.680 ;
        RECT 1293.130 19.480 1613.150 19.620 ;
        RECT 1293.130 19.420 1293.450 19.480 ;
        RECT 1612.830 19.420 1613.150 19.480 ;
      LAYER via ;
        RECT 1808.360 1677.940 1808.620 1678.200 ;
        RECT 1812.500 1677.940 1812.760 1678.200 ;
        RECT 1612.860 45.600 1613.120 45.860 ;
        RECT 1808.360 46.280 1808.620 46.540 ;
        RECT 1293.160 19.420 1293.420 19.680 ;
        RECT 1612.860 19.420 1613.120 19.680 ;
      LAYER met2 ;
        RECT 1814.260 1700.410 1814.540 1702.400 ;
        RECT 1812.560 1700.270 1814.540 1700.410 ;
        RECT 1812.560 1678.230 1812.700 1700.270 ;
        RECT 1814.260 1700.000 1814.540 1700.270 ;
        RECT 1808.360 1677.910 1808.620 1678.230 ;
        RECT 1812.500 1677.910 1812.760 1678.230 ;
        RECT 1808.420 46.570 1808.560 1677.910 ;
        RECT 1808.360 46.250 1808.620 46.570 ;
        RECT 1612.860 45.570 1613.120 45.890 ;
        RECT 1612.920 19.710 1613.060 45.570 ;
        RECT 1293.160 19.390 1293.420 19.710 ;
        RECT 1612.860 19.390 1613.120 19.710 ;
        RECT 1293.220 2.400 1293.360 19.390 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1613.290 29.140 1613.610 29.200 ;
        RECT 1821.670 29.140 1821.990 29.200 ;
        RECT 1613.290 29.000 1821.990 29.140 ;
        RECT 1613.290 28.940 1613.610 29.000 ;
        RECT 1821.670 28.940 1821.990 29.000 ;
        RECT 1311.070 20.300 1311.390 20.360 ;
        RECT 1613.290 20.300 1613.610 20.360 ;
        RECT 1311.070 20.160 1613.610 20.300 ;
        RECT 1311.070 20.100 1311.390 20.160 ;
        RECT 1613.290 20.100 1613.610 20.160 ;
      LAYER via ;
        RECT 1613.320 28.940 1613.580 29.200 ;
        RECT 1821.700 28.940 1821.960 29.200 ;
        RECT 1311.100 20.100 1311.360 20.360 ;
        RECT 1613.320 20.100 1613.580 20.360 ;
      LAYER met2 ;
        RECT 1823.460 1700.410 1823.740 1702.400 ;
        RECT 1821.760 1700.270 1823.740 1700.410 ;
        RECT 1821.760 29.230 1821.900 1700.270 ;
        RECT 1823.460 1700.000 1823.740 1700.270 ;
        RECT 1613.320 28.910 1613.580 29.230 ;
        RECT 1821.700 28.910 1821.960 29.230 ;
        RECT 1613.380 20.390 1613.520 28.910 ;
        RECT 1311.100 20.070 1311.360 20.390 ;
        RECT 1613.320 20.070 1613.580 20.390 ;
        RECT 1311.160 2.400 1311.300 20.070 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1829.030 1531.940 1829.350 1532.000 ;
        RECT 1829.950 1531.940 1830.270 1532.000 ;
        RECT 1829.030 1531.800 1830.270 1531.940 ;
        RECT 1829.030 1531.740 1829.350 1531.800 ;
        RECT 1829.950 1531.740 1830.270 1531.800 ;
        RECT 1829.490 1490.260 1829.810 1490.520 ;
        RECT 1829.580 1489.840 1829.720 1490.260 ;
        RECT 1829.490 1489.580 1829.810 1489.840 ;
        RECT 1438.030 52.600 1438.350 52.660 ;
        RECT 1828.110 52.600 1828.430 52.660 ;
        RECT 1438.030 52.460 1828.430 52.600 ;
        RECT 1438.030 52.400 1438.350 52.460 ;
        RECT 1828.110 52.400 1828.430 52.460 ;
        RECT 1329.010 17.580 1329.330 17.640 ;
        RECT 1438.030 17.580 1438.350 17.640 ;
        RECT 1329.010 17.440 1438.350 17.580 ;
        RECT 1329.010 17.380 1329.330 17.440 ;
        RECT 1438.030 17.380 1438.350 17.440 ;
      LAYER via ;
        RECT 1829.060 1531.740 1829.320 1532.000 ;
        RECT 1829.980 1531.740 1830.240 1532.000 ;
        RECT 1829.520 1490.260 1829.780 1490.520 ;
        RECT 1829.520 1489.580 1829.780 1489.840 ;
        RECT 1438.060 52.400 1438.320 52.660 ;
        RECT 1828.140 52.400 1828.400 52.660 ;
        RECT 1329.040 17.380 1329.300 17.640 ;
        RECT 1438.060 17.380 1438.320 17.640 ;
      LAYER met2 ;
        RECT 1832.660 1701.090 1832.940 1702.400 ;
        RECT 1830.040 1700.950 1832.940 1701.090 ;
        RECT 1830.040 1656.210 1830.180 1700.950 ;
        RECT 1832.660 1700.000 1832.940 1700.950 ;
        RECT 1829.580 1656.070 1830.180 1656.210 ;
        RECT 1829.580 1587.530 1829.720 1656.070 ;
        RECT 1829.120 1587.390 1829.720 1587.530 ;
        RECT 1829.120 1580.165 1829.260 1587.390 ;
        RECT 1829.050 1579.795 1829.330 1580.165 ;
        RECT 1829.970 1579.795 1830.250 1580.165 ;
        RECT 1830.040 1532.030 1830.180 1579.795 ;
        RECT 1829.060 1531.710 1829.320 1532.030 ;
        RECT 1829.980 1531.710 1830.240 1532.030 ;
        RECT 1829.120 1497.090 1829.260 1531.710 ;
        RECT 1829.120 1496.950 1829.720 1497.090 ;
        RECT 1829.580 1490.550 1829.720 1496.950 ;
        RECT 1829.520 1490.230 1829.780 1490.550 ;
        RECT 1829.520 1489.550 1829.780 1489.870 ;
        RECT 1829.580 980.290 1829.720 1489.550 ;
        RECT 1829.120 980.150 1829.720 980.290 ;
        RECT 1829.120 979.610 1829.260 980.150 ;
        RECT 1829.120 979.470 1829.720 979.610 ;
        RECT 1829.580 303.690 1829.720 979.470 ;
        RECT 1829.120 303.550 1829.720 303.690 ;
        RECT 1829.120 303.010 1829.260 303.550 ;
        RECT 1829.120 302.870 1829.720 303.010 ;
        RECT 1829.580 207.130 1829.720 302.870 ;
        RECT 1829.120 206.990 1829.720 207.130 ;
        RECT 1829.120 206.450 1829.260 206.990 ;
        RECT 1829.120 206.310 1829.720 206.450 ;
        RECT 1829.580 96.970 1829.720 206.310 ;
        RECT 1829.120 96.830 1829.720 96.970 ;
        RECT 1829.120 62.970 1829.260 96.830 ;
        RECT 1828.200 62.830 1829.260 62.970 ;
        RECT 1828.200 52.690 1828.340 62.830 ;
        RECT 1438.060 52.370 1438.320 52.690 ;
        RECT 1828.140 52.370 1828.400 52.690 ;
        RECT 1438.120 17.670 1438.260 52.370 ;
        RECT 1329.040 17.350 1329.300 17.670 ;
        RECT 1438.060 17.350 1438.320 17.670 ;
        RECT 1329.100 2.400 1329.240 17.350 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
      LAYER via2 ;
        RECT 1829.050 1579.840 1829.330 1580.120 ;
        RECT 1829.970 1579.840 1830.250 1580.120 ;
      LAYER met3 ;
        RECT 1829.025 1580.130 1829.355 1580.145 ;
        RECT 1829.945 1580.130 1830.275 1580.145 ;
        RECT 1829.025 1579.830 1830.275 1580.130 ;
        RECT 1829.025 1579.815 1829.355 1579.830 ;
        RECT 1829.945 1579.815 1830.275 1579.830 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1497.370 1678.140 1497.690 1678.200 ;
        RECT 1500.590 1678.140 1500.910 1678.200 ;
        RECT 1497.370 1678.000 1500.910 1678.140 ;
        RECT 1497.370 1677.940 1497.690 1678.000 ;
        RECT 1500.590 1677.940 1500.910 1678.000 ;
        RECT 686.390 27.440 686.710 27.500 ;
        RECT 1497.370 27.440 1497.690 27.500 ;
        RECT 686.390 27.300 1497.690 27.440 ;
        RECT 686.390 27.240 686.710 27.300 ;
        RECT 1497.370 27.240 1497.690 27.300 ;
      LAYER via ;
        RECT 1497.400 1677.940 1497.660 1678.200 ;
        RECT 1500.620 1677.940 1500.880 1678.200 ;
        RECT 686.420 27.240 686.680 27.500 ;
        RECT 1497.400 27.240 1497.660 27.500 ;
      LAYER met2 ;
        RECT 1501.920 1700.410 1502.200 1702.400 ;
        RECT 1500.680 1700.270 1502.200 1700.410 ;
        RECT 1500.680 1678.230 1500.820 1700.270 ;
        RECT 1501.920 1700.000 1502.200 1700.270 ;
        RECT 1497.400 1677.910 1497.660 1678.230 ;
        RECT 1500.620 1677.910 1500.880 1678.230 ;
        RECT 1497.460 27.530 1497.600 1677.910 ;
        RECT 686.420 27.210 686.680 27.530 ;
        RECT 1497.400 27.210 1497.660 27.530 ;
        RECT 686.480 2.400 686.620 27.210 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1835.930 1678.140 1836.250 1678.200 ;
        RECT 1840.070 1678.140 1840.390 1678.200 ;
        RECT 1835.930 1678.000 1840.390 1678.140 ;
        RECT 1835.930 1677.940 1836.250 1678.000 ;
        RECT 1840.070 1677.940 1840.390 1678.000 ;
        RECT 1449.070 53.280 1449.390 53.340 ;
        RECT 1835.930 53.280 1836.250 53.340 ;
        RECT 1449.070 53.140 1836.250 53.280 ;
        RECT 1449.070 53.080 1449.390 53.140 ;
        RECT 1835.930 53.080 1836.250 53.140 ;
        RECT 1346.490 18.260 1346.810 18.320 ;
        RECT 1449.070 18.260 1449.390 18.320 ;
        RECT 1346.490 18.120 1449.390 18.260 ;
        RECT 1346.490 18.060 1346.810 18.120 ;
        RECT 1449.070 18.060 1449.390 18.120 ;
      LAYER via ;
        RECT 1835.960 1677.940 1836.220 1678.200 ;
        RECT 1840.100 1677.940 1840.360 1678.200 ;
        RECT 1449.100 53.080 1449.360 53.340 ;
        RECT 1835.960 53.080 1836.220 53.340 ;
        RECT 1346.520 18.060 1346.780 18.320 ;
        RECT 1449.100 18.060 1449.360 18.320 ;
      LAYER met2 ;
        RECT 1841.860 1700.410 1842.140 1702.400 ;
        RECT 1840.160 1700.270 1842.140 1700.410 ;
        RECT 1840.160 1678.230 1840.300 1700.270 ;
        RECT 1841.860 1700.000 1842.140 1700.270 ;
        RECT 1835.960 1677.910 1836.220 1678.230 ;
        RECT 1840.100 1677.910 1840.360 1678.230 ;
        RECT 1836.020 53.370 1836.160 1677.910 ;
        RECT 1449.100 53.050 1449.360 53.370 ;
        RECT 1835.960 53.050 1836.220 53.370 ;
        RECT 1449.160 18.350 1449.300 53.050 ;
        RECT 1346.520 18.030 1346.780 18.350 ;
        RECT 1449.100 18.030 1449.360 18.350 ;
        RECT 1346.580 2.400 1346.720 18.030 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1582.930 29.820 1583.250 29.880 ;
        RECT 1849.270 29.820 1849.590 29.880 ;
        RECT 1582.930 29.680 1849.590 29.820 ;
        RECT 1582.930 29.620 1583.250 29.680 ;
        RECT 1849.270 29.620 1849.590 29.680 ;
        RECT 1364.430 18.940 1364.750 19.000 ;
        RECT 1582.930 18.940 1583.250 19.000 ;
        RECT 1364.430 18.800 1583.250 18.940 ;
        RECT 1364.430 18.740 1364.750 18.800 ;
        RECT 1582.930 18.740 1583.250 18.800 ;
      LAYER via ;
        RECT 1582.960 29.620 1583.220 29.880 ;
        RECT 1849.300 29.620 1849.560 29.880 ;
        RECT 1364.460 18.740 1364.720 19.000 ;
        RECT 1582.960 18.740 1583.220 19.000 ;
      LAYER met2 ;
        RECT 1851.060 1700.410 1851.340 1702.400 ;
        RECT 1849.360 1700.270 1851.340 1700.410 ;
        RECT 1849.360 29.910 1849.500 1700.270 ;
        RECT 1851.060 1700.000 1851.340 1700.270 ;
        RECT 1582.960 29.590 1583.220 29.910 ;
        RECT 1849.300 29.590 1849.560 29.910 ;
        RECT 1583.020 19.030 1583.160 29.590 ;
        RECT 1364.460 18.710 1364.720 19.030 ;
        RECT 1582.960 18.710 1583.220 19.030 ;
        RECT 1364.520 2.400 1364.660 18.710 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1856.705 1546.405 1856.875 1593.835 ;
        RECT 1857.165 1352.605 1857.335 1400.715 ;
        RECT 1857.165 1256.045 1857.335 1304.155 ;
        RECT 1857.165 283.305 1857.335 303.195 ;
        RECT 1857.165 235.025 1857.335 282.795 ;
        RECT 1400.845 16.405 1401.015 20.655 ;
      LAYER mcon ;
        RECT 1856.705 1593.665 1856.875 1593.835 ;
        RECT 1857.165 1400.545 1857.335 1400.715 ;
        RECT 1857.165 1303.985 1857.335 1304.155 ;
        RECT 1857.165 303.025 1857.335 303.195 ;
        RECT 1857.165 282.625 1857.335 282.795 ;
        RECT 1400.845 20.485 1401.015 20.655 ;
      LAYER met1 ;
        RECT 1856.645 1593.820 1856.935 1593.865 ;
        RECT 1857.090 1593.820 1857.410 1593.880 ;
        RECT 1856.645 1593.680 1857.410 1593.820 ;
        RECT 1856.645 1593.635 1856.935 1593.680 ;
        RECT 1857.090 1593.620 1857.410 1593.680 ;
        RECT 1856.630 1546.560 1856.950 1546.620 ;
        RECT 1856.435 1546.420 1856.950 1546.560 ;
        RECT 1856.630 1546.360 1856.950 1546.420 ;
        RECT 1856.170 1490.800 1856.490 1490.860 ;
        RECT 1858.010 1490.800 1858.330 1490.860 ;
        RECT 1856.170 1490.660 1858.330 1490.800 ;
        RECT 1856.170 1490.600 1856.490 1490.660 ;
        RECT 1858.010 1490.600 1858.330 1490.660 ;
        RECT 1857.090 1400.700 1857.410 1400.760 ;
        RECT 1856.895 1400.560 1857.410 1400.700 ;
        RECT 1857.090 1400.500 1857.410 1400.560 ;
        RECT 1857.090 1352.760 1857.410 1352.820 ;
        RECT 1856.895 1352.620 1857.410 1352.760 ;
        RECT 1857.090 1352.560 1857.410 1352.620 ;
        RECT 1857.090 1304.140 1857.410 1304.200 ;
        RECT 1856.895 1304.000 1857.410 1304.140 ;
        RECT 1857.090 1303.940 1857.410 1304.000 ;
        RECT 1857.090 1256.200 1857.410 1256.260 ;
        RECT 1856.895 1256.060 1857.410 1256.200 ;
        RECT 1857.090 1256.000 1857.410 1256.060 ;
        RECT 1857.090 1172.700 1857.410 1172.960 ;
        RECT 1857.180 1172.280 1857.320 1172.700 ;
        RECT 1857.090 1172.020 1857.410 1172.280 ;
        RECT 1857.090 1076.140 1857.410 1076.400 ;
        RECT 1857.180 1075.720 1857.320 1076.140 ;
        RECT 1857.090 1075.460 1857.410 1075.720 ;
        RECT 1857.090 979.580 1857.410 979.840 ;
        RECT 1857.180 979.160 1857.320 979.580 ;
        RECT 1857.090 978.900 1857.410 979.160 ;
        RECT 1857.090 883.020 1857.410 883.280 ;
        RECT 1857.180 882.600 1857.320 883.020 ;
        RECT 1857.090 882.340 1857.410 882.600 ;
        RECT 1857.090 786.460 1857.410 786.720 ;
        RECT 1857.180 786.040 1857.320 786.460 ;
        RECT 1857.090 785.780 1857.410 786.040 ;
        RECT 1857.090 400.220 1857.410 400.480 ;
        RECT 1857.180 399.800 1857.320 400.220 ;
        RECT 1857.090 399.540 1857.410 399.800 ;
        RECT 1857.090 303.180 1857.410 303.240 ;
        RECT 1856.895 303.040 1857.410 303.180 ;
        RECT 1857.090 302.980 1857.410 303.040 ;
        RECT 1857.090 283.460 1857.410 283.520 ;
        RECT 1856.895 283.320 1857.410 283.460 ;
        RECT 1857.090 283.260 1857.410 283.320 ;
        RECT 1857.090 282.780 1857.410 282.840 ;
        RECT 1857.090 282.640 1857.605 282.780 ;
        RECT 1857.090 282.580 1857.410 282.640 ;
        RECT 1856.630 235.180 1856.950 235.240 ;
        RECT 1857.105 235.180 1857.395 235.225 ;
        RECT 1856.630 235.040 1857.395 235.180 ;
        RECT 1856.630 234.980 1856.950 235.040 ;
        RECT 1857.105 234.995 1857.395 235.040 ;
        RECT 1856.630 234.300 1856.950 234.560 ;
        RECT 1856.720 234.160 1856.860 234.300 ;
        RECT 1857.550 234.160 1857.870 234.220 ;
        RECT 1856.720 234.020 1857.870 234.160 ;
        RECT 1857.550 233.960 1857.870 234.020 ;
        RECT 1856.630 96.800 1856.950 96.860 ;
        RECT 1857.550 96.800 1857.870 96.860 ;
        RECT 1856.630 96.660 1857.870 96.800 ;
        RECT 1856.630 96.600 1856.950 96.660 ;
        RECT 1857.550 96.600 1857.870 96.660 ;
        RECT 1573.270 30.500 1573.590 30.560 ;
        RECT 1856.630 30.500 1856.950 30.560 ;
        RECT 1573.270 30.360 1856.950 30.500 ;
        RECT 1573.270 30.300 1573.590 30.360 ;
        RECT 1856.630 30.300 1856.950 30.360 ;
        RECT 1573.270 20.980 1573.590 21.040 ;
        RECT 1572.440 20.840 1573.590 20.980 ;
        RECT 1400.785 20.640 1401.075 20.685 ;
        RECT 1572.440 20.640 1572.580 20.840 ;
        RECT 1573.270 20.780 1573.590 20.840 ;
        RECT 1400.785 20.500 1572.580 20.640 ;
        RECT 1400.785 20.455 1401.075 20.500 ;
        RECT 1382.370 16.560 1382.690 16.620 ;
        RECT 1400.785 16.560 1401.075 16.605 ;
        RECT 1382.370 16.420 1401.075 16.560 ;
        RECT 1382.370 16.360 1382.690 16.420 ;
        RECT 1400.785 16.375 1401.075 16.420 ;
      LAYER via ;
        RECT 1857.120 1593.620 1857.380 1593.880 ;
        RECT 1856.660 1546.360 1856.920 1546.620 ;
        RECT 1856.200 1490.600 1856.460 1490.860 ;
        RECT 1858.040 1490.600 1858.300 1490.860 ;
        RECT 1857.120 1400.500 1857.380 1400.760 ;
        RECT 1857.120 1352.560 1857.380 1352.820 ;
        RECT 1857.120 1303.940 1857.380 1304.200 ;
        RECT 1857.120 1256.000 1857.380 1256.260 ;
        RECT 1857.120 1172.700 1857.380 1172.960 ;
        RECT 1857.120 1172.020 1857.380 1172.280 ;
        RECT 1857.120 1076.140 1857.380 1076.400 ;
        RECT 1857.120 1075.460 1857.380 1075.720 ;
        RECT 1857.120 979.580 1857.380 979.840 ;
        RECT 1857.120 978.900 1857.380 979.160 ;
        RECT 1857.120 883.020 1857.380 883.280 ;
        RECT 1857.120 882.340 1857.380 882.600 ;
        RECT 1857.120 786.460 1857.380 786.720 ;
        RECT 1857.120 785.780 1857.380 786.040 ;
        RECT 1857.120 400.220 1857.380 400.480 ;
        RECT 1857.120 399.540 1857.380 399.800 ;
        RECT 1857.120 302.980 1857.380 303.240 ;
        RECT 1857.120 283.260 1857.380 283.520 ;
        RECT 1857.120 282.580 1857.380 282.840 ;
        RECT 1856.660 234.980 1856.920 235.240 ;
        RECT 1856.660 234.300 1856.920 234.560 ;
        RECT 1857.580 233.960 1857.840 234.220 ;
        RECT 1856.660 96.600 1856.920 96.860 ;
        RECT 1857.580 96.600 1857.840 96.860 ;
        RECT 1573.300 30.300 1573.560 30.560 ;
        RECT 1856.660 30.300 1856.920 30.560 ;
        RECT 1573.300 20.780 1573.560 21.040 ;
        RECT 1382.400 16.360 1382.660 16.620 ;
      LAYER met2 ;
        RECT 1859.800 1700.410 1860.080 1702.400 ;
        RECT 1858.100 1700.270 1860.080 1700.410 ;
        RECT 1858.100 1656.210 1858.240 1700.270 ;
        RECT 1859.800 1700.000 1860.080 1700.270 ;
        RECT 1857.180 1656.070 1858.240 1656.210 ;
        RECT 1857.180 1608.610 1857.320 1656.070 ;
        RECT 1857.180 1608.470 1857.780 1608.610 ;
        RECT 1857.640 1594.330 1857.780 1608.470 ;
        RECT 1857.180 1594.190 1857.780 1594.330 ;
        RECT 1857.180 1593.910 1857.320 1594.190 ;
        RECT 1857.120 1593.590 1857.380 1593.910 ;
        RECT 1856.660 1546.330 1856.920 1546.650 ;
        RECT 1856.720 1537.890 1856.860 1546.330 ;
        RECT 1856.260 1537.750 1856.860 1537.890 ;
        RECT 1856.260 1490.890 1856.400 1537.750 ;
        RECT 1856.200 1490.570 1856.460 1490.890 ;
        RECT 1858.040 1490.570 1858.300 1490.890 ;
        RECT 1858.100 1463.090 1858.240 1490.570 ;
        RECT 1857.180 1462.950 1858.240 1463.090 ;
        RECT 1857.180 1400.790 1857.320 1462.950 ;
        RECT 1857.120 1400.470 1857.380 1400.790 ;
        RECT 1857.120 1352.530 1857.380 1352.850 ;
        RECT 1857.180 1304.230 1857.320 1352.530 ;
        RECT 1857.120 1303.910 1857.380 1304.230 ;
        RECT 1857.120 1255.970 1857.380 1256.290 ;
        RECT 1857.180 1172.990 1857.320 1255.970 ;
        RECT 1857.120 1172.670 1857.380 1172.990 ;
        RECT 1857.120 1171.990 1857.380 1172.310 ;
        RECT 1857.180 1076.430 1857.320 1171.990 ;
        RECT 1857.120 1076.110 1857.380 1076.430 ;
        RECT 1857.120 1075.430 1857.380 1075.750 ;
        RECT 1857.180 979.870 1857.320 1075.430 ;
        RECT 1857.120 979.550 1857.380 979.870 ;
        RECT 1857.120 978.870 1857.380 979.190 ;
        RECT 1857.180 883.310 1857.320 978.870 ;
        RECT 1857.120 882.990 1857.380 883.310 ;
        RECT 1857.120 882.310 1857.380 882.630 ;
        RECT 1857.180 786.750 1857.320 882.310 ;
        RECT 1857.120 786.430 1857.380 786.750 ;
        RECT 1857.120 785.750 1857.380 786.070 ;
        RECT 1857.180 400.510 1857.320 785.750 ;
        RECT 1857.120 400.190 1857.380 400.510 ;
        RECT 1857.120 399.510 1857.380 399.830 ;
        RECT 1857.180 303.270 1857.320 399.510 ;
        RECT 1857.120 302.950 1857.380 303.270 ;
        RECT 1857.120 283.230 1857.380 283.550 ;
        RECT 1857.180 282.870 1857.320 283.230 ;
        RECT 1857.120 282.550 1857.380 282.870 ;
        RECT 1856.660 234.950 1856.920 235.270 ;
        RECT 1856.720 234.590 1856.860 234.950 ;
        RECT 1856.660 234.270 1856.920 234.590 ;
        RECT 1857.580 233.930 1857.840 234.250 ;
        RECT 1857.640 96.890 1857.780 233.930 ;
        RECT 1856.660 96.570 1856.920 96.890 ;
        RECT 1857.580 96.570 1857.840 96.890 ;
        RECT 1856.720 30.590 1856.860 96.570 ;
        RECT 1573.300 30.270 1573.560 30.590 ;
        RECT 1856.660 30.270 1856.920 30.590 ;
        RECT 1573.360 21.070 1573.500 30.270 ;
        RECT 1573.300 20.750 1573.560 21.070 ;
        RECT 1382.400 16.330 1382.660 16.650 ;
        RECT 1382.460 2.400 1382.600 16.330 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1399.850 30.840 1400.170 30.900 ;
        RECT 1863.990 30.840 1864.310 30.900 ;
        RECT 1399.850 30.700 1864.310 30.840 ;
        RECT 1399.850 30.640 1400.170 30.700 ;
        RECT 1863.990 30.640 1864.310 30.700 ;
      LAYER via ;
        RECT 1399.880 30.640 1400.140 30.900 ;
        RECT 1864.020 30.640 1864.280 30.900 ;
      LAYER met2 ;
        RECT 1869.000 1701.090 1869.280 1702.400 ;
        RECT 1866.840 1700.950 1869.280 1701.090 ;
        RECT 1866.840 1656.210 1866.980 1700.950 ;
        RECT 1869.000 1700.000 1869.280 1700.950 ;
        RECT 1864.080 1656.070 1866.980 1656.210 ;
        RECT 1864.080 30.930 1864.220 1656.070 ;
        RECT 1399.880 30.610 1400.140 30.930 ;
        RECT 1864.020 30.610 1864.280 30.930 ;
        RECT 1399.940 14.010 1400.080 30.610 ;
        RECT 1399.940 13.870 1400.540 14.010 ;
        RECT 1400.400 2.400 1400.540 13.870 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1418.250 31.180 1418.570 31.240 ;
        RECT 1876.870 31.180 1877.190 31.240 ;
        RECT 1418.250 31.040 1877.190 31.180 ;
        RECT 1418.250 30.980 1418.570 31.040 ;
        RECT 1876.870 30.980 1877.190 31.040 ;
      LAYER via ;
        RECT 1418.280 30.980 1418.540 31.240 ;
        RECT 1876.900 30.980 1877.160 31.240 ;
      LAYER met2 ;
        RECT 1878.200 1700.410 1878.480 1702.400 ;
        RECT 1876.960 1700.270 1878.480 1700.410 ;
        RECT 1876.960 31.270 1877.100 1700.270 ;
        RECT 1878.200 1700.000 1878.480 1700.270 ;
        RECT 1418.280 30.950 1418.540 31.270 ;
        RECT 1876.900 30.950 1877.160 31.270 ;
        RECT 1418.340 2.400 1418.480 30.950 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1884.305 1546.405 1884.475 1593.835 ;
        RECT 1884.305 1497.445 1884.475 1545.555 ;
        RECT 1884.765 1352.605 1884.935 1400.715 ;
        RECT 1884.765 1256.045 1884.935 1304.155 ;
        RECT 1884.765 579.785 1884.935 627.895 ;
        RECT 1884.765 483.225 1884.935 531.335 ;
      LAYER mcon ;
        RECT 1884.305 1593.665 1884.475 1593.835 ;
        RECT 1884.305 1545.385 1884.475 1545.555 ;
        RECT 1884.765 1400.545 1884.935 1400.715 ;
        RECT 1884.765 1303.985 1884.935 1304.155 ;
        RECT 1884.765 627.725 1884.935 627.895 ;
        RECT 1884.765 531.165 1884.935 531.335 ;
      LAYER met1 ;
        RECT 1884.245 1593.820 1884.535 1593.865 ;
        RECT 1884.690 1593.820 1885.010 1593.880 ;
        RECT 1884.245 1593.680 1885.010 1593.820 ;
        RECT 1884.245 1593.635 1884.535 1593.680 ;
        RECT 1884.690 1593.620 1885.010 1593.680 ;
        RECT 1884.230 1546.560 1884.550 1546.620 ;
        RECT 1884.035 1546.420 1884.550 1546.560 ;
        RECT 1884.230 1546.360 1884.550 1546.420 ;
        RECT 1884.230 1545.540 1884.550 1545.600 ;
        RECT 1884.035 1545.400 1884.550 1545.540 ;
        RECT 1884.230 1545.340 1884.550 1545.400 ;
        RECT 1884.245 1497.600 1884.535 1497.645 ;
        RECT 1884.690 1497.600 1885.010 1497.660 ;
        RECT 1884.245 1497.460 1885.010 1497.600 ;
        RECT 1884.245 1497.415 1884.535 1497.460 ;
        RECT 1884.690 1497.400 1885.010 1497.460 ;
        RECT 1884.230 1449.660 1884.550 1449.720 ;
        RECT 1884.230 1449.520 1884.920 1449.660 ;
        RECT 1884.230 1449.460 1884.550 1449.520 ;
        RECT 1884.780 1449.380 1884.920 1449.520 ;
        RECT 1884.690 1449.120 1885.010 1449.380 ;
        RECT 1884.690 1400.700 1885.010 1400.760 ;
        RECT 1884.495 1400.560 1885.010 1400.700 ;
        RECT 1884.690 1400.500 1885.010 1400.560 ;
        RECT 1884.690 1352.760 1885.010 1352.820 ;
        RECT 1884.495 1352.620 1885.010 1352.760 ;
        RECT 1884.690 1352.560 1885.010 1352.620 ;
        RECT 1884.690 1304.140 1885.010 1304.200 ;
        RECT 1884.495 1304.000 1885.010 1304.140 ;
        RECT 1884.690 1303.940 1885.010 1304.000 ;
        RECT 1884.690 1256.200 1885.010 1256.260 ;
        RECT 1884.495 1256.060 1885.010 1256.200 ;
        RECT 1884.690 1256.000 1885.010 1256.060 ;
        RECT 1883.770 1159.300 1884.090 1159.360 ;
        RECT 1884.690 1159.300 1885.010 1159.360 ;
        RECT 1883.770 1159.160 1885.010 1159.300 ;
        RECT 1883.770 1159.100 1884.090 1159.160 ;
        RECT 1884.690 1159.100 1885.010 1159.160 ;
        RECT 1883.770 1062.740 1884.090 1062.800 ;
        RECT 1884.690 1062.740 1885.010 1062.800 ;
        RECT 1883.770 1062.600 1885.010 1062.740 ;
        RECT 1883.770 1062.540 1884.090 1062.600 ;
        RECT 1884.690 1062.540 1885.010 1062.600 ;
        RECT 1883.770 966.180 1884.090 966.240 ;
        RECT 1884.690 966.180 1885.010 966.240 ;
        RECT 1883.770 966.040 1885.010 966.180 ;
        RECT 1883.770 965.980 1884.090 966.040 ;
        RECT 1884.690 965.980 1885.010 966.040 ;
        RECT 1883.770 869.620 1884.090 869.680 ;
        RECT 1884.690 869.620 1885.010 869.680 ;
        RECT 1883.770 869.480 1885.010 869.620 ;
        RECT 1883.770 869.420 1884.090 869.480 ;
        RECT 1884.690 869.420 1885.010 869.480 ;
        RECT 1883.770 821.000 1884.090 821.060 ;
        RECT 1884.690 821.000 1885.010 821.060 ;
        RECT 1883.770 820.860 1885.010 821.000 ;
        RECT 1883.770 820.800 1884.090 820.860 ;
        RECT 1884.690 820.800 1885.010 820.860 ;
        RECT 1883.770 724.440 1884.090 724.500 ;
        RECT 1884.690 724.440 1885.010 724.500 ;
        RECT 1883.770 724.300 1885.010 724.440 ;
        RECT 1883.770 724.240 1884.090 724.300 ;
        RECT 1884.690 724.240 1885.010 724.300 ;
        RECT 1884.690 627.880 1885.010 627.940 ;
        RECT 1884.495 627.740 1885.010 627.880 ;
        RECT 1884.690 627.680 1885.010 627.740 ;
        RECT 1884.690 579.940 1885.010 580.000 ;
        RECT 1884.495 579.800 1885.010 579.940 ;
        RECT 1884.690 579.740 1885.010 579.800 ;
        RECT 1884.690 531.320 1885.010 531.380 ;
        RECT 1884.495 531.180 1885.010 531.320 ;
        RECT 1884.690 531.120 1885.010 531.180 ;
        RECT 1884.690 483.380 1885.010 483.440 ;
        RECT 1884.495 483.240 1885.010 483.380 ;
        RECT 1884.690 483.180 1885.010 483.240 ;
        RECT 1884.690 400.220 1885.010 400.480 ;
        RECT 1884.780 399.800 1884.920 400.220 ;
        RECT 1884.690 399.540 1885.010 399.800 ;
        RECT 1884.690 289.580 1885.010 289.640 ;
        RECT 1885.150 289.580 1885.470 289.640 ;
        RECT 1884.690 289.440 1885.470 289.580 ;
        RECT 1884.690 289.380 1885.010 289.440 ;
        RECT 1885.150 289.380 1885.470 289.440 ;
        RECT 1884.690 193.360 1885.010 193.420 ;
        RECT 1885.150 193.360 1885.470 193.420 ;
        RECT 1884.690 193.220 1885.470 193.360 ;
        RECT 1884.690 193.160 1885.010 193.220 ;
        RECT 1885.150 193.160 1885.470 193.220 ;
        RECT 1435.730 31.520 1436.050 31.580 ;
        RECT 1884.690 31.520 1885.010 31.580 ;
        RECT 1435.730 31.380 1885.010 31.520 ;
        RECT 1435.730 31.320 1436.050 31.380 ;
        RECT 1884.690 31.320 1885.010 31.380 ;
      LAYER via ;
        RECT 1884.720 1593.620 1884.980 1593.880 ;
        RECT 1884.260 1546.360 1884.520 1546.620 ;
        RECT 1884.260 1545.340 1884.520 1545.600 ;
        RECT 1884.720 1497.400 1884.980 1497.660 ;
        RECT 1884.260 1449.460 1884.520 1449.720 ;
        RECT 1884.720 1449.120 1884.980 1449.380 ;
        RECT 1884.720 1400.500 1884.980 1400.760 ;
        RECT 1884.720 1352.560 1884.980 1352.820 ;
        RECT 1884.720 1303.940 1884.980 1304.200 ;
        RECT 1884.720 1256.000 1884.980 1256.260 ;
        RECT 1883.800 1159.100 1884.060 1159.360 ;
        RECT 1884.720 1159.100 1884.980 1159.360 ;
        RECT 1883.800 1062.540 1884.060 1062.800 ;
        RECT 1884.720 1062.540 1884.980 1062.800 ;
        RECT 1883.800 965.980 1884.060 966.240 ;
        RECT 1884.720 965.980 1884.980 966.240 ;
        RECT 1883.800 869.420 1884.060 869.680 ;
        RECT 1884.720 869.420 1884.980 869.680 ;
        RECT 1883.800 820.800 1884.060 821.060 ;
        RECT 1884.720 820.800 1884.980 821.060 ;
        RECT 1883.800 724.240 1884.060 724.500 ;
        RECT 1884.720 724.240 1884.980 724.500 ;
        RECT 1884.720 627.680 1884.980 627.940 ;
        RECT 1884.720 579.740 1884.980 580.000 ;
        RECT 1884.720 531.120 1884.980 531.380 ;
        RECT 1884.720 483.180 1884.980 483.440 ;
        RECT 1884.720 400.220 1884.980 400.480 ;
        RECT 1884.720 399.540 1884.980 399.800 ;
        RECT 1884.720 289.380 1884.980 289.640 ;
        RECT 1885.180 289.380 1885.440 289.640 ;
        RECT 1884.720 193.160 1884.980 193.420 ;
        RECT 1885.180 193.160 1885.440 193.420 ;
        RECT 1435.760 31.320 1436.020 31.580 ;
        RECT 1884.720 31.320 1884.980 31.580 ;
      LAYER met2 ;
        RECT 1887.400 1700.410 1887.680 1702.400 ;
        RECT 1886.160 1700.270 1887.680 1700.410 ;
        RECT 1886.160 1677.970 1886.300 1700.270 ;
        RECT 1887.400 1700.000 1887.680 1700.270 ;
        RECT 1884.780 1677.830 1886.300 1677.970 ;
        RECT 1884.780 1608.610 1884.920 1677.830 ;
        RECT 1884.780 1608.470 1885.380 1608.610 ;
        RECT 1885.240 1594.330 1885.380 1608.470 ;
        RECT 1884.780 1594.190 1885.380 1594.330 ;
        RECT 1884.780 1593.910 1884.920 1594.190 ;
        RECT 1884.720 1593.590 1884.980 1593.910 ;
        RECT 1884.260 1546.330 1884.520 1546.650 ;
        RECT 1884.320 1545.630 1884.460 1546.330 ;
        RECT 1884.260 1545.310 1884.520 1545.630 ;
        RECT 1884.720 1497.370 1884.980 1497.690 ;
        RECT 1884.780 1463.090 1884.920 1497.370 ;
        RECT 1884.320 1462.950 1884.920 1463.090 ;
        RECT 1884.320 1449.750 1884.460 1462.950 ;
        RECT 1884.260 1449.430 1884.520 1449.750 ;
        RECT 1884.720 1449.090 1884.980 1449.410 ;
        RECT 1884.780 1400.790 1884.920 1449.090 ;
        RECT 1884.720 1400.470 1884.980 1400.790 ;
        RECT 1884.720 1352.530 1884.980 1352.850 ;
        RECT 1884.780 1304.230 1884.920 1352.530 ;
        RECT 1884.720 1303.910 1884.980 1304.230 ;
        RECT 1884.720 1255.970 1884.980 1256.290 ;
        RECT 1884.780 1207.525 1884.920 1255.970 ;
        RECT 1883.790 1207.155 1884.070 1207.525 ;
        RECT 1884.710 1207.155 1884.990 1207.525 ;
        RECT 1883.860 1159.390 1884.000 1207.155 ;
        RECT 1883.800 1159.070 1884.060 1159.390 ;
        RECT 1884.720 1159.070 1884.980 1159.390 ;
        RECT 1884.780 1110.965 1884.920 1159.070 ;
        RECT 1883.790 1110.595 1884.070 1110.965 ;
        RECT 1884.710 1110.595 1884.990 1110.965 ;
        RECT 1883.860 1062.830 1884.000 1110.595 ;
        RECT 1883.800 1062.510 1884.060 1062.830 ;
        RECT 1884.720 1062.510 1884.980 1062.830 ;
        RECT 1884.780 1014.405 1884.920 1062.510 ;
        RECT 1883.790 1014.035 1884.070 1014.405 ;
        RECT 1884.710 1014.035 1884.990 1014.405 ;
        RECT 1883.860 966.270 1884.000 1014.035 ;
        RECT 1883.800 965.950 1884.060 966.270 ;
        RECT 1884.720 965.950 1884.980 966.270 ;
        RECT 1884.780 917.845 1884.920 965.950 ;
        RECT 1883.790 917.475 1884.070 917.845 ;
        RECT 1884.710 917.475 1884.990 917.845 ;
        RECT 1883.860 869.710 1884.000 917.475 ;
        RECT 1883.800 869.390 1884.060 869.710 ;
        RECT 1884.720 869.390 1884.980 869.710 ;
        RECT 1884.780 821.090 1884.920 869.390 ;
        RECT 1883.800 820.770 1884.060 821.090 ;
        RECT 1884.720 820.770 1884.980 821.090 ;
        RECT 1883.860 773.005 1884.000 820.770 ;
        RECT 1883.790 772.635 1884.070 773.005 ;
        RECT 1884.710 772.635 1884.990 773.005 ;
        RECT 1884.780 724.530 1884.920 772.635 ;
        RECT 1883.800 724.210 1884.060 724.530 ;
        RECT 1884.720 724.210 1884.980 724.530 ;
        RECT 1883.860 676.445 1884.000 724.210 ;
        RECT 1883.790 676.075 1884.070 676.445 ;
        RECT 1884.710 676.075 1884.990 676.445 ;
        RECT 1884.780 627.970 1884.920 676.075 ;
        RECT 1884.720 627.650 1884.980 627.970 ;
        RECT 1884.720 579.710 1884.980 580.030 ;
        RECT 1884.780 531.410 1884.920 579.710 ;
        RECT 1884.720 531.090 1884.980 531.410 ;
        RECT 1884.720 483.150 1884.980 483.470 ;
        RECT 1884.780 400.510 1884.920 483.150 ;
        RECT 1884.720 400.190 1884.980 400.510 ;
        RECT 1884.720 399.510 1884.980 399.830 ;
        RECT 1884.780 303.690 1884.920 399.510 ;
        RECT 1884.320 303.550 1884.920 303.690 ;
        RECT 1884.320 303.010 1884.460 303.550 ;
        RECT 1884.320 302.870 1884.920 303.010 ;
        RECT 1884.780 289.670 1884.920 302.870 ;
        RECT 1884.720 289.350 1884.980 289.670 ;
        RECT 1885.180 289.350 1885.440 289.670 ;
        RECT 1885.240 193.450 1885.380 289.350 ;
        RECT 1884.720 193.130 1884.980 193.450 ;
        RECT 1885.180 193.130 1885.440 193.450 ;
        RECT 1884.780 169.050 1884.920 193.130 ;
        RECT 1884.320 168.910 1884.920 169.050 ;
        RECT 1884.320 130.970 1884.460 168.910 ;
        RECT 1884.320 130.830 1884.920 130.970 ;
        RECT 1884.780 31.610 1884.920 130.830 ;
        RECT 1435.760 31.290 1436.020 31.610 ;
        RECT 1884.720 31.290 1884.980 31.610 ;
        RECT 1435.820 2.400 1435.960 31.290 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
      LAYER via2 ;
        RECT 1883.790 1207.200 1884.070 1207.480 ;
        RECT 1884.710 1207.200 1884.990 1207.480 ;
        RECT 1883.790 1110.640 1884.070 1110.920 ;
        RECT 1884.710 1110.640 1884.990 1110.920 ;
        RECT 1883.790 1014.080 1884.070 1014.360 ;
        RECT 1884.710 1014.080 1884.990 1014.360 ;
        RECT 1883.790 917.520 1884.070 917.800 ;
        RECT 1884.710 917.520 1884.990 917.800 ;
        RECT 1883.790 772.680 1884.070 772.960 ;
        RECT 1884.710 772.680 1884.990 772.960 ;
        RECT 1883.790 676.120 1884.070 676.400 ;
        RECT 1884.710 676.120 1884.990 676.400 ;
      LAYER met3 ;
        RECT 1883.765 1207.490 1884.095 1207.505 ;
        RECT 1884.685 1207.490 1885.015 1207.505 ;
        RECT 1883.765 1207.190 1885.015 1207.490 ;
        RECT 1883.765 1207.175 1884.095 1207.190 ;
        RECT 1884.685 1207.175 1885.015 1207.190 ;
        RECT 1883.765 1110.930 1884.095 1110.945 ;
        RECT 1884.685 1110.930 1885.015 1110.945 ;
        RECT 1883.765 1110.630 1885.015 1110.930 ;
        RECT 1883.765 1110.615 1884.095 1110.630 ;
        RECT 1884.685 1110.615 1885.015 1110.630 ;
        RECT 1883.765 1014.370 1884.095 1014.385 ;
        RECT 1884.685 1014.370 1885.015 1014.385 ;
        RECT 1883.765 1014.070 1885.015 1014.370 ;
        RECT 1883.765 1014.055 1884.095 1014.070 ;
        RECT 1884.685 1014.055 1885.015 1014.070 ;
        RECT 1883.765 917.810 1884.095 917.825 ;
        RECT 1884.685 917.810 1885.015 917.825 ;
        RECT 1883.765 917.510 1885.015 917.810 ;
        RECT 1883.765 917.495 1884.095 917.510 ;
        RECT 1884.685 917.495 1885.015 917.510 ;
        RECT 1883.765 772.970 1884.095 772.985 ;
        RECT 1884.685 772.970 1885.015 772.985 ;
        RECT 1883.765 772.670 1885.015 772.970 ;
        RECT 1883.765 772.655 1884.095 772.670 ;
        RECT 1884.685 772.655 1885.015 772.670 ;
        RECT 1883.765 676.410 1884.095 676.425 ;
        RECT 1884.685 676.410 1885.015 676.425 ;
        RECT 1883.765 676.110 1885.015 676.410 ;
        RECT 1883.765 676.095 1884.095 676.110 ;
        RECT 1884.685 676.095 1885.015 676.110 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1891.130 1678.140 1891.450 1678.200 ;
        RECT 1895.270 1678.140 1895.590 1678.200 ;
        RECT 1891.130 1678.000 1895.590 1678.140 ;
        RECT 1891.130 1677.940 1891.450 1678.000 ;
        RECT 1895.270 1677.940 1895.590 1678.000 ;
        RECT 1453.670 31.860 1453.990 31.920 ;
        RECT 1891.130 31.860 1891.450 31.920 ;
        RECT 1453.670 31.720 1891.450 31.860 ;
        RECT 1453.670 31.660 1453.990 31.720 ;
        RECT 1891.130 31.660 1891.450 31.720 ;
      LAYER via ;
        RECT 1891.160 1677.940 1891.420 1678.200 ;
        RECT 1895.300 1677.940 1895.560 1678.200 ;
        RECT 1453.700 31.660 1453.960 31.920 ;
        RECT 1891.160 31.660 1891.420 31.920 ;
      LAYER met2 ;
        RECT 1896.600 1700.410 1896.880 1702.400 ;
        RECT 1895.360 1700.270 1896.880 1700.410 ;
        RECT 1895.360 1678.230 1895.500 1700.270 ;
        RECT 1896.600 1700.000 1896.880 1700.270 ;
        RECT 1891.160 1677.910 1891.420 1678.230 ;
        RECT 1895.300 1677.910 1895.560 1678.230 ;
        RECT 1891.220 31.950 1891.360 1677.910 ;
        RECT 1453.700 31.630 1453.960 31.950 ;
        RECT 1891.160 31.630 1891.420 31.950 ;
        RECT 1453.760 2.400 1453.900 31.630 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1471.610 26.420 1471.930 26.480 ;
        RECT 1904.470 26.420 1904.790 26.480 ;
        RECT 1471.610 26.280 1904.790 26.420 ;
        RECT 1471.610 26.220 1471.930 26.280 ;
        RECT 1904.470 26.220 1904.790 26.280 ;
      LAYER via ;
        RECT 1471.640 26.220 1471.900 26.480 ;
        RECT 1904.500 26.220 1904.760 26.480 ;
      LAYER met2 ;
        RECT 1905.800 1700.410 1906.080 1702.400 ;
        RECT 1904.560 1700.270 1906.080 1700.410 ;
        RECT 1904.560 26.510 1904.700 1700.270 ;
        RECT 1905.800 1700.000 1906.080 1700.270 ;
        RECT 1471.640 26.190 1471.900 26.510 ;
        RECT 1904.500 26.190 1904.760 26.510 ;
        RECT 1471.700 2.400 1471.840 26.190 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1911.445 1510.365 1911.615 1587.035 ;
        RECT 1912.365 1449.165 1912.535 1497.275 ;
        RECT 1911.905 241.485 1912.075 289.595 ;
        RECT 1911.905 41.565 1912.075 89.675 ;
      LAYER mcon ;
        RECT 1911.445 1586.865 1911.615 1587.035 ;
        RECT 1912.365 1497.105 1912.535 1497.275 ;
        RECT 1911.905 289.425 1912.075 289.595 ;
        RECT 1911.905 89.505 1912.075 89.675 ;
      LAYER met1 ;
        RECT 1911.370 1593.820 1911.690 1593.880 ;
        RECT 1912.290 1593.820 1912.610 1593.880 ;
        RECT 1911.370 1593.680 1912.610 1593.820 ;
        RECT 1911.370 1593.620 1911.690 1593.680 ;
        RECT 1912.290 1593.620 1912.610 1593.680 ;
        RECT 1911.370 1587.020 1911.690 1587.080 ;
        RECT 1911.175 1586.880 1911.690 1587.020 ;
        RECT 1911.370 1586.820 1911.690 1586.880 ;
        RECT 1911.385 1510.520 1911.675 1510.565 ;
        RECT 1912.290 1510.520 1912.610 1510.580 ;
        RECT 1911.385 1510.380 1912.610 1510.520 ;
        RECT 1911.385 1510.335 1911.675 1510.380 ;
        RECT 1912.290 1510.320 1912.610 1510.380 ;
        RECT 1912.290 1497.260 1912.610 1497.320 ;
        RECT 1912.095 1497.120 1912.610 1497.260 ;
        RECT 1912.290 1497.060 1912.610 1497.120 ;
        RECT 1912.290 1449.320 1912.610 1449.380 ;
        RECT 1912.095 1449.180 1912.610 1449.320 ;
        RECT 1912.290 1449.120 1912.610 1449.180 ;
        RECT 1912.290 1365.820 1912.610 1366.080 ;
        RECT 1912.380 1365.400 1912.520 1365.820 ;
        RECT 1912.290 1365.140 1912.610 1365.400 ;
        RECT 1912.290 1269.260 1912.610 1269.520 ;
        RECT 1912.380 1268.840 1912.520 1269.260 ;
        RECT 1912.290 1268.580 1912.610 1268.840 ;
        RECT 1912.290 1172.700 1912.610 1172.960 ;
        RECT 1912.380 1172.280 1912.520 1172.700 ;
        RECT 1912.290 1172.020 1912.610 1172.280 ;
        RECT 1912.290 1076.140 1912.610 1076.400 ;
        RECT 1912.380 1075.720 1912.520 1076.140 ;
        RECT 1912.290 1075.460 1912.610 1075.720 ;
        RECT 1912.290 979.580 1912.610 979.840 ;
        RECT 1912.380 979.160 1912.520 979.580 ;
        RECT 1912.290 978.900 1912.610 979.160 ;
        RECT 1912.290 883.020 1912.610 883.280 ;
        RECT 1912.380 882.600 1912.520 883.020 ;
        RECT 1912.290 882.340 1912.610 882.600 ;
        RECT 1912.290 786.460 1912.610 786.720 ;
        RECT 1912.380 786.040 1912.520 786.460 ;
        RECT 1912.290 785.780 1912.610 786.040 ;
        RECT 1912.290 400.220 1912.610 400.480 ;
        RECT 1912.380 399.800 1912.520 400.220 ;
        RECT 1912.290 399.540 1912.610 399.800 ;
        RECT 1911.845 289.580 1912.135 289.625 ;
        RECT 1912.290 289.580 1912.610 289.640 ;
        RECT 1911.845 289.440 1912.610 289.580 ;
        RECT 1911.845 289.395 1912.135 289.440 ;
        RECT 1912.290 289.380 1912.610 289.440 ;
        RECT 1911.830 241.640 1912.150 241.700 ;
        RECT 1911.635 241.500 1912.150 241.640 ;
        RECT 1911.830 241.440 1912.150 241.500 ;
        RECT 1911.830 193.500 1912.150 193.760 ;
        RECT 1911.920 193.080 1912.060 193.500 ;
        RECT 1911.830 192.820 1912.150 193.080 ;
        RECT 1911.370 96.800 1911.690 96.860 ;
        RECT 1912.290 96.800 1912.610 96.860 ;
        RECT 1911.370 96.660 1912.610 96.800 ;
        RECT 1911.370 96.600 1911.690 96.660 ;
        RECT 1912.290 96.600 1912.610 96.660 ;
        RECT 1911.845 89.660 1912.135 89.705 ;
        RECT 1912.290 89.660 1912.610 89.720 ;
        RECT 1911.845 89.520 1912.610 89.660 ;
        RECT 1911.845 89.475 1912.135 89.520 ;
        RECT 1912.290 89.460 1912.610 89.520 ;
        RECT 1911.830 41.720 1912.150 41.780 ;
        RECT 1911.635 41.580 1912.150 41.720 ;
        RECT 1911.830 41.520 1912.150 41.580 ;
        RECT 1489.550 26.760 1489.870 26.820 ;
        RECT 1911.830 26.760 1912.150 26.820 ;
        RECT 1489.550 26.620 1912.150 26.760 ;
        RECT 1489.550 26.560 1489.870 26.620 ;
        RECT 1911.830 26.560 1912.150 26.620 ;
      LAYER via ;
        RECT 1911.400 1593.620 1911.660 1593.880 ;
        RECT 1912.320 1593.620 1912.580 1593.880 ;
        RECT 1911.400 1586.820 1911.660 1587.080 ;
        RECT 1912.320 1510.320 1912.580 1510.580 ;
        RECT 1912.320 1497.060 1912.580 1497.320 ;
        RECT 1912.320 1449.120 1912.580 1449.380 ;
        RECT 1912.320 1365.820 1912.580 1366.080 ;
        RECT 1912.320 1365.140 1912.580 1365.400 ;
        RECT 1912.320 1269.260 1912.580 1269.520 ;
        RECT 1912.320 1268.580 1912.580 1268.840 ;
        RECT 1912.320 1172.700 1912.580 1172.960 ;
        RECT 1912.320 1172.020 1912.580 1172.280 ;
        RECT 1912.320 1076.140 1912.580 1076.400 ;
        RECT 1912.320 1075.460 1912.580 1075.720 ;
        RECT 1912.320 979.580 1912.580 979.840 ;
        RECT 1912.320 978.900 1912.580 979.160 ;
        RECT 1912.320 883.020 1912.580 883.280 ;
        RECT 1912.320 882.340 1912.580 882.600 ;
        RECT 1912.320 786.460 1912.580 786.720 ;
        RECT 1912.320 785.780 1912.580 786.040 ;
        RECT 1912.320 400.220 1912.580 400.480 ;
        RECT 1912.320 399.540 1912.580 399.800 ;
        RECT 1912.320 289.380 1912.580 289.640 ;
        RECT 1911.860 241.440 1912.120 241.700 ;
        RECT 1911.860 193.500 1912.120 193.760 ;
        RECT 1911.860 192.820 1912.120 193.080 ;
        RECT 1911.400 96.600 1911.660 96.860 ;
        RECT 1912.320 96.600 1912.580 96.860 ;
        RECT 1912.320 89.460 1912.580 89.720 ;
        RECT 1911.860 41.520 1912.120 41.780 ;
        RECT 1489.580 26.560 1489.840 26.820 ;
        RECT 1911.860 26.560 1912.120 26.820 ;
      LAYER met2 ;
        RECT 1915.000 1701.090 1915.280 1702.400 ;
        RECT 1913.300 1700.950 1915.280 1701.090 ;
        RECT 1913.300 1656.210 1913.440 1700.950 ;
        RECT 1915.000 1700.000 1915.280 1700.950 ;
        RECT 1912.380 1656.070 1913.440 1656.210 ;
        RECT 1912.380 1593.910 1912.520 1656.070 ;
        RECT 1911.400 1593.590 1911.660 1593.910 ;
        RECT 1912.320 1593.590 1912.580 1593.910 ;
        RECT 1911.460 1587.110 1911.600 1593.590 ;
        RECT 1911.400 1586.790 1911.660 1587.110 ;
        RECT 1912.320 1510.290 1912.580 1510.610 ;
        RECT 1912.380 1497.350 1912.520 1510.290 ;
        RECT 1912.320 1497.030 1912.580 1497.350 ;
        RECT 1912.320 1449.090 1912.580 1449.410 ;
        RECT 1912.380 1366.110 1912.520 1449.090 ;
        RECT 1912.320 1365.790 1912.580 1366.110 ;
        RECT 1912.320 1365.110 1912.580 1365.430 ;
        RECT 1912.380 1269.550 1912.520 1365.110 ;
        RECT 1912.320 1269.230 1912.580 1269.550 ;
        RECT 1912.320 1268.550 1912.580 1268.870 ;
        RECT 1912.380 1172.990 1912.520 1268.550 ;
        RECT 1912.320 1172.670 1912.580 1172.990 ;
        RECT 1912.320 1171.990 1912.580 1172.310 ;
        RECT 1912.380 1076.430 1912.520 1171.990 ;
        RECT 1912.320 1076.110 1912.580 1076.430 ;
        RECT 1912.320 1075.430 1912.580 1075.750 ;
        RECT 1912.380 979.870 1912.520 1075.430 ;
        RECT 1912.320 979.550 1912.580 979.870 ;
        RECT 1912.320 978.870 1912.580 979.190 ;
        RECT 1912.380 883.310 1912.520 978.870 ;
        RECT 1912.320 882.990 1912.580 883.310 ;
        RECT 1912.320 882.310 1912.580 882.630 ;
        RECT 1912.380 786.750 1912.520 882.310 ;
        RECT 1912.320 786.430 1912.580 786.750 ;
        RECT 1912.320 785.750 1912.580 786.070 ;
        RECT 1912.380 400.510 1912.520 785.750 ;
        RECT 1912.320 400.190 1912.580 400.510 ;
        RECT 1912.320 399.510 1912.580 399.830 ;
        RECT 1912.380 303.690 1912.520 399.510 ;
        RECT 1911.920 303.550 1912.520 303.690 ;
        RECT 1911.920 303.010 1912.060 303.550 ;
        RECT 1911.920 302.870 1912.520 303.010 ;
        RECT 1912.380 289.670 1912.520 302.870 ;
        RECT 1912.320 289.350 1912.580 289.670 ;
        RECT 1911.860 241.410 1912.120 241.730 ;
        RECT 1911.920 193.790 1912.060 241.410 ;
        RECT 1911.860 193.470 1912.120 193.790 ;
        RECT 1911.860 192.790 1912.120 193.110 ;
        RECT 1911.920 169.050 1912.060 192.790 ;
        RECT 1911.460 168.910 1912.060 169.050 ;
        RECT 1911.460 96.890 1911.600 168.910 ;
        RECT 1911.400 96.570 1911.660 96.890 ;
        RECT 1912.320 96.570 1912.580 96.890 ;
        RECT 1912.380 89.750 1912.520 96.570 ;
        RECT 1912.320 89.430 1912.580 89.750 ;
        RECT 1911.860 41.490 1912.120 41.810 ;
        RECT 1911.920 26.850 1912.060 41.490 ;
        RECT 1489.580 26.530 1489.840 26.850 ;
        RECT 1911.860 26.530 1912.120 26.850 ;
        RECT 1489.640 2.400 1489.780 26.530 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1507.030 27.100 1507.350 27.160 ;
        RECT 1919.190 27.100 1919.510 27.160 ;
        RECT 1507.030 26.960 1919.510 27.100 ;
        RECT 1507.030 26.900 1507.350 26.960 ;
        RECT 1919.190 26.900 1919.510 26.960 ;
      LAYER via ;
        RECT 1507.060 26.900 1507.320 27.160 ;
        RECT 1919.220 26.900 1919.480 27.160 ;
      LAYER met2 ;
        RECT 1924.200 1701.090 1924.480 1702.400 ;
        RECT 1922.040 1700.950 1924.480 1701.090 ;
        RECT 1922.040 1656.210 1922.180 1700.950 ;
        RECT 1924.200 1700.000 1924.480 1700.950 ;
        RECT 1919.280 1656.070 1922.180 1656.210 ;
        RECT 1919.280 27.190 1919.420 1656.070 ;
        RECT 1507.060 26.870 1507.320 27.190 ;
        RECT 1919.220 26.870 1919.480 27.190 ;
        RECT 1507.120 2.400 1507.260 26.870 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 710.310 59.740 710.630 59.800 ;
        RECT 1512.090 59.740 1512.410 59.800 ;
        RECT 710.310 59.600 1512.410 59.740 ;
        RECT 710.310 59.540 710.630 59.600 ;
        RECT 1512.090 59.540 1512.410 59.600 ;
        RECT 704.330 20.980 704.650 21.040 ;
        RECT 710.310 20.980 710.630 21.040 ;
        RECT 704.330 20.840 710.630 20.980 ;
        RECT 704.330 20.780 704.650 20.840 ;
        RECT 710.310 20.780 710.630 20.840 ;
      LAYER via ;
        RECT 710.340 59.540 710.600 59.800 ;
        RECT 1512.120 59.540 1512.380 59.800 ;
        RECT 704.360 20.780 704.620 21.040 ;
        RECT 710.340 20.780 710.600 21.040 ;
      LAYER met2 ;
        RECT 1511.120 1700.410 1511.400 1702.400 ;
        RECT 1511.120 1700.270 1512.320 1700.410 ;
        RECT 1511.120 1700.000 1511.400 1700.270 ;
        RECT 1512.180 59.830 1512.320 1700.270 ;
        RECT 710.340 59.510 710.600 59.830 ;
        RECT 1512.120 59.510 1512.380 59.830 ;
        RECT 710.400 21.070 710.540 59.510 ;
        RECT 704.360 20.750 704.620 21.070 ;
        RECT 710.340 20.750 710.600 21.070 ;
        RECT 704.420 2.400 704.560 20.750 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.970 32.200 1525.290 32.260 ;
        RECT 1932.070 32.200 1932.390 32.260 ;
        RECT 1524.970 32.060 1932.390 32.200 ;
        RECT 1524.970 32.000 1525.290 32.060 ;
        RECT 1932.070 32.000 1932.390 32.060 ;
      LAYER via ;
        RECT 1525.000 32.000 1525.260 32.260 ;
        RECT 1932.100 32.000 1932.360 32.260 ;
      LAYER met2 ;
        RECT 1933.400 1700.410 1933.680 1702.400 ;
        RECT 1932.160 1700.270 1933.680 1700.410 ;
        RECT 1932.160 32.290 1932.300 1700.270 ;
        RECT 1933.400 1700.000 1933.680 1700.270 ;
        RECT 1525.000 31.970 1525.260 32.290 ;
        RECT 1932.100 31.970 1932.360 32.290 ;
        RECT 1525.060 2.400 1525.200 31.970 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1939.505 1538.925 1939.675 1587.035 ;
        RECT 1939.505 1490.645 1939.675 1524.475 ;
        RECT 1939.965 789.905 1940.135 814.215 ;
        RECT 1939.965 524.365 1940.135 572.475 ;
        RECT 1939.965 427.805 1940.135 475.915 ;
        RECT 1939.965 282.965 1940.135 331.075 ;
        RECT 1939.505 186.405 1939.675 234.515 ;
        RECT 1939.045 138.125 1939.215 138.975 ;
      LAYER mcon ;
        RECT 1939.505 1586.865 1939.675 1587.035 ;
        RECT 1939.505 1524.305 1939.675 1524.475 ;
        RECT 1939.965 814.045 1940.135 814.215 ;
        RECT 1939.965 572.305 1940.135 572.475 ;
        RECT 1939.965 475.745 1940.135 475.915 ;
        RECT 1939.965 330.905 1940.135 331.075 ;
        RECT 1939.505 234.345 1939.675 234.515 ;
        RECT 1939.045 138.805 1939.215 138.975 ;
      LAYER met1 ;
        RECT 1939.430 1593.820 1939.750 1593.880 ;
        RECT 1939.890 1593.820 1940.210 1593.880 ;
        RECT 1939.430 1593.680 1940.210 1593.820 ;
        RECT 1939.430 1593.620 1939.750 1593.680 ;
        RECT 1939.890 1593.620 1940.210 1593.680 ;
        RECT 1939.430 1587.020 1939.750 1587.080 ;
        RECT 1939.235 1586.880 1939.750 1587.020 ;
        RECT 1939.430 1586.820 1939.750 1586.880 ;
        RECT 1939.430 1539.080 1939.750 1539.140 ;
        RECT 1939.235 1538.940 1939.750 1539.080 ;
        RECT 1939.430 1538.880 1939.750 1538.940 ;
        RECT 1939.430 1524.460 1939.750 1524.520 ;
        RECT 1939.235 1524.320 1939.750 1524.460 ;
        RECT 1939.430 1524.260 1939.750 1524.320 ;
        RECT 1939.445 1490.800 1939.735 1490.845 ;
        RECT 1939.890 1490.800 1940.210 1490.860 ;
        RECT 1939.445 1490.660 1940.210 1490.800 ;
        RECT 1939.445 1490.615 1939.735 1490.660 ;
        RECT 1939.890 1490.600 1940.210 1490.660 ;
        RECT 1939.890 1463.060 1940.210 1463.320 ;
        RECT 1939.980 1462.640 1940.120 1463.060 ;
        RECT 1939.890 1462.380 1940.210 1462.640 ;
        RECT 1939.890 1400.700 1940.210 1400.760 ;
        RECT 1940.350 1400.700 1940.670 1400.760 ;
        RECT 1939.890 1400.560 1940.670 1400.700 ;
        RECT 1939.890 1400.500 1940.210 1400.560 ;
        RECT 1940.350 1400.500 1940.670 1400.560 ;
        RECT 1939.890 814.200 1940.210 814.260 ;
        RECT 1939.695 814.060 1940.210 814.200 ;
        RECT 1939.890 814.000 1940.210 814.060 ;
        RECT 1939.890 790.060 1940.210 790.120 ;
        RECT 1939.695 789.920 1940.210 790.060 ;
        RECT 1939.890 789.860 1940.210 789.920 ;
        RECT 1939.890 627.880 1940.210 627.940 ;
        RECT 1940.350 627.880 1940.670 627.940 ;
        RECT 1939.890 627.740 1940.670 627.880 ;
        RECT 1939.890 627.680 1940.210 627.740 ;
        RECT 1940.350 627.680 1940.670 627.740 ;
        RECT 1939.890 593.200 1940.210 593.260 ;
        RECT 1940.350 593.200 1940.670 593.260 ;
        RECT 1939.890 593.060 1940.670 593.200 ;
        RECT 1939.890 593.000 1940.210 593.060 ;
        RECT 1940.350 593.000 1940.670 593.060 ;
        RECT 1939.890 572.460 1940.210 572.520 ;
        RECT 1939.695 572.320 1940.210 572.460 ;
        RECT 1939.890 572.260 1940.210 572.320 ;
        RECT 1939.890 524.520 1940.210 524.580 ;
        RECT 1939.695 524.380 1940.210 524.520 ;
        RECT 1939.890 524.320 1940.210 524.380 ;
        RECT 1939.890 475.900 1940.210 475.960 ;
        RECT 1939.695 475.760 1940.210 475.900 ;
        RECT 1939.890 475.700 1940.210 475.760 ;
        RECT 1939.890 427.960 1940.210 428.020 ;
        RECT 1939.695 427.820 1940.210 427.960 ;
        RECT 1939.890 427.760 1940.210 427.820 ;
        RECT 1939.890 379.340 1940.210 379.400 ;
        RECT 1940.810 379.340 1941.130 379.400 ;
        RECT 1939.890 379.200 1941.130 379.340 ;
        RECT 1939.890 379.140 1940.210 379.200 ;
        RECT 1940.810 379.140 1941.130 379.200 ;
        RECT 1939.890 331.060 1940.210 331.120 ;
        RECT 1939.695 330.920 1940.210 331.060 ;
        RECT 1939.890 330.860 1940.210 330.920 ;
        RECT 1939.905 283.120 1940.195 283.165 ;
        RECT 1940.350 283.120 1940.670 283.180 ;
        RECT 1939.905 282.980 1940.670 283.120 ;
        RECT 1939.905 282.935 1940.195 282.980 ;
        RECT 1940.350 282.920 1940.670 282.980 ;
        RECT 1939.430 241.640 1939.750 241.700 ;
        RECT 1940.350 241.640 1940.670 241.700 ;
        RECT 1939.430 241.500 1940.670 241.640 ;
        RECT 1939.430 241.440 1939.750 241.500 ;
        RECT 1940.350 241.440 1940.670 241.500 ;
        RECT 1939.430 234.500 1939.750 234.560 ;
        RECT 1939.235 234.360 1939.750 234.500 ;
        RECT 1939.430 234.300 1939.750 234.360 ;
        RECT 1939.430 186.560 1939.750 186.620 ;
        RECT 1939.235 186.420 1939.750 186.560 ;
        RECT 1939.430 186.360 1939.750 186.420 ;
        RECT 1938.985 138.960 1939.275 139.005 ;
        RECT 1939.430 138.960 1939.750 139.020 ;
        RECT 1938.985 138.820 1939.750 138.960 ;
        RECT 1938.985 138.775 1939.275 138.820 ;
        RECT 1939.430 138.760 1939.750 138.820 ;
        RECT 1938.970 138.280 1939.290 138.340 ;
        RECT 1938.775 138.140 1939.290 138.280 ;
        RECT 1938.970 138.080 1939.290 138.140 ;
        RECT 1939.430 48.520 1939.750 48.580 ;
        RECT 1940.350 48.520 1940.670 48.580 ;
        RECT 1939.430 48.380 1940.670 48.520 ;
        RECT 1939.430 48.320 1939.750 48.380 ;
        RECT 1940.350 48.320 1940.670 48.380 ;
        RECT 1542.910 32.540 1543.230 32.600 ;
        RECT 1939.430 32.540 1939.750 32.600 ;
        RECT 1542.910 32.400 1939.750 32.540 ;
        RECT 1542.910 32.340 1543.230 32.400 ;
        RECT 1939.430 32.340 1939.750 32.400 ;
      LAYER via ;
        RECT 1939.460 1593.620 1939.720 1593.880 ;
        RECT 1939.920 1593.620 1940.180 1593.880 ;
        RECT 1939.460 1586.820 1939.720 1587.080 ;
        RECT 1939.460 1538.880 1939.720 1539.140 ;
        RECT 1939.460 1524.260 1939.720 1524.520 ;
        RECT 1939.920 1490.600 1940.180 1490.860 ;
        RECT 1939.920 1463.060 1940.180 1463.320 ;
        RECT 1939.920 1462.380 1940.180 1462.640 ;
        RECT 1939.920 1400.500 1940.180 1400.760 ;
        RECT 1940.380 1400.500 1940.640 1400.760 ;
        RECT 1939.920 814.000 1940.180 814.260 ;
        RECT 1939.920 789.860 1940.180 790.120 ;
        RECT 1939.920 627.680 1940.180 627.940 ;
        RECT 1940.380 627.680 1940.640 627.940 ;
        RECT 1939.920 593.000 1940.180 593.260 ;
        RECT 1940.380 593.000 1940.640 593.260 ;
        RECT 1939.920 572.260 1940.180 572.520 ;
        RECT 1939.920 524.320 1940.180 524.580 ;
        RECT 1939.920 475.700 1940.180 475.960 ;
        RECT 1939.920 427.760 1940.180 428.020 ;
        RECT 1939.920 379.140 1940.180 379.400 ;
        RECT 1940.840 379.140 1941.100 379.400 ;
        RECT 1939.920 330.860 1940.180 331.120 ;
        RECT 1940.380 282.920 1940.640 283.180 ;
        RECT 1939.460 241.440 1939.720 241.700 ;
        RECT 1940.380 241.440 1940.640 241.700 ;
        RECT 1939.460 234.300 1939.720 234.560 ;
        RECT 1939.460 186.360 1939.720 186.620 ;
        RECT 1939.460 138.760 1939.720 139.020 ;
        RECT 1939.000 138.080 1939.260 138.340 ;
        RECT 1939.460 48.320 1939.720 48.580 ;
        RECT 1940.380 48.320 1940.640 48.580 ;
        RECT 1542.940 32.340 1543.200 32.600 ;
        RECT 1939.460 32.340 1939.720 32.600 ;
      LAYER met2 ;
        RECT 1942.600 1700.410 1942.880 1702.400 ;
        RECT 1940.900 1700.270 1942.880 1700.410 ;
        RECT 1940.900 1656.210 1941.040 1700.270 ;
        RECT 1942.600 1700.000 1942.880 1700.270 ;
        RECT 1939.980 1656.070 1941.040 1656.210 ;
        RECT 1939.980 1593.910 1940.120 1656.070 ;
        RECT 1939.460 1593.590 1939.720 1593.910 ;
        RECT 1939.920 1593.590 1940.180 1593.910 ;
        RECT 1939.520 1587.110 1939.660 1593.590 ;
        RECT 1939.460 1586.790 1939.720 1587.110 ;
        RECT 1939.460 1538.850 1939.720 1539.170 ;
        RECT 1939.520 1524.550 1939.660 1538.850 ;
        RECT 1939.460 1524.230 1939.720 1524.550 ;
        RECT 1939.920 1490.570 1940.180 1490.890 ;
        RECT 1939.980 1463.350 1940.120 1490.570 ;
        RECT 1939.920 1463.030 1940.180 1463.350 ;
        RECT 1939.920 1462.350 1940.180 1462.670 ;
        RECT 1939.980 1400.790 1940.120 1462.350 ;
        RECT 1939.920 1400.470 1940.180 1400.790 ;
        RECT 1940.380 1400.470 1940.640 1400.790 ;
        RECT 1940.440 1365.850 1940.580 1400.470 ;
        RECT 1939.980 1365.710 1940.580 1365.850 ;
        RECT 1939.980 1269.970 1940.120 1365.710 ;
        RECT 1939.520 1269.830 1940.120 1269.970 ;
        RECT 1939.520 1269.290 1939.660 1269.830 ;
        RECT 1939.520 1269.150 1940.120 1269.290 ;
        RECT 1939.980 883.730 1940.120 1269.150 ;
        RECT 1939.520 883.590 1940.120 883.730 ;
        RECT 1939.520 883.050 1939.660 883.590 ;
        RECT 1939.520 882.910 1940.120 883.050 ;
        RECT 1939.980 814.290 1940.120 882.910 ;
        RECT 1939.920 813.970 1940.180 814.290 ;
        RECT 1939.920 789.830 1940.180 790.150 ;
        RECT 1939.980 690.610 1940.120 789.830 ;
        RECT 1939.520 690.470 1940.120 690.610 ;
        RECT 1939.520 688.570 1939.660 690.470 ;
        RECT 1939.520 688.430 1940.120 688.570 ;
        RECT 1939.980 627.970 1940.120 688.430 ;
        RECT 1939.920 627.650 1940.180 627.970 ;
        RECT 1940.380 627.650 1940.640 627.970 ;
        RECT 1940.440 593.290 1940.580 627.650 ;
        RECT 1939.920 592.970 1940.180 593.290 ;
        RECT 1940.380 592.970 1940.640 593.290 ;
        RECT 1939.980 572.550 1940.120 592.970 ;
        RECT 1939.920 572.230 1940.180 572.550 ;
        RECT 1939.920 524.290 1940.180 524.610 ;
        RECT 1939.980 475.990 1940.120 524.290 ;
        RECT 1939.920 475.670 1940.180 475.990 ;
        RECT 1939.920 427.730 1940.180 428.050 ;
        RECT 1939.980 379.430 1940.120 427.730 ;
        RECT 1939.920 379.110 1940.180 379.430 ;
        RECT 1940.840 379.110 1941.100 379.430 ;
        RECT 1940.900 331.685 1941.040 379.110 ;
        RECT 1939.910 331.315 1940.190 331.685 ;
        RECT 1940.830 331.315 1941.110 331.685 ;
        RECT 1939.980 331.150 1940.120 331.315 ;
        RECT 1939.920 330.830 1940.180 331.150 ;
        RECT 1940.380 282.890 1940.640 283.210 ;
        RECT 1940.440 241.730 1940.580 282.890 ;
        RECT 1939.460 241.410 1939.720 241.730 ;
        RECT 1940.380 241.410 1940.640 241.730 ;
        RECT 1939.520 234.590 1939.660 241.410 ;
        RECT 1939.460 234.270 1939.720 234.590 ;
        RECT 1939.460 186.330 1939.720 186.650 ;
        RECT 1939.520 139.050 1939.660 186.330 ;
        RECT 1939.460 138.730 1939.720 139.050 ;
        RECT 1939.000 138.050 1939.260 138.370 ;
        RECT 1939.060 95.610 1939.200 138.050 ;
        RECT 1939.060 95.470 1940.580 95.610 ;
        RECT 1940.440 48.610 1940.580 95.470 ;
        RECT 1939.460 48.290 1939.720 48.610 ;
        RECT 1940.380 48.290 1940.640 48.610 ;
        RECT 1939.520 32.630 1939.660 48.290 ;
        RECT 1542.940 32.310 1543.200 32.630 ;
        RECT 1939.460 32.310 1939.720 32.630 ;
        RECT 1543.000 2.400 1543.140 32.310 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
      LAYER via2 ;
        RECT 1939.910 331.360 1940.190 331.640 ;
        RECT 1940.830 331.360 1941.110 331.640 ;
      LAYER met3 ;
        RECT 1939.885 331.650 1940.215 331.665 ;
        RECT 1940.805 331.650 1941.135 331.665 ;
        RECT 1939.885 331.350 1941.135 331.650 ;
        RECT 1939.885 331.335 1940.215 331.350 ;
        RECT 1940.805 331.335 1941.135 331.350 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1560.850 32.880 1561.170 32.940 ;
        RECT 1946.790 32.880 1947.110 32.940 ;
        RECT 1560.850 32.740 1947.110 32.880 ;
        RECT 1560.850 32.680 1561.170 32.740 ;
        RECT 1946.790 32.680 1947.110 32.740 ;
      LAYER via ;
        RECT 1560.880 32.680 1561.140 32.940 ;
        RECT 1946.820 32.680 1947.080 32.940 ;
      LAYER met2 ;
        RECT 1951.800 1700.410 1952.080 1702.400 ;
        RECT 1949.180 1700.270 1952.080 1700.410 ;
        RECT 1949.180 1678.650 1949.320 1700.270 ;
        RECT 1951.800 1700.000 1952.080 1700.270 ;
        RECT 1946.880 1678.510 1949.320 1678.650 ;
        RECT 1946.880 32.970 1947.020 1678.510 ;
        RECT 1560.880 32.650 1561.140 32.970 ;
        RECT 1946.820 32.650 1947.080 32.970 ;
        RECT 1560.940 2.400 1561.080 32.650 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1578.790 27.440 1579.110 27.500 ;
        RECT 1959.670 27.440 1959.990 27.500 ;
        RECT 1578.790 27.300 1959.990 27.440 ;
        RECT 1578.790 27.240 1579.110 27.300 ;
        RECT 1959.670 27.240 1959.990 27.300 ;
      LAYER via ;
        RECT 1578.820 27.240 1579.080 27.500 ;
        RECT 1959.700 27.240 1959.960 27.500 ;
      LAYER met2 ;
        RECT 1961.000 1700.410 1961.280 1702.400 ;
        RECT 1959.760 1700.270 1961.280 1700.410 ;
        RECT 1959.760 27.530 1959.900 1700.270 ;
        RECT 1961.000 1700.000 1961.280 1700.270 ;
        RECT 1578.820 27.210 1579.080 27.530 ;
        RECT 1959.700 27.210 1959.960 27.530 ;
        RECT 1578.880 2.400 1579.020 27.210 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1596.270 22.680 1596.590 22.740 ;
        RECT 1967.490 22.680 1967.810 22.740 ;
        RECT 1596.270 22.540 1967.810 22.680 ;
        RECT 1596.270 22.480 1596.590 22.540 ;
        RECT 1967.490 22.480 1967.810 22.540 ;
      LAYER via ;
        RECT 1596.300 22.480 1596.560 22.740 ;
        RECT 1967.520 22.480 1967.780 22.740 ;
      LAYER met2 ;
        RECT 1970.200 1700.410 1970.480 1702.400 ;
        RECT 1967.580 1700.270 1970.480 1700.410 ;
        RECT 1967.580 22.770 1967.720 1700.270 ;
        RECT 1970.200 1700.000 1970.480 1700.270 ;
        RECT 1596.300 22.450 1596.560 22.770 ;
        RECT 1967.520 22.450 1967.780 22.770 ;
        RECT 1596.360 2.400 1596.500 22.450 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1614.210 22.340 1614.530 22.400 ;
        RECT 1974.390 22.340 1974.710 22.400 ;
        RECT 1614.210 22.200 1974.710 22.340 ;
        RECT 1614.210 22.140 1614.530 22.200 ;
        RECT 1974.390 22.140 1974.710 22.200 ;
      LAYER via ;
        RECT 1614.240 22.140 1614.500 22.400 ;
        RECT 1974.420 22.140 1974.680 22.400 ;
      LAYER met2 ;
        RECT 1979.400 1700.410 1979.680 1702.400 ;
        RECT 1976.780 1700.270 1979.680 1700.410 ;
        RECT 1976.780 1678.650 1976.920 1700.270 ;
        RECT 1979.400 1700.000 1979.680 1700.270 ;
        RECT 1974.480 1678.510 1976.920 1678.650 ;
        RECT 1974.480 22.430 1974.620 1678.510 ;
        RECT 1614.240 22.110 1614.500 22.430 ;
        RECT 1974.420 22.110 1974.680 22.430 ;
        RECT 1614.300 2.400 1614.440 22.110 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1632.150 22.000 1632.470 22.060 ;
        RECT 1987.270 22.000 1987.590 22.060 ;
        RECT 1632.150 21.860 1987.590 22.000 ;
        RECT 1632.150 21.800 1632.470 21.860 ;
        RECT 1987.270 21.800 1987.590 21.860 ;
      LAYER via ;
        RECT 1632.180 21.800 1632.440 22.060 ;
        RECT 1987.300 21.800 1987.560 22.060 ;
      LAYER met2 ;
        RECT 1988.600 1700.410 1988.880 1702.400 ;
        RECT 1987.360 1700.270 1988.880 1700.410 ;
        RECT 1987.360 22.090 1987.500 1700.270 ;
        RECT 1988.600 1700.000 1988.880 1700.270 ;
        RECT 1632.180 21.770 1632.440 22.090 ;
        RECT 1987.300 21.770 1987.560 22.090 ;
        RECT 1632.240 2.400 1632.380 21.770 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1650.090 21.660 1650.410 21.720 ;
        RECT 1995.090 21.660 1995.410 21.720 ;
        RECT 1650.090 21.520 1995.410 21.660 ;
        RECT 1650.090 21.460 1650.410 21.520 ;
        RECT 1995.090 21.460 1995.410 21.520 ;
      LAYER via ;
        RECT 1650.120 21.460 1650.380 21.720 ;
        RECT 1995.120 21.460 1995.380 21.720 ;
      LAYER met2 ;
        RECT 1997.800 1700.410 1998.080 1702.400 ;
        RECT 1995.180 1700.270 1998.080 1700.410 ;
        RECT 1995.180 21.750 1995.320 1700.270 ;
        RECT 1997.800 1700.000 1998.080 1700.270 ;
        RECT 1650.120 21.430 1650.380 21.750 ;
        RECT 1995.120 21.430 1995.380 21.750 ;
        RECT 1650.180 2.400 1650.320 21.430 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2002.525 1352.605 2002.695 1400.715 ;
        RECT 2002.525 1256.045 2002.695 1304.155 ;
        RECT 2002.525 737.885 2002.695 765.935 ;
        RECT 2001.605 572.645 2001.775 620.755 ;
        RECT 2001.605 386.325 2001.775 434.775 ;
        RECT 2002.065 241.825 2002.235 255.935 ;
        RECT 2003.445 145.265 2003.615 159.035 ;
        RECT 2002.985 89.845 2003.155 137.955 ;
        RECT 2002.065 41.565 2002.235 89.335 ;
      LAYER mcon ;
        RECT 2002.525 1400.545 2002.695 1400.715 ;
        RECT 2002.525 1303.985 2002.695 1304.155 ;
        RECT 2002.525 765.765 2002.695 765.935 ;
        RECT 2001.605 620.585 2001.775 620.755 ;
        RECT 2001.605 434.605 2001.775 434.775 ;
        RECT 2002.065 255.765 2002.235 255.935 ;
        RECT 2003.445 158.865 2003.615 159.035 ;
        RECT 2002.985 137.785 2003.155 137.955 ;
        RECT 2002.065 89.165 2002.235 89.335 ;
      LAYER met1 ;
        RECT 2001.990 1607.760 2002.310 1607.820 ;
        RECT 2002.910 1607.760 2003.230 1607.820 ;
        RECT 2001.990 1607.620 2003.230 1607.760 ;
        RECT 2001.990 1607.560 2002.310 1607.620 ;
        RECT 2002.910 1607.560 2003.230 1607.620 ;
        RECT 2001.530 1545.880 2001.850 1545.940 ;
        RECT 2001.990 1545.880 2002.310 1545.940 ;
        RECT 2001.530 1545.740 2002.310 1545.880 ;
        RECT 2001.530 1545.680 2001.850 1545.740 ;
        RECT 2001.990 1545.680 2002.310 1545.740 ;
        RECT 2001.990 1511.340 2002.310 1511.600 ;
        RECT 2002.080 1510.520 2002.220 1511.340 ;
        RECT 2002.450 1510.520 2002.770 1510.580 ;
        RECT 2002.080 1510.380 2002.770 1510.520 ;
        RECT 2002.450 1510.320 2002.770 1510.380 ;
        RECT 2002.450 1490.460 2002.770 1490.520 ;
        RECT 2002.910 1490.460 2003.230 1490.520 ;
        RECT 2002.450 1490.320 2003.230 1490.460 ;
        RECT 2002.450 1490.260 2002.770 1490.320 ;
        RECT 2002.910 1490.260 2003.230 1490.320 ;
        RECT 2002.450 1400.700 2002.770 1400.760 ;
        RECT 2002.255 1400.560 2002.770 1400.700 ;
        RECT 2002.450 1400.500 2002.770 1400.560 ;
        RECT 2002.465 1352.760 2002.755 1352.805 ;
        RECT 2002.910 1352.760 2003.230 1352.820 ;
        RECT 2002.465 1352.620 2003.230 1352.760 ;
        RECT 2002.465 1352.575 2002.755 1352.620 ;
        RECT 2002.910 1352.560 2003.230 1352.620 ;
        RECT 2002.450 1304.140 2002.770 1304.200 ;
        RECT 2002.255 1304.000 2002.770 1304.140 ;
        RECT 2002.450 1303.940 2002.770 1304.000 ;
        RECT 2002.465 1256.200 2002.755 1256.245 ;
        RECT 2002.910 1256.200 2003.230 1256.260 ;
        RECT 2002.465 1256.060 2003.230 1256.200 ;
        RECT 2002.465 1256.015 2002.755 1256.060 ;
        RECT 2002.910 1256.000 2003.230 1256.060 ;
        RECT 2001.530 1159.300 2001.850 1159.360 ;
        RECT 2002.910 1159.300 2003.230 1159.360 ;
        RECT 2001.530 1159.160 2003.230 1159.300 ;
        RECT 2001.530 1159.100 2001.850 1159.160 ;
        RECT 2002.910 1159.100 2003.230 1159.160 ;
        RECT 2001.530 1062.740 2001.850 1062.800 ;
        RECT 2002.910 1062.740 2003.230 1062.800 ;
        RECT 2001.530 1062.600 2003.230 1062.740 ;
        RECT 2001.530 1062.540 2001.850 1062.600 ;
        RECT 2002.910 1062.540 2003.230 1062.600 ;
        RECT 2001.530 966.180 2001.850 966.240 ;
        RECT 2002.910 966.180 2003.230 966.240 ;
        RECT 2001.530 966.040 2003.230 966.180 ;
        RECT 2001.530 965.980 2001.850 966.040 ;
        RECT 2002.910 965.980 2003.230 966.040 ;
        RECT 2001.990 883.220 2002.310 883.280 ;
        RECT 2002.910 883.220 2003.230 883.280 ;
        RECT 2001.990 883.080 2003.230 883.220 ;
        RECT 2001.990 883.020 2002.310 883.080 ;
        RECT 2002.910 883.020 2003.230 883.080 ;
        RECT 2001.530 821.340 2001.850 821.400 ;
        RECT 2001.990 821.340 2002.310 821.400 ;
        RECT 2001.530 821.200 2002.310 821.340 ;
        RECT 2001.530 821.140 2001.850 821.200 ;
        RECT 2001.990 821.140 2002.310 821.200 ;
        RECT 2002.450 765.920 2002.770 765.980 ;
        RECT 2002.255 765.780 2002.770 765.920 ;
        RECT 2002.450 765.720 2002.770 765.780 ;
        RECT 2002.450 738.040 2002.770 738.100 ;
        RECT 2002.255 737.900 2002.770 738.040 ;
        RECT 2002.450 737.840 2002.770 737.900 ;
        RECT 2001.990 717.640 2002.310 717.700 ;
        RECT 2002.450 717.640 2002.770 717.700 ;
        RECT 2001.990 717.500 2002.770 717.640 ;
        RECT 2001.990 717.440 2002.310 717.500 ;
        RECT 2002.450 717.440 2002.770 717.500 ;
        RECT 2001.990 641.620 2002.310 641.880 ;
        RECT 2002.080 641.480 2002.220 641.620 ;
        RECT 2002.450 641.480 2002.770 641.540 ;
        RECT 2002.080 641.340 2002.770 641.480 ;
        RECT 2002.450 641.280 2002.770 641.340 ;
        RECT 2001.545 620.740 2001.835 620.785 ;
        RECT 2002.450 620.740 2002.770 620.800 ;
        RECT 2001.545 620.600 2002.770 620.740 ;
        RECT 2001.545 620.555 2001.835 620.600 ;
        RECT 2002.450 620.540 2002.770 620.600 ;
        RECT 2001.530 572.800 2001.850 572.860 ;
        RECT 2001.335 572.660 2001.850 572.800 ;
        RECT 2001.530 572.600 2001.850 572.660 ;
        RECT 2001.545 434.760 2001.835 434.805 ;
        RECT 2001.990 434.760 2002.310 434.820 ;
        RECT 2001.545 434.620 2002.310 434.760 ;
        RECT 2001.545 434.575 2001.835 434.620 ;
        RECT 2001.990 434.560 2002.310 434.620 ;
        RECT 2001.530 386.480 2001.850 386.540 ;
        RECT 2001.335 386.340 2001.850 386.480 ;
        RECT 2001.530 386.280 2001.850 386.340 ;
        RECT 2002.005 255.920 2002.295 255.965 ;
        RECT 2002.450 255.920 2002.770 255.980 ;
        RECT 2002.005 255.780 2002.770 255.920 ;
        RECT 2002.005 255.735 2002.295 255.780 ;
        RECT 2002.450 255.720 2002.770 255.780 ;
        RECT 2001.990 241.980 2002.310 242.040 ;
        RECT 2001.795 241.840 2002.310 241.980 ;
        RECT 2001.990 241.780 2002.310 241.840 ;
        RECT 2001.990 241.300 2002.310 241.360 ;
        RECT 2003.830 241.300 2004.150 241.360 ;
        RECT 2001.990 241.160 2004.150 241.300 ;
        RECT 2001.990 241.100 2002.310 241.160 ;
        RECT 2003.830 241.100 2004.150 241.160 ;
        RECT 2003.370 159.020 2003.690 159.080 ;
        RECT 2003.175 158.880 2003.690 159.020 ;
        RECT 2003.370 158.820 2003.690 158.880 ;
        RECT 2003.370 145.420 2003.690 145.480 ;
        RECT 2003.175 145.280 2003.690 145.420 ;
        RECT 2003.370 145.220 2003.690 145.280 ;
        RECT 2002.910 137.940 2003.230 138.000 ;
        RECT 2002.715 137.800 2003.230 137.940 ;
        RECT 2002.910 137.740 2003.230 137.800 ;
        RECT 2002.910 90.000 2003.230 90.060 ;
        RECT 2002.715 89.860 2003.230 90.000 ;
        RECT 2002.910 89.800 2003.230 89.860 ;
        RECT 2002.005 89.320 2002.295 89.365 ;
        RECT 2002.910 89.320 2003.230 89.380 ;
        RECT 2002.005 89.180 2003.230 89.320 ;
        RECT 2002.005 89.135 2002.295 89.180 ;
        RECT 2002.910 89.120 2003.230 89.180 ;
        RECT 2001.990 41.720 2002.310 41.780 ;
        RECT 2001.795 41.580 2002.310 41.720 ;
        RECT 2001.990 41.520 2002.310 41.580 ;
        RECT 1668.030 21.320 1668.350 21.380 ;
        RECT 2001.990 21.320 2002.310 21.380 ;
        RECT 1668.030 21.180 2002.310 21.320 ;
        RECT 1668.030 21.120 1668.350 21.180 ;
        RECT 2001.990 21.120 2002.310 21.180 ;
      LAYER via ;
        RECT 2002.020 1607.560 2002.280 1607.820 ;
        RECT 2002.940 1607.560 2003.200 1607.820 ;
        RECT 2001.560 1545.680 2001.820 1545.940 ;
        RECT 2002.020 1545.680 2002.280 1545.940 ;
        RECT 2002.020 1511.340 2002.280 1511.600 ;
        RECT 2002.480 1510.320 2002.740 1510.580 ;
        RECT 2002.480 1490.260 2002.740 1490.520 ;
        RECT 2002.940 1490.260 2003.200 1490.520 ;
        RECT 2002.480 1400.500 2002.740 1400.760 ;
        RECT 2002.940 1352.560 2003.200 1352.820 ;
        RECT 2002.480 1303.940 2002.740 1304.200 ;
        RECT 2002.940 1256.000 2003.200 1256.260 ;
        RECT 2001.560 1159.100 2001.820 1159.360 ;
        RECT 2002.940 1159.100 2003.200 1159.360 ;
        RECT 2001.560 1062.540 2001.820 1062.800 ;
        RECT 2002.940 1062.540 2003.200 1062.800 ;
        RECT 2001.560 965.980 2001.820 966.240 ;
        RECT 2002.940 965.980 2003.200 966.240 ;
        RECT 2002.020 883.020 2002.280 883.280 ;
        RECT 2002.940 883.020 2003.200 883.280 ;
        RECT 2001.560 821.140 2001.820 821.400 ;
        RECT 2002.020 821.140 2002.280 821.400 ;
        RECT 2002.480 765.720 2002.740 765.980 ;
        RECT 2002.480 737.840 2002.740 738.100 ;
        RECT 2002.020 717.440 2002.280 717.700 ;
        RECT 2002.480 717.440 2002.740 717.700 ;
        RECT 2002.020 641.620 2002.280 641.880 ;
        RECT 2002.480 641.280 2002.740 641.540 ;
        RECT 2002.480 620.540 2002.740 620.800 ;
        RECT 2001.560 572.600 2001.820 572.860 ;
        RECT 2002.020 434.560 2002.280 434.820 ;
        RECT 2001.560 386.280 2001.820 386.540 ;
        RECT 2002.480 255.720 2002.740 255.980 ;
        RECT 2002.020 241.780 2002.280 242.040 ;
        RECT 2002.020 241.100 2002.280 241.360 ;
        RECT 2003.860 241.100 2004.120 241.360 ;
        RECT 2003.400 158.820 2003.660 159.080 ;
        RECT 2003.400 145.220 2003.660 145.480 ;
        RECT 2002.940 137.740 2003.200 138.000 ;
        RECT 2002.940 89.800 2003.200 90.060 ;
        RECT 2002.940 89.120 2003.200 89.380 ;
        RECT 2002.020 41.520 2002.280 41.780 ;
        RECT 1668.060 21.120 1668.320 21.380 ;
        RECT 2002.020 21.120 2002.280 21.380 ;
      LAYER met2 ;
        RECT 2007.000 1700.410 2007.280 1702.400 ;
        RECT 2004.380 1700.270 2007.280 1700.410 ;
        RECT 2004.380 1677.970 2004.520 1700.270 ;
        RECT 2007.000 1700.000 2007.280 1700.270 ;
        RECT 2003.000 1677.830 2004.520 1677.970 ;
        RECT 2003.000 1607.850 2003.140 1677.830 ;
        RECT 2002.020 1607.530 2002.280 1607.850 ;
        RECT 2002.940 1607.530 2003.200 1607.850 ;
        RECT 2002.080 1559.650 2002.220 1607.530 ;
        RECT 2001.620 1559.510 2002.220 1559.650 ;
        RECT 2001.620 1545.970 2001.760 1559.510 ;
        RECT 2001.560 1545.650 2001.820 1545.970 ;
        RECT 2002.020 1545.650 2002.280 1545.970 ;
        RECT 2002.080 1511.630 2002.220 1545.650 ;
        RECT 2002.020 1511.310 2002.280 1511.630 ;
        RECT 2002.480 1510.290 2002.740 1510.610 ;
        RECT 2002.540 1490.550 2002.680 1510.290 ;
        RECT 2002.480 1490.230 2002.740 1490.550 ;
        RECT 2002.940 1490.230 2003.200 1490.550 ;
        RECT 2003.000 1401.210 2003.140 1490.230 ;
        RECT 2002.540 1401.070 2003.140 1401.210 ;
        RECT 2002.540 1400.790 2002.680 1401.070 ;
        RECT 2002.480 1400.470 2002.740 1400.790 ;
        RECT 2002.940 1352.530 2003.200 1352.850 ;
        RECT 2003.000 1317.570 2003.140 1352.530 ;
        RECT 2002.540 1317.430 2003.140 1317.570 ;
        RECT 2002.540 1304.230 2002.680 1317.430 ;
        RECT 2002.480 1303.910 2002.740 1304.230 ;
        RECT 2002.940 1255.970 2003.200 1256.290 ;
        RECT 2003.000 1221.010 2003.140 1255.970 ;
        RECT 2002.540 1220.870 2003.140 1221.010 ;
        RECT 2002.540 1207.525 2002.680 1220.870 ;
        RECT 2001.550 1207.155 2001.830 1207.525 ;
        RECT 2002.470 1207.155 2002.750 1207.525 ;
        RECT 2001.620 1159.390 2001.760 1207.155 ;
        RECT 2001.560 1159.070 2001.820 1159.390 ;
        RECT 2002.940 1159.070 2003.200 1159.390 ;
        RECT 2003.000 1124.450 2003.140 1159.070 ;
        RECT 2002.540 1124.310 2003.140 1124.450 ;
        RECT 2002.540 1110.965 2002.680 1124.310 ;
        RECT 2001.550 1110.595 2001.830 1110.965 ;
        RECT 2002.470 1110.595 2002.750 1110.965 ;
        RECT 2001.620 1062.830 2001.760 1110.595 ;
        RECT 2001.560 1062.510 2001.820 1062.830 ;
        RECT 2002.940 1062.510 2003.200 1062.830 ;
        RECT 2003.000 1027.890 2003.140 1062.510 ;
        RECT 2002.540 1027.750 2003.140 1027.890 ;
        RECT 2002.540 1014.405 2002.680 1027.750 ;
        RECT 2001.550 1014.035 2001.830 1014.405 ;
        RECT 2002.470 1014.035 2002.750 1014.405 ;
        RECT 2001.620 966.270 2001.760 1014.035 ;
        RECT 2001.560 965.950 2001.820 966.270 ;
        RECT 2002.940 965.950 2003.200 966.270 ;
        RECT 2003.000 931.330 2003.140 965.950 ;
        RECT 2002.540 931.190 2003.140 931.330 ;
        RECT 2002.540 883.730 2002.680 931.190 ;
        RECT 2002.080 883.590 2002.680 883.730 ;
        RECT 2002.080 883.310 2002.220 883.590 ;
        RECT 2002.020 882.990 2002.280 883.310 ;
        RECT 2002.940 882.990 2003.200 883.310 ;
        RECT 2003.000 869.450 2003.140 882.990 ;
        RECT 2002.080 869.310 2003.140 869.450 ;
        RECT 2002.080 821.430 2002.220 869.310 ;
        RECT 2001.560 821.110 2001.820 821.430 ;
        RECT 2002.020 821.110 2002.280 821.430 ;
        RECT 2001.620 773.685 2001.760 821.110 ;
        RECT 2001.550 773.315 2001.830 773.685 ;
        RECT 2002.470 772.635 2002.750 773.005 ;
        RECT 2002.540 766.010 2002.680 772.635 ;
        RECT 2002.480 765.690 2002.740 766.010 ;
        RECT 2002.480 737.810 2002.740 738.130 ;
        RECT 2002.540 717.730 2002.680 737.810 ;
        RECT 2002.020 717.410 2002.280 717.730 ;
        RECT 2002.480 717.410 2002.740 717.730 ;
        RECT 2002.080 641.910 2002.220 717.410 ;
        RECT 2002.020 641.590 2002.280 641.910 ;
        RECT 2002.480 641.250 2002.740 641.570 ;
        RECT 2002.540 620.830 2002.680 641.250 ;
        RECT 2002.480 620.510 2002.740 620.830 ;
        RECT 2001.560 572.570 2001.820 572.890 ;
        RECT 2001.620 531.605 2001.760 572.570 ;
        RECT 2001.550 531.235 2001.830 531.605 ;
        RECT 2002.470 531.235 2002.750 531.605 ;
        RECT 2002.540 507.010 2002.680 531.235 ;
        RECT 2001.620 506.870 2002.680 507.010 ;
        RECT 2001.620 483.325 2001.760 506.870 ;
        RECT 2001.550 482.955 2001.830 483.325 ;
        RECT 2002.930 482.955 2003.210 483.325 ;
        RECT 2003.000 448.530 2003.140 482.955 ;
        RECT 2002.080 448.390 2003.140 448.530 ;
        RECT 2002.080 434.850 2002.220 448.390 ;
        RECT 2002.020 434.530 2002.280 434.850 ;
        RECT 2001.560 386.250 2001.820 386.570 ;
        RECT 2001.620 351.970 2001.760 386.250 ;
        RECT 2001.620 351.830 2002.680 351.970 ;
        RECT 2002.540 256.010 2002.680 351.830 ;
        RECT 2002.480 255.690 2002.740 256.010 ;
        RECT 2002.020 241.750 2002.280 242.070 ;
        RECT 2002.080 241.390 2002.220 241.750 ;
        RECT 2002.020 241.070 2002.280 241.390 ;
        RECT 2003.860 241.070 2004.120 241.390 ;
        RECT 2003.920 193.530 2004.060 241.070 ;
        RECT 2003.460 193.390 2004.060 193.530 ;
        RECT 2003.460 159.110 2003.600 193.390 ;
        RECT 2003.400 158.790 2003.660 159.110 ;
        RECT 2003.400 145.250 2003.660 145.510 ;
        RECT 2003.000 145.190 2003.660 145.250 ;
        RECT 2003.000 145.110 2003.600 145.190 ;
        RECT 2003.000 138.030 2003.140 145.110 ;
        RECT 2002.940 137.710 2003.200 138.030 ;
        RECT 2002.940 89.770 2003.200 90.090 ;
        RECT 2003.000 89.410 2003.140 89.770 ;
        RECT 2002.940 89.090 2003.200 89.410 ;
        RECT 2002.020 41.490 2002.280 41.810 ;
        RECT 2002.080 21.410 2002.220 41.490 ;
        RECT 1668.060 21.090 1668.320 21.410 ;
        RECT 2002.020 21.090 2002.280 21.410 ;
        RECT 1668.120 2.400 1668.260 21.090 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
      LAYER via2 ;
        RECT 2001.550 1207.200 2001.830 1207.480 ;
        RECT 2002.470 1207.200 2002.750 1207.480 ;
        RECT 2001.550 1110.640 2001.830 1110.920 ;
        RECT 2002.470 1110.640 2002.750 1110.920 ;
        RECT 2001.550 1014.080 2001.830 1014.360 ;
        RECT 2002.470 1014.080 2002.750 1014.360 ;
        RECT 2001.550 773.360 2001.830 773.640 ;
        RECT 2002.470 772.680 2002.750 772.960 ;
        RECT 2001.550 531.280 2001.830 531.560 ;
        RECT 2002.470 531.280 2002.750 531.560 ;
        RECT 2001.550 483.000 2001.830 483.280 ;
        RECT 2002.930 483.000 2003.210 483.280 ;
      LAYER met3 ;
        RECT 2001.525 1207.490 2001.855 1207.505 ;
        RECT 2002.445 1207.490 2002.775 1207.505 ;
        RECT 2001.525 1207.190 2002.775 1207.490 ;
        RECT 2001.525 1207.175 2001.855 1207.190 ;
        RECT 2002.445 1207.175 2002.775 1207.190 ;
        RECT 2001.525 1110.930 2001.855 1110.945 ;
        RECT 2002.445 1110.930 2002.775 1110.945 ;
        RECT 2001.525 1110.630 2002.775 1110.930 ;
        RECT 2001.525 1110.615 2001.855 1110.630 ;
        RECT 2002.445 1110.615 2002.775 1110.630 ;
        RECT 2001.525 1014.370 2001.855 1014.385 ;
        RECT 2002.445 1014.370 2002.775 1014.385 ;
        RECT 2001.525 1014.070 2002.775 1014.370 ;
        RECT 2001.525 1014.055 2001.855 1014.070 ;
        RECT 2002.445 1014.055 2002.775 1014.070 ;
        RECT 2001.525 773.650 2001.855 773.665 ;
        RECT 2001.525 773.350 2003.450 773.650 ;
        RECT 2001.525 773.335 2001.855 773.350 ;
        RECT 2002.445 772.970 2002.775 772.985 ;
        RECT 2003.150 772.970 2003.450 773.350 ;
        RECT 2002.445 772.670 2003.450 772.970 ;
        RECT 2002.445 772.655 2002.775 772.670 ;
        RECT 2001.525 531.570 2001.855 531.585 ;
        RECT 2002.445 531.570 2002.775 531.585 ;
        RECT 2001.525 531.270 2002.775 531.570 ;
        RECT 2001.525 531.255 2001.855 531.270 ;
        RECT 2002.445 531.255 2002.775 531.270 ;
        RECT 2001.525 483.290 2001.855 483.305 ;
        RECT 2002.905 483.290 2003.235 483.305 ;
        RECT 2001.525 482.990 2003.235 483.290 ;
        RECT 2001.525 482.975 2001.855 482.990 ;
        RECT 2002.905 482.975 2003.235 482.990 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.510 20.980 1685.830 21.040 ;
        RECT 2015.330 20.980 2015.650 21.040 ;
        RECT 1685.510 20.840 2015.650 20.980 ;
        RECT 1685.510 20.780 1685.830 20.840 ;
        RECT 2015.330 20.780 2015.650 20.840 ;
      LAYER via ;
        RECT 1685.540 20.780 1685.800 21.040 ;
        RECT 2015.360 20.780 2015.620 21.040 ;
      LAYER met2 ;
        RECT 2016.200 1700.410 2016.480 1702.400 ;
        RECT 2015.420 1700.270 2016.480 1700.410 ;
        RECT 2015.420 21.070 2015.560 1700.270 ;
        RECT 2016.200 1700.000 2016.480 1700.270 ;
        RECT 1685.540 20.750 1685.800 21.070 ;
        RECT 2015.360 20.750 2015.620 21.070 ;
        RECT 1685.600 2.400 1685.740 20.750 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.110 66.200 724.430 66.260 ;
        RECT 1518.530 66.200 1518.850 66.260 ;
        RECT 724.110 66.060 1518.850 66.200 ;
        RECT 724.110 66.000 724.430 66.060 ;
        RECT 1518.530 66.000 1518.850 66.060 ;
      LAYER via ;
        RECT 724.140 66.000 724.400 66.260 ;
        RECT 1518.560 66.000 1518.820 66.260 ;
      LAYER met2 ;
        RECT 1520.320 1700.410 1520.600 1702.400 ;
        RECT 1518.620 1700.270 1520.600 1700.410 ;
        RECT 1518.620 66.290 1518.760 1700.270 ;
        RECT 1520.320 1700.000 1520.600 1700.270 ;
        RECT 724.140 65.970 724.400 66.290 ;
        RECT 1518.560 65.970 1518.820 66.290 ;
        RECT 724.200 16.730 724.340 65.970 ;
        RECT 722.360 16.590 724.340 16.730 ;
        RECT 722.360 2.400 722.500 16.590 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.450 23.700 1703.770 23.760 ;
        RECT 2022.690 23.700 2023.010 23.760 ;
        RECT 1703.450 23.560 2023.010 23.700 ;
        RECT 1703.450 23.500 1703.770 23.560 ;
        RECT 2022.690 23.500 2023.010 23.560 ;
      LAYER via ;
        RECT 1703.480 23.500 1703.740 23.760 ;
        RECT 2022.720 23.500 2022.980 23.760 ;
      LAYER met2 ;
        RECT 2025.400 1700.410 2025.680 1702.400 ;
        RECT 2022.780 1700.270 2025.680 1700.410 ;
        RECT 2022.780 23.790 2022.920 1700.270 ;
        RECT 2025.400 1700.000 2025.680 1700.270 ;
        RECT 1703.480 23.470 1703.740 23.790 ;
        RECT 2022.720 23.470 2022.980 23.790 ;
        RECT 1703.540 2.400 1703.680 23.470 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2029.590 1678.140 2029.910 1678.200 ;
        RECT 2033.270 1678.140 2033.590 1678.200 ;
        RECT 2029.590 1678.000 2033.590 1678.140 ;
        RECT 2029.590 1677.940 2029.910 1678.000 ;
        RECT 2033.270 1677.940 2033.590 1678.000 ;
        RECT 1721.390 23.360 1721.710 23.420 ;
        RECT 2029.590 23.360 2029.910 23.420 ;
        RECT 1721.390 23.220 2029.910 23.360 ;
        RECT 1721.390 23.160 1721.710 23.220 ;
        RECT 2029.590 23.160 2029.910 23.220 ;
      LAYER via ;
        RECT 2029.620 1677.940 2029.880 1678.200 ;
        RECT 2033.300 1677.940 2033.560 1678.200 ;
        RECT 1721.420 23.160 1721.680 23.420 ;
        RECT 2029.620 23.160 2029.880 23.420 ;
      LAYER met2 ;
        RECT 2034.600 1700.410 2034.880 1702.400 ;
        RECT 2033.360 1700.270 2034.880 1700.410 ;
        RECT 2033.360 1678.230 2033.500 1700.270 ;
        RECT 2034.600 1700.000 2034.880 1700.270 ;
        RECT 2029.620 1677.910 2029.880 1678.230 ;
        RECT 2033.300 1677.910 2033.560 1678.230 ;
        RECT 2029.680 23.450 2029.820 1677.910 ;
        RECT 1721.420 23.130 1721.680 23.450 ;
        RECT 2029.620 23.130 2029.880 23.450 ;
        RECT 1721.480 2.400 1721.620 23.130 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1739.330 24.380 1739.650 24.440 ;
        RECT 2042.470 24.380 2042.790 24.440 ;
        RECT 1739.330 24.240 2042.790 24.380 ;
        RECT 1739.330 24.180 1739.650 24.240 ;
        RECT 2042.470 24.180 2042.790 24.240 ;
      LAYER via ;
        RECT 1739.360 24.180 1739.620 24.440 ;
        RECT 2042.500 24.180 2042.760 24.440 ;
      LAYER met2 ;
        RECT 2043.800 1700.410 2044.080 1702.400 ;
        RECT 2042.560 1700.270 2044.080 1700.410 ;
        RECT 2042.560 24.470 2042.700 1700.270 ;
        RECT 2043.800 1700.000 2044.080 1700.270 ;
        RECT 1739.360 24.150 1739.620 24.470 ;
        RECT 2042.500 24.150 2042.760 24.470 ;
        RECT 1739.420 2.400 1739.560 24.150 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1756.810 24.040 1757.130 24.100 ;
        RECT 2050.290 24.040 2050.610 24.100 ;
        RECT 1756.810 23.900 2050.610 24.040 ;
        RECT 1756.810 23.840 1757.130 23.900 ;
        RECT 2050.290 23.840 2050.610 23.900 ;
      LAYER via ;
        RECT 1756.840 23.840 1757.100 24.100 ;
        RECT 2050.320 23.840 2050.580 24.100 ;
      LAYER met2 ;
        RECT 2053.000 1700.410 2053.280 1702.400 ;
        RECT 2050.380 1700.270 2053.280 1700.410 ;
        RECT 2050.380 24.130 2050.520 1700.270 ;
        RECT 2053.000 1700.000 2053.280 1700.270 ;
        RECT 1756.840 23.810 1757.100 24.130 ;
        RECT 2050.320 23.810 2050.580 24.130 ;
        RECT 1756.900 2.400 1757.040 23.810 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1774.750 30.160 1775.070 30.220 ;
        RECT 2056.730 30.160 2057.050 30.220 ;
        RECT 1774.750 30.020 2057.050 30.160 ;
        RECT 1774.750 29.960 1775.070 30.020 ;
        RECT 2056.730 29.960 2057.050 30.020 ;
      LAYER via ;
        RECT 1774.780 29.960 1775.040 30.220 ;
        RECT 2056.760 29.960 2057.020 30.220 ;
      LAYER met2 ;
        RECT 2062.200 1700.410 2062.480 1702.400 ;
        RECT 2059.580 1700.270 2062.480 1700.410 ;
        RECT 2059.580 1677.970 2059.720 1700.270 ;
        RECT 2062.200 1700.000 2062.480 1700.270 ;
        RECT 2056.820 1677.830 2059.720 1677.970 ;
        RECT 2056.820 30.250 2056.960 1677.830 ;
        RECT 1774.780 29.930 1775.040 30.250 ;
        RECT 2056.760 29.930 2057.020 30.250 ;
        RECT 1774.840 2.400 1774.980 29.930 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1792.690 24.720 1793.010 24.780 ;
        RECT 2070.530 24.720 2070.850 24.780 ;
        RECT 1792.690 24.580 2070.850 24.720 ;
        RECT 1792.690 24.520 1793.010 24.580 ;
        RECT 2070.530 24.520 2070.850 24.580 ;
      LAYER via ;
        RECT 1792.720 24.520 1792.980 24.780 ;
        RECT 2070.560 24.520 2070.820 24.780 ;
      LAYER met2 ;
        RECT 2071.400 1700.410 2071.680 1702.400 ;
        RECT 2070.620 1700.270 2071.680 1700.410 ;
        RECT 2070.620 24.810 2070.760 1700.270 ;
        RECT 2071.400 1700.000 2071.680 1700.270 ;
        RECT 1792.720 24.490 1792.980 24.810 ;
        RECT 2070.560 24.490 2070.820 24.810 ;
        RECT 1792.780 2.400 1792.920 24.490 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1810.630 29.480 1810.950 29.540 ;
        RECT 2077.890 29.480 2078.210 29.540 ;
        RECT 1810.630 29.340 2078.210 29.480 ;
        RECT 1810.630 29.280 1810.950 29.340 ;
        RECT 2077.890 29.280 2078.210 29.340 ;
      LAYER via ;
        RECT 1810.660 29.280 1810.920 29.540 ;
        RECT 2077.920 29.280 2078.180 29.540 ;
      LAYER met2 ;
        RECT 2080.600 1700.410 2080.880 1702.400 ;
        RECT 2077.980 1700.270 2080.880 1700.410 ;
        RECT 2077.980 29.570 2078.120 1700.270 ;
        RECT 2080.600 1700.000 2080.880 1700.270 ;
        RECT 1810.660 29.250 1810.920 29.570 ;
        RECT 2077.920 29.250 2078.180 29.570 ;
        RECT 1810.720 2.400 1810.860 29.250 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2084.405 1594.005 2084.575 1642.115 ;
        RECT 2084.405 1497.445 2084.575 1545.555 ;
        RECT 2084.405 1352.605 2084.575 1400.715 ;
        RECT 2084.405 1256.045 2084.575 1304.155 ;
        RECT 2084.405 338.045 2084.575 386.155 ;
        RECT 2084.405 241.825 2084.575 289.595 ;
        RECT 2084.405 144.925 2084.575 193.035 ;
        RECT 2084.865 61.285 2085.035 96.475 ;
      LAYER mcon ;
        RECT 2084.405 1641.945 2084.575 1642.115 ;
        RECT 2084.405 1545.385 2084.575 1545.555 ;
        RECT 2084.405 1400.545 2084.575 1400.715 ;
        RECT 2084.405 1303.985 2084.575 1304.155 ;
        RECT 2084.405 385.985 2084.575 386.155 ;
        RECT 2084.405 289.425 2084.575 289.595 ;
        RECT 2084.405 192.865 2084.575 193.035 ;
        RECT 2084.865 96.305 2085.035 96.475 ;
      LAYER met1 ;
        RECT 2083.870 1656.040 2084.190 1656.100 ;
        RECT 2084.790 1656.040 2085.110 1656.100 ;
        RECT 2083.870 1655.900 2085.110 1656.040 ;
        RECT 2083.870 1655.840 2084.190 1655.900 ;
        RECT 2084.790 1655.840 2085.110 1655.900 ;
        RECT 2084.345 1642.100 2084.635 1642.145 ;
        RECT 2084.790 1642.100 2085.110 1642.160 ;
        RECT 2084.345 1641.960 2085.110 1642.100 ;
        RECT 2084.345 1641.915 2084.635 1641.960 ;
        RECT 2084.790 1641.900 2085.110 1641.960 ;
        RECT 2084.330 1594.160 2084.650 1594.220 ;
        RECT 2084.135 1594.020 2084.650 1594.160 ;
        RECT 2084.330 1593.960 2084.650 1594.020 ;
        RECT 2083.870 1559.140 2084.190 1559.200 ;
        RECT 2084.790 1559.140 2085.110 1559.200 ;
        RECT 2083.870 1559.000 2085.110 1559.140 ;
        RECT 2083.870 1558.940 2084.190 1559.000 ;
        RECT 2084.790 1558.940 2085.110 1559.000 ;
        RECT 2084.345 1545.540 2084.635 1545.585 ;
        RECT 2084.790 1545.540 2085.110 1545.600 ;
        RECT 2084.345 1545.400 2085.110 1545.540 ;
        RECT 2084.345 1545.355 2084.635 1545.400 ;
        RECT 2084.790 1545.340 2085.110 1545.400 ;
        RECT 2084.330 1497.600 2084.650 1497.660 ;
        RECT 2084.135 1497.460 2084.650 1497.600 ;
        RECT 2084.330 1497.400 2084.650 1497.460 ;
        RECT 2084.330 1400.700 2084.650 1400.760 ;
        RECT 2084.135 1400.560 2084.650 1400.700 ;
        RECT 2084.330 1400.500 2084.650 1400.560 ;
        RECT 2084.345 1352.760 2084.635 1352.805 ;
        RECT 2084.790 1352.760 2085.110 1352.820 ;
        RECT 2084.345 1352.620 2085.110 1352.760 ;
        RECT 2084.345 1352.575 2084.635 1352.620 ;
        RECT 2084.790 1352.560 2085.110 1352.620 ;
        RECT 2084.330 1304.140 2084.650 1304.200 ;
        RECT 2084.135 1304.000 2084.650 1304.140 ;
        RECT 2084.330 1303.940 2084.650 1304.000 ;
        RECT 2084.345 1256.200 2084.635 1256.245 ;
        RECT 2084.790 1256.200 2085.110 1256.260 ;
        RECT 2084.345 1256.060 2085.110 1256.200 ;
        RECT 2084.345 1256.015 2084.635 1256.060 ;
        RECT 2084.790 1256.000 2085.110 1256.060 ;
        RECT 2084.790 1159.300 2085.110 1159.360 ;
        RECT 2085.710 1159.300 2086.030 1159.360 ;
        RECT 2084.790 1159.160 2086.030 1159.300 ;
        RECT 2084.790 1159.100 2085.110 1159.160 ;
        RECT 2085.710 1159.100 2086.030 1159.160 ;
        RECT 2084.790 1062.740 2085.110 1062.800 ;
        RECT 2085.710 1062.740 2086.030 1062.800 ;
        RECT 2084.790 1062.600 2086.030 1062.740 ;
        RECT 2084.790 1062.540 2085.110 1062.600 ;
        RECT 2085.710 1062.540 2086.030 1062.600 ;
        RECT 2084.790 966.180 2085.110 966.240 ;
        RECT 2085.710 966.180 2086.030 966.240 ;
        RECT 2084.790 966.040 2086.030 966.180 ;
        RECT 2084.790 965.980 2085.110 966.040 ;
        RECT 2085.710 965.980 2086.030 966.040 ;
        RECT 2084.790 869.620 2085.110 869.680 ;
        RECT 2085.710 869.620 2086.030 869.680 ;
        RECT 2084.790 869.480 2086.030 869.620 ;
        RECT 2084.790 869.420 2085.110 869.480 ;
        RECT 2085.710 869.420 2086.030 869.480 ;
        RECT 2084.330 821.000 2084.650 821.060 ;
        RECT 2085.710 821.000 2086.030 821.060 ;
        RECT 2084.330 820.860 2086.030 821.000 ;
        RECT 2084.330 820.800 2084.650 820.860 ;
        RECT 2085.710 820.800 2086.030 820.860 ;
        RECT 2084.330 689.900 2084.650 690.160 ;
        RECT 2083.870 689.760 2084.190 689.820 ;
        RECT 2084.420 689.760 2084.560 689.900 ;
        RECT 2083.870 689.620 2084.560 689.760 ;
        RECT 2083.870 689.560 2084.190 689.620 ;
        RECT 2084.330 593.340 2084.650 593.600 ;
        RECT 2083.870 593.200 2084.190 593.260 ;
        RECT 2084.420 593.200 2084.560 593.340 ;
        RECT 2083.870 593.060 2084.560 593.200 ;
        RECT 2083.870 593.000 2084.190 593.060 ;
        RECT 2084.330 496.780 2084.650 497.040 ;
        RECT 2083.870 496.640 2084.190 496.700 ;
        RECT 2084.420 496.640 2084.560 496.780 ;
        RECT 2083.870 496.500 2084.560 496.640 ;
        RECT 2083.870 496.440 2084.190 496.500 ;
        RECT 2083.870 386.820 2084.190 386.880 ;
        RECT 2084.790 386.820 2085.110 386.880 ;
        RECT 2083.870 386.680 2085.110 386.820 ;
        RECT 2083.870 386.620 2084.190 386.680 ;
        RECT 2084.790 386.620 2085.110 386.680 ;
        RECT 2084.345 386.140 2084.635 386.185 ;
        RECT 2084.790 386.140 2085.110 386.200 ;
        RECT 2084.345 386.000 2085.110 386.140 ;
        RECT 2084.345 385.955 2084.635 386.000 ;
        RECT 2084.790 385.940 2085.110 386.000 ;
        RECT 2084.330 338.200 2084.650 338.260 ;
        RECT 2084.135 338.060 2084.650 338.200 ;
        RECT 2084.330 338.000 2084.650 338.060 ;
        RECT 2083.870 303.520 2084.190 303.580 ;
        RECT 2084.790 303.520 2085.110 303.580 ;
        RECT 2083.870 303.380 2085.110 303.520 ;
        RECT 2083.870 303.320 2084.190 303.380 ;
        RECT 2084.790 303.320 2085.110 303.380 ;
        RECT 2084.345 289.580 2084.635 289.625 ;
        RECT 2084.790 289.580 2085.110 289.640 ;
        RECT 2084.345 289.440 2085.110 289.580 ;
        RECT 2084.345 289.395 2084.635 289.440 ;
        RECT 2084.790 289.380 2085.110 289.440 ;
        RECT 2084.330 241.980 2084.650 242.040 ;
        RECT 2084.135 241.840 2084.650 241.980 ;
        RECT 2084.330 241.780 2084.650 241.840 ;
        RECT 2084.330 241.300 2084.650 241.360 ;
        RECT 2085.250 241.300 2085.570 241.360 ;
        RECT 2084.330 241.160 2085.570 241.300 ;
        RECT 2084.330 241.100 2084.650 241.160 ;
        RECT 2085.250 241.100 2085.570 241.160 ;
        RECT 2084.345 193.020 2084.635 193.065 ;
        RECT 2084.790 193.020 2085.110 193.080 ;
        RECT 2084.345 192.880 2085.110 193.020 ;
        RECT 2084.345 192.835 2084.635 192.880 ;
        RECT 2084.790 192.820 2085.110 192.880 ;
        RECT 2084.330 145.080 2084.650 145.140 ;
        RECT 2084.135 144.940 2084.650 145.080 ;
        RECT 2084.330 144.880 2084.650 144.940 ;
        RECT 2083.870 110.400 2084.190 110.460 ;
        RECT 2084.790 110.400 2085.110 110.460 ;
        RECT 2083.870 110.260 2085.110 110.400 ;
        RECT 2083.870 110.200 2084.190 110.260 ;
        RECT 2084.790 110.200 2085.110 110.260 ;
        RECT 2084.790 96.460 2085.110 96.520 ;
        RECT 2084.595 96.320 2085.110 96.460 ;
        RECT 2084.790 96.260 2085.110 96.320 ;
        RECT 2084.790 61.440 2085.110 61.500 ;
        RECT 2084.595 61.300 2085.110 61.440 ;
        RECT 2084.790 61.240 2085.110 61.300 ;
        RECT 1828.570 25.060 1828.890 25.120 ;
        RECT 2084.790 25.060 2085.110 25.120 ;
        RECT 1828.570 24.920 2085.110 25.060 ;
        RECT 1828.570 24.860 1828.890 24.920 ;
        RECT 2084.790 24.860 2085.110 24.920 ;
      LAYER via ;
        RECT 2083.900 1655.840 2084.160 1656.100 ;
        RECT 2084.820 1655.840 2085.080 1656.100 ;
        RECT 2084.820 1641.900 2085.080 1642.160 ;
        RECT 2084.360 1593.960 2084.620 1594.220 ;
        RECT 2083.900 1558.940 2084.160 1559.200 ;
        RECT 2084.820 1558.940 2085.080 1559.200 ;
        RECT 2084.820 1545.340 2085.080 1545.600 ;
        RECT 2084.360 1497.400 2084.620 1497.660 ;
        RECT 2084.360 1400.500 2084.620 1400.760 ;
        RECT 2084.820 1352.560 2085.080 1352.820 ;
        RECT 2084.360 1303.940 2084.620 1304.200 ;
        RECT 2084.820 1256.000 2085.080 1256.260 ;
        RECT 2084.820 1159.100 2085.080 1159.360 ;
        RECT 2085.740 1159.100 2086.000 1159.360 ;
        RECT 2084.820 1062.540 2085.080 1062.800 ;
        RECT 2085.740 1062.540 2086.000 1062.800 ;
        RECT 2084.820 965.980 2085.080 966.240 ;
        RECT 2085.740 965.980 2086.000 966.240 ;
        RECT 2084.820 869.420 2085.080 869.680 ;
        RECT 2085.740 869.420 2086.000 869.680 ;
        RECT 2084.360 820.800 2084.620 821.060 ;
        RECT 2085.740 820.800 2086.000 821.060 ;
        RECT 2084.360 689.900 2084.620 690.160 ;
        RECT 2083.900 689.560 2084.160 689.820 ;
        RECT 2084.360 593.340 2084.620 593.600 ;
        RECT 2083.900 593.000 2084.160 593.260 ;
        RECT 2084.360 496.780 2084.620 497.040 ;
        RECT 2083.900 496.440 2084.160 496.700 ;
        RECT 2083.900 386.620 2084.160 386.880 ;
        RECT 2084.820 386.620 2085.080 386.880 ;
        RECT 2084.820 385.940 2085.080 386.200 ;
        RECT 2084.360 338.000 2084.620 338.260 ;
        RECT 2083.900 303.320 2084.160 303.580 ;
        RECT 2084.820 303.320 2085.080 303.580 ;
        RECT 2084.820 289.380 2085.080 289.640 ;
        RECT 2084.360 241.780 2084.620 242.040 ;
        RECT 2084.360 241.100 2084.620 241.360 ;
        RECT 2085.280 241.100 2085.540 241.360 ;
        RECT 2084.820 192.820 2085.080 193.080 ;
        RECT 2084.360 144.880 2084.620 145.140 ;
        RECT 2083.900 110.200 2084.160 110.460 ;
        RECT 2084.820 110.200 2085.080 110.460 ;
        RECT 2084.820 96.260 2085.080 96.520 ;
        RECT 2084.820 61.240 2085.080 61.500 ;
        RECT 1828.600 24.860 1828.860 25.120 ;
        RECT 2084.820 24.860 2085.080 25.120 ;
      LAYER met2 ;
        RECT 2089.800 1700.410 2090.080 1702.400 ;
        RECT 2087.180 1700.270 2090.080 1700.410 ;
        RECT 2087.180 1677.970 2087.320 1700.270 ;
        RECT 2089.800 1700.000 2090.080 1700.270 ;
        RECT 2083.960 1677.830 2087.320 1677.970 ;
        RECT 2083.960 1656.130 2084.100 1677.830 ;
        RECT 2083.900 1655.810 2084.160 1656.130 ;
        RECT 2084.820 1655.810 2085.080 1656.130 ;
        RECT 2084.880 1642.190 2085.020 1655.810 ;
        RECT 2084.820 1641.870 2085.080 1642.190 ;
        RECT 2084.360 1593.930 2084.620 1594.250 ;
        RECT 2084.420 1559.650 2084.560 1593.930 ;
        RECT 2083.960 1559.510 2084.560 1559.650 ;
        RECT 2083.960 1559.230 2084.100 1559.510 ;
        RECT 2083.900 1558.910 2084.160 1559.230 ;
        RECT 2084.820 1558.910 2085.080 1559.230 ;
        RECT 2084.880 1545.630 2085.020 1558.910 ;
        RECT 2084.820 1545.310 2085.080 1545.630 ;
        RECT 2084.360 1497.370 2084.620 1497.690 ;
        RECT 2084.420 1473.290 2084.560 1497.370 ;
        RECT 2084.420 1473.150 2085.020 1473.290 ;
        RECT 2084.880 1414.130 2085.020 1473.150 ;
        RECT 2084.420 1413.990 2085.020 1414.130 ;
        RECT 2084.420 1400.790 2084.560 1413.990 ;
        RECT 2084.360 1400.470 2084.620 1400.790 ;
        RECT 2084.820 1352.530 2085.080 1352.850 ;
        RECT 2084.880 1317.570 2085.020 1352.530 ;
        RECT 2084.420 1317.430 2085.020 1317.570 ;
        RECT 2084.420 1304.230 2084.560 1317.430 ;
        RECT 2084.360 1303.910 2084.620 1304.230 ;
        RECT 2084.820 1255.970 2085.080 1256.290 ;
        RECT 2084.880 1221.010 2085.020 1255.970 ;
        RECT 2084.420 1220.870 2085.020 1221.010 ;
        RECT 2084.420 1207.525 2084.560 1220.870 ;
        RECT 2084.350 1207.155 2084.630 1207.525 ;
        RECT 2085.730 1207.155 2086.010 1207.525 ;
        RECT 2085.800 1159.390 2085.940 1207.155 ;
        RECT 2084.820 1159.070 2085.080 1159.390 ;
        RECT 2085.740 1159.070 2086.000 1159.390 ;
        RECT 2084.880 1124.450 2085.020 1159.070 ;
        RECT 2084.420 1124.310 2085.020 1124.450 ;
        RECT 2084.420 1110.965 2084.560 1124.310 ;
        RECT 2084.350 1110.595 2084.630 1110.965 ;
        RECT 2085.730 1110.595 2086.010 1110.965 ;
        RECT 2085.800 1062.830 2085.940 1110.595 ;
        RECT 2084.820 1062.510 2085.080 1062.830 ;
        RECT 2085.740 1062.510 2086.000 1062.830 ;
        RECT 2084.880 1027.890 2085.020 1062.510 ;
        RECT 2084.420 1027.750 2085.020 1027.890 ;
        RECT 2084.420 1014.405 2084.560 1027.750 ;
        RECT 2084.350 1014.035 2084.630 1014.405 ;
        RECT 2085.730 1014.035 2086.010 1014.405 ;
        RECT 2085.800 966.270 2085.940 1014.035 ;
        RECT 2084.820 965.950 2085.080 966.270 ;
        RECT 2085.740 965.950 2086.000 966.270 ;
        RECT 2084.880 931.330 2085.020 965.950 ;
        RECT 2084.420 931.190 2085.020 931.330 ;
        RECT 2084.420 917.845 2084.560 931.190 ;
        RECT 2084.350 917.475 2084.630 917.845 ;
        RECT 2085.730 917.475 2086.010 917.845 ;
        RECT 2085.800 869.710 2085.940 917.475 ;
        RECT 2084.820 869.390 2085.080 869.710 ;
        RECT 2085.740 869.390 2086.000 869.710 ;
        RECT 2084.880 834.770 2085.020 869.390 ;
        RECT 2084.420 834.630 2085.020 834.770 ;
        RECT 2084.420 821.090 2084.560 834.630 ;
        RECT 2084.360 820.770 2084.620 821.090 ;
        RECT 2085.740 820.770 2086.000 821.090 ;
        RECT 2085.800 773.005 2085.940 820.770 ;
        RECT 2084.810 772.635 2085.090 773.005 ;
        RECT 2085.730 772.635 2086.010 773.005 ;
        RECT 2084.880 738.210 2085.020 772.635 ;
        RECT 2084.420 738.070 2085.020 738.210 ;
        RECT 2084.420 690.190 2084.560 738.070 ;
        RECT 2084.360 689.870 2084.620 690.190 ;
        RECT 2083.900 689.530 2084.160 689.850 ;
        RECT 2083.960 676.445 2084.100 689.530 ;
        RECT 2083.890 676.075 2084.170 676.445 ;
        RECT 2084.810 676.075 2085.090 676.445 ;
        RECT 2084.880 641.650 2085.020 676.075 ;
        RECT 2084.420 641.510 2085.020 641.650 ;
        RECT 2084.420 593.630 2084.560 641.510 ;
        RECT 2084.360 593.310 2084.620 593.630 ;
        RECT 2083.900 592.970 2084.160 593.290 ;
        RECT 2083.960 579.885 2084.100 592.970 ;
        RECT 2083.890 579.515 2084.170 579.885 ;
        RECT 2084.810 579.515 2085.090 579.885 ;
        RECT 2084.880 545.090 2085.020 579.515 ;
        RECT 2084.420 544.950 2085.020 545.090 ;
        RECT 2084.420 497.070 2084.560 544.950 ;
        RECT 2084.360 496.750 2084.620 497.070 ;
        RECT 2083.900 496.410 2084.160 496.730 ;
        RECT 2083.960 483.325 2084.100 496.410 ;
        RECT 2083.890 482.955 2084.170 483.325 ;
        RECT 2084.810 482.955 2085.090 483.325 ;
        RECT 2084.880 448.530 2085.020 482.955 ;
        RECT 2084.420 448.390 2085.020 448.530 ;
        RECT 2084.420 410.450 2084.560 448.390 ;
        RECT 2083.960 410.310 2084.560 410.450 ;
        RECT 2083.960 386.910 2084.100 410.310 ;
        RECT 2083.900 386.590 2084.160 386.910 ;
        RECT 2084.820 386.590 2085.080 386.910 ;
        RECT 2084.880 386.230 2085.020 386.590 ;
        RECT 2084.820 385.910 2085.080 386.230 ;
        RECT 2084.360 337.970 2084.620 338.290 ;
        RECT 2084.420 303.690 2084.560 337.970 ;
        RECT 2083.960 303.610 2084.560 303.690 ;
        RECT 2083.900 303.550 2084.560 303.610 ;
        RECT 2083.900 303.290 2084.160 303.550 ;
        RECT 2084.820 303.290 2085.080 303.610 ;
        RECT 2084.880 289.670 2085.020 303.290 ;
        RECT 2084.820 289.350 2085.080 289.670 ;
        RECT 2084.360 241.750 2084.620 242.070 ;
        RECT 2084.420 241.390 2084.560 241.750 ;
        RECT 2084.360 241.070 2084.620 241.390 ;
        RECT 2085.280 241.070 2085.540 241.390 ;
        RECT 2085.340 193.530 2085.480 241.070 ;
        RECT 2084.880 193.390 2085.480 193.530 ;
        RECT 2084.880 193.110 2085.020 193.390 ;
        RECT 2084.820 192.790 2085.080 193.110 ;
        RECT 2084.360 144.850 2084.620 145.170 ;
        RECT 2084.420 110.570 2084.560 144.850 ;
        RECT 2083.960 110.490 2084.560 110.570 ;
        RECT 2083.900 110.430 2084.560 110.490 ;
        RECT 2083.900 110.170 2084.160 110.430 ;
        RECT 2084.820 110.170 2085.080 110.490 ;
        RECT 2084.880 96.550 2085.020 110.170 ;
        RECT 2084.820 96.230 2085.080 96.550 ;
        RECT 2084.820 61.210 2085.080 61.530 ;
        RECT 2084.880 25.150 2085.020 61.210 ;
        RECT 1828.600 24.830 1828.860 25.150 ;
        RECT 2084.820 24.830 2085.080 25.150 ;
        RECT 1828.660 2.400 1828.800 24.830 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
      LAYER via2 ;
        RECT 2084.350 1207.200 2084.630 1207.480 ;
        RECT 2085.730 1207.200 2086.010 1207.480 ;
        RECT 2084.350 1110.640 2084.630 1110.920 ;
        RECT 2085.730 1110.640 2086.010 1110.920 ;
        RECT 2084.350 1014.080 2084.630 1014.360 ;
        RECT 2085.730 1014.080 2086.010 1014.360 ;
        RECT 2084.350 917.520 2084.630 917.800 ;
        RECT 2085.730 917.520 2086.010 917.800 ;
        RECT 2084.810 772.680 2085.090 772.960 ;
        RECT 2085.730 772.680 2086.010 772.960 ;
        RECT 2083.890 676.120 2084.170 676.400 ;
        RECT 2084.810 676.120 2085.090 676.400 ;
        RECT 2083.890 579.560 2084.170 579.840 ;
        RECT 2084.810 579.560 2085.090 579.840 ;
        RECT 2083.890 483.000 2084.170 483.280 ;
        RECT 2084.810 483.000 2085.090 483.280 ;
      LAYER met3 ;
        RECT 2084.325 1207.490 2084.655 1207.505 ;
        RECT 2085.705 1207.490 2086.035 1207.505 ;
        RECT 2084.325 1207.190 2086.035 1207.490 ;
        RECT 2084.325 1207.175 2084.655 1207.190 ;
        RECT 2085.705 1207.175 2086.035 1207.190 ;
        RECT 2084.325 1110.930 2084.655 1110.945 ;
        RECT 2085.705 1110.930 2086.035 1110.945 ;
        RECT 2084.325 1110.630 2086.035 1110.930 ;
        RECT 2084.325 1110.615 2084.655 1110.630 ;
        RECT 2085.705 1110.615 2086.035 1110.630 ;
        RECT 2084.325 1014.370 2084.655 1014.385 ;
        RECT 2085.705 1014.370 2086.035 1014.385 ;
        RECT 2084.325 1014.070 2086.035 1014.370 ;
        RECT 2084.325 1014.055 2084.655 1014.070 ;
        RECT 2085.705 1014.055 2086.035 1014.070 ;
        RECT 2084.325 917.810 2084.655 917.825 ;
        RECT 2085.705 917.810 2086.035 917.825 ;
        RECT 2084.325 917.510 2086.035 917.810 ;
        RECT 2084.325 917.495 2084.655 917.510 ;
        RECT 2085.705 917.495 2086.035 917.510 ;
        RECT 2084.785 772.970 2085.115 772.985 ;
        RECT 2085.705 772.970 2086.035 772.985 ;
        RECT 2084.785 772.670 2086.035 772.970 ;
        RECT 2084.785 772.655 2085.115 772.670 ;
        RECT 2085.705 772.655 2086.035 772.670 ;
        RECT 2083.865 676.410 2084.195 676.425 ;
        RECT 2084.785 676.410 2085.115 676.425 ;
        RECT 2083.865 676.110 2085.115 676.410 ;
        RECT 2083.865 676.095 2084.195 676.110 ;
        RECT 2084.785 676.095 2085.115 676.110 ;
        RECT 2083.865 579.850 2084.195 579.865 ;
        RECT 2084.785 579.850 2085.115 579.865 ;
        RECT 2083.865 579.550 2085.115 579.850 ;
        RECT 2083.865 579.535 2084.195 579.550 ;
        RECT 2084.785 579.535 2085.115 579.550 ;
        RECT 2083.865 483.290 2084.195 483.305 ;
        RECT 2084.785 483.290 2085.115 483.305 ;
        RECT 2083.865 482.990 2085.115 483.290 ;
        RECT 2083.865 482.975 2084.195 482.990 ;
        RECT 2084.785 482.975 2085.115 482.990 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1846.050 29.140 1846.370 29.200 ;
        RECT 2098.130 29.140 2098.450 29.200 ;
        RECT 1846.050 29.000 2098.450 29.140 ;
        RECT 1846.050 28.940 1846.370 29.000 ;
        RECT 2098.130 28.940 2098.450 29.000 ;
      LAYER via ;
        RECT 1846.080 28.940 1846.340 29.200 ;
        RECT 2098.160 28.940 2098.420 29.200 ;
      LAYER met2 ;
        RECT 2099.000 1700.410 2099.280 1702.400 ;
        RECT 2098.220 1700.270 2099.280 1700.410 ;
        RECT 2098.220 29.230 2098.360 1700.270 ;
        RECT 2099.000 1700.000 2099.280 1700.270 ;
        RECT 1846.080 28.910 1846.340 29.230 ;
        RECT 2098.160 28.910 2098.420 29.230 ;
        RECT 1846.140 2.400 1846.280 28.910 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1864.450 30.840 1864.770 30.900 ;
        RECT 2105.490 30.840 2105.810 30.900 ;
        RECT 1864.450 30.700 2105.810 30.840 ;
        RECT 1864.450 30.640 1864.770 30.700 ;
        RECT 2105.490 30.640 2105.810 30.700 ;
      LAYER via ;
        RECT 1864.480 30.640 1864.740 30.900 ;
        RECT 2105.520 30.640 2105.780 30.900 ;
      LAYER met2 ;
        RECT 2108.200 1700.410 2108.480 1702.400 ;
        RECT 2105.580 1700.270 2108.480 1700.410 ;
        RECT 2105.580 30.930 2105.720 1700.270 ;
        RECT 2108.200 1700.000 2108.480 1700.270 ;
        RECT 1864.480 30.610 1864.740 30.930 ;
        RECT 2105.520 30.610 2105.780 30.930 ;
        RECT 1864.540 22.170 1864.680 30.610 ;
        RECT 1864.080 22.030 1864.680 22.170 ;
        RECT 1864.080 2.400 1864.220 22.030 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1525.965 1449.165 1526.135 1497.275 ;
        RECT 1525.965 1352.605 1526.135 1400.715 ;
        RECT 1525.965 1256.045 1526.135 1304.155 ;
        RECT 1525.965 579.785 1526.135 603.755 ;
        RECT 1525.965 483.225 1526.135 531.335 ;
        RECT 1525.965 386.325 1526.135 434.775 ;
        RECT 1525.505 96.645 1525.675 111.095 ;
      LAYER mcon ;
        RECT 1525.965 1497.105 1526.135 1497.275 ;
        RECT 1525.965 1400.545 1526.135 1400.715 ;
        RECT 1525.965 1303.985 1526.135 1304.155 ;
        RECT 1525.965 603.585 1526.135 603.755 ;
        RECT 1525.965 531.165 1526.135 531.335 ;
        RECT 1525.965 434.605 1526.135 434.775 ;
        RECT 1525.505 110.925 1525.675 111.095 ;
      LAYER met1 ;
        RECT 1525.890 1655.840 1526.210 1656.100 ;
        RECT 1525.980 1655.700 1526.120 1655.840 ;
        RECT 1526.350 1655.700 1526.670 1655.760 ;
        RECT 1525.980 1655.560 1526.670 1655.700 ;
        RECT 1526.350 1655.500 1526.670 1655.560 ;
        RECT 1525.890 1545.880 1526.210 1545.940 ;
        RECT 1526.350 1545.880 1526.670 1545.940 ;
        RECT 1525.890 1545.740 1526.670 1545.880 ;
        RECT 1525.890 1545.680 1526.210 1545.740 ;
        RECT 1526.350 1545.680 1526.670 1545.740 ;
        RECT 1525.890 1497.260 1526.210 1497.320 ;
        RECT 1525.695 1497.120 1526.210 1497.260 ;
        RECT 1525.890 1497.060 1526.210 1497.120 ;
        RECT 1525.890 1449.320 1526.210 1449.380 ;
        RECT 1525.695 1449.180 1526.210 1449.320 ;
        RECT 1525.890 1449.120 1526.210 1449.180 ;
        RECT 1525.890 1400.700 1526.210 1400.760 ;
        RECT 1525.695 1400.560 1526.210 1400.700 ;
        RECT 1525.890 1400.500 1526.210 1400.560 ;
        RECT 1525.890 1352.760 1526.210 1352.820 ;
        RECT 1525.695 1352.620 1526.210 1352.760 ;
        RECT 1525.890 1352.560 1526.210 1352.620 ;
        RECT 1525.890 1304.140 1526.210 1304.200 ;
        RECT 1525.695 1304.000 1526.210 1304.140 ;
        RECT 1525.890 1303.940 1526.210 1304.000 ;
        RECT 1525.890 1256.200 1526.210 1256.260 ;
        RECT 1525.695 1256.060 1526.210 1256.200 ;
        RECT 1525.890 1256.000 1526.210 1256.060 ;
        RECT 1525.890 1159.300 1526.210 1159.360 ;
        RECT 1526.810 1159.300 1527.130 1159.360 ;
        RECT 1525.890 1159.160 1527.130 1159.300 ;
        RECT 1525.890 1159.100 1526.210 1159.160 ;
        RECT 1526.810 1159.100 1527.130 1159.160 ;
        RECT 1525.890 1062.740 1526.210 1062.800 ;
        RECT 1526.810 1062.740 1527.130 1062.800 ;
        RECT 1525.890 1062.600 1527.130 1062.740 ;
        RECT 1525.890 1062.540 1526.210 1062.600 ;
        RECT 1526.810 1062.540 1527.130 1062.600 ;
        RECT 1525.890 966.180 1526.210 966.240 ;
        RECT 1526.810 966.180 1527.130 966.240 ;
        RECT 1525.890 966.040 1527.130 966.180 ;
        RECT 1525.890 965.980 1526.210 966.040 ;
        RECT 1526.810 965.980 1527.130 966.040 ;
        RECT 1525.890 869.620 1526.210 869.680 ;
        RECT 1526.810 869.620 1527.130 869.680 ;
        RECT 1525.890 869.480 1527.130 869.620 ;
        RECT 1525.890 869.420 1526.210 869.480 ;
        RECT 1526.810 869.420 1527.130 869.480 ;
        RECT 1525.890 821.000 1526.210 821.060 ;
        RECT 1526.350 821.000 1526.670 821.060 ;
        RECT 1525.890 820.860 1526.670 821.000 ;
        RECT 1525.890 820.800 1526.210 820.860 ;
        RECT 1526.350 820.800 1526.670 820.860 ;
        RECT 1525.905 603.740 1526.195 603.785 ;
        RECT 1526.350 603.740 1526.670 603.800 ;
        RECT 1525.905 603.600 1526.670 603.740 ;
        RECT 1525.905 603.555 1526.195 603.600 ;
        RECT 1526.350 603.540 1526.670 603.600 ;
        RECT 1525.890 579.940 1526.210 580.000 ;
        RECT 1525.695 579.800 1526.210 579.940 ;
        RECT 1525.890 579.740 1526.210 579.800 ;
        RECT 1525.890 531.320 1526.210 531.380 ;
        RECT 1525.695 531.180 1526.210 531.320 ;
        RECT 1525.890 531.120 1526.210 531.180 ;
        RECT 1525.890 483.380 1526.210 483.440 ;
        RECT 1525.695 483.240 1526.210 483.380 ;
        RECT 1525.890 483.180 1526.210 483.240 ;
        RECT 1525.890 434.760 1526.210 434.820 ;
        RECT 1525.695 434.620 1526.210 434.760 ;
        RECT 1525.890 434.560 1526.210 434.620 ;
        RECT 1525.890 386.480 1526.210 386.540 ;
        RECT 1525.695 386.340 1526.210 386.480 ;
        RECT 1525.890 386.280 1526.210 386.340 ;
        RECT 1525.890 337.860 1526.210 337.920 ;
        RECT 1526.350 337.860 1526.670 337.920 ;
        RECT 1525.890 337.720 1526.670 337.860 ;
        RECT 1525.890 337.660 1526.210 337.720 ;
        RECT 1526.350 337.660 1526.670 337.720 ;
        RECT 1525.445 111.080 1525.735 111.125 ;
        RECT 1526.350 111.080 1526.670 111.140 ;
        RECT 1525.445 110.940 1526.670 111.080 ;
        RECT 1525.445 110.895 1525.735 110.940 ;
        RECT 1526.350 110.880 1526.670 110.940 ;
        RECT 1525.430 96.800 1525.750 96.860 ;
        RECT 1525.235 96.660 1525.750 96.800 ;
        RECT 1525.430 96.600 1525.750 96.660 ;
        RECT 744.810 67.560 745.130 67.620 ;
        RECT 1525.430 67.560 1525.750 67.620 ;
        RECT 744.810 67.420 1525.750 67.560 ;
        RECT 744.810 67.360 745.130 67.420 ;
        RECT 1525.430 67.360 1525.750 67.420 ;
      LAYER via ;
        RECT 1525.920 1655.840 1526.180 1656.100 ;
        RECT 1526.380 1655.500 1526.640 1655.760 ;
        RECT 1525.920 1545.680 1526.180 1545.940 ;
        RECT 1526.380 1545.680 1526.640 1545.940 ;
        RECT 1525.920 1497.060 1526.180 1497.320 ;
        RECT 1525.920 1449.120 1526.180 1449.380 ;
        RECT 1525.920 1400.500 1526.180 1400.760 ;
        RECT 1525.920 1352.560 1526.180 1352.820 ;
        RECT 1525.920 1303.940 1526.180 1304.200 ;
        RECT 1525.920 1256.000 1526.180 1256.260 ;
        RECT 1525.920 1159.100 1526.180 1159.360 ;
        RECT 1526.840 1159.100 1527.100 1159.360 ;
        RECT 1525.920 1062.540 1526.180 1062.800 ;
        RECT 1526.840 1062.540 1527.100 1062.800 ;
        RECT 1525.920 965.980 1526.180 966.240 ;
        RECT 1526.840 965.980 1527.100 966.240 ;
        RECT 1525.920 869.420 1526.180 869.680 ;
        RECT 1526.840 869.420 1527.100 869.680 ;
        RECT 1525.920 820.800 1526.180 821.060 ;
        RECT 1526.380 820.800 1526.640 821.060 ;
        RECT 1526.380 603.540 1526.640 603.800 ;
        RECT 1525.920 579.740 1526.180 580.000 ;
        RECT 1525.920 531.120 1526.180 531.380 ;
        RECT 1525.920 483.180 1526.180 483.440 ;
        RECT 1525.920 434.560 1526.180 434.820 ;
        RECT 1525.920 386.280 1526.180 386.540 ;
        RECT 1525.920 337.660 1526.180 337.920 ;
        RECT 1526.380 337.660 1526.640 337.920 ;
        RECT 1526.380 110.880 1526.640 111.140 ;
        RECT 1525.460 96.600 1525.720 96.860 ;
        RECT 744.840 67.360 745.100 67.620 ;
        RECT 1525.460 67.360 1525.720 67.620 ;
      LAYER met2 ;
        RECT 1529.520 1700.410 1529.800 1702.400 ;
        RECT 1526.900 1700.270 1529.800 1700.410 ;
        RECT 1526.900 1677.970 1527.040 1700.270 ;
        RECT 1529.520 1700.000 1529.800 1700.270 ;
        RECT 1525.980 1677.830 1527.040 1677.970 ;
        RECT 1525.980 1656.130 1526.120 1677.830 ;
        RECT 1525.920 1655.810 1526.180 1656.130 ;
        RECT 1526.380 1655.470 1526.640 1655.790 ;
        RECT 1526.440 1545.970 1526.580 1655.470 ;
        RECT 1525.920 1545.650 1526.180 1545.970 ;
        RECT 1526.380 1545.650 1526.640 1545.970 ;
        RECT 1525.980 1497.350 1526.120 1545.650 ;
        RECT 1525.920 1497.030 1526.180 1497.350 ;
        RECT 1525.920 1449.090 1526.180 1449.410 ;
        RECT 1525.980 1400.790 1526.120 1449.090 ;
        RECT 1525.920 1400.470 1526.180 1400.790 ;
        RECT 1525.920 1352.530 1526.180 1352.850 ;
        RECT 1525.980 1304.230 1526.120 1352.530 ;
        RECT 1525.920 1303.910 1526.180 1304.230 ;
        RECT 1525.920 1255.970 1526.180 1256.290 ;
        RECT 1525.980 1207.525 1526.120 1255.970 ;
        RECT 1525.910 1207.155 1526.190 1207.525 ;
        RECT 1526.830 1207.155 1527.110 1207.525 ;
        RECT 1526.900 1159.390 1527.040 1207.155 ;
        RECT 1525.920 1159.070 1526.180 1159.390 ;
        RECT 1526.840 1159.070 1527.100 1159.390 ;
        RECT 1525.980 1110.965 1526.120 1159.070 ;
        RECT 1525.910 1110.595 1526.190 1110.965 ;
        RECT 1526.830 1110.595 1527.110 1110.965 ;
        RECT 1526.900 1062.830 1527.040 1110.595 ;
        RECT 1525.920 1062.510 1526.180 1062.830 ;
        RECT 1526.840 1062.510 1527.100 1062.830 ;
        RECT 1525.980 1014.405 1526.120 1062.510 ;
        RECT 1525.910 1014.035 1526.190 1014.405 ;
        RECT 1526.830 1014.035 1527.110 1014.405 ;
        RECT 1526.900 966.270 1527.040 1014.035 ;
        RECT 1525.920 965.950 1526.180 966.270 ;
        RECT 1526.840 965.950 1527.100 966.270 ;
        RECT 1525.980 917.845 1526.120 965.950 ;
        RECT 1525.910 917.475 1526.190 917.845 ;
        RECT 1526.830 917.475 1527.110 917.845 ;
        RECT 1526.900 869.710 1527.040 917.475 ;
        RECT 1525.920 869.390 1526.180 869.710 ;
        RECT 1526.840 869.390 1527.100 869.710 ;
        RECT 1525.980 821.090 1526.120 869.390 ;
        RECT 1525.920 820.770 1526.180 821.090 ;
        RECT 1526.380 820.770 1526.640 821.090 ;
        RECT 1526.440 603.830 1526.580 820.770 ;
        RECT 1526.380 603.510 1526.640 603.830 ;
        RECT 1525.920 579.710 1526.180 580.030 ;
        RECT 1525.980 531.410 1526.120 579.710 ;
        RECT 1525.920 531.090 1526.180 531.410 ;
        RECT 1525.920 483.150 1526.180 483.470 ;
        RECT 1525.980 434.850 1526.120 483.150 ;
        RECT 1525.920 434.530 1526.180 434.850 ;
        RECT 1525.920 386.250 1526.180 386.570 ;
        RECT 1525.980 337.950 1526.120 386.250 ;
        RECT 1525.920 337.630 1526.180 337.950 ;
        RECT 1526.380 337.630 1526.640 337.950 ;
        RECT 1526.440 111.170 1526.580 337.630 ;
        RECT 1526.380 110.850 1526.640 111.170 ;
        RECT 1525.460 96.570 1525.720 96.890 ;
        RECT 1525.520 67.650 1525.660 96.570 ;
        RECT 744.840 67.330 745.100 67.650 ;
        RECT 1525.460 67.330 1525.720 67.650 ;
        RECT 744.900 16.730 745.040 67.330 ;
        RECT 740.300 16.590 745.040 16.730 ;
        RECT 740.300 2.400 740.440 16.590 ;
        RECT 740.090 -4.800 740.650 2.400 ;
      LAYER via2 ;
        RECT 1525.910 1207.200 1526.190 1207.480 ;
        RECT 1526.830 1207.200 1527.110 1207.480 ;
        RECT 1525.910 1110.640 1526.190 1110.920 ;
        RECT 1526.830 1110.640 1527.110 1110.920 ;
        RECT 1525.910 1014.080 1526.190 1014.360 ;
        RECT 1526.830 1014.080 1527.110 1014.360 ;
        RECT 1525.910 917.520 1526.190 917.800 ;
        RECT 1526.830 917.520 1527.110 917.800 ;
      LAYER met3 ;
        RECT 1525.885 1207.490 1526.215 1207.505 ;
        RECT 1526.805 1207.490 1527.135 1207.505 ;
        RECT 1525.885 1207.190 1527.135 1207.490 ;
        RECT 1525.885 1207.175 1526.215 1207.190 ;
        RECT 1526.805 1207.175 1527.135 1207.190 ;
        RECT 1525.885 1110.930 1526.215 1110.945 ;
        RECT 1526.805 1110.930 1527.135 1110.945 ;
        RECT 1525.885 1110.630 1527.135 1110.930 ;
        RECT 1525.885 1110.615 1526.215 1110.630 ;
        RECT 1526.805 1110.615 1527.135 1110.630 ;
        RECT 1525.885 1014.370 1526.215 1014.385 ;
        RECT 1526.805 1014.370 1527.135 1014.385 ;
        RECT 1525.885 1014.070 1527.135 1014.370 ;
        RECT 1525.885 1014.055 1526.215 1014.070 ;
        RECT 1526.805 1014.055 1527.135 1014.070 ;
        RECT 1525.885 917.810 1526.215 917.825 ;
        RECT 1526.805 917.810 1527.135 917.825 ;
        RECT 1525.885 917.510 1527.135 917.810 ;
        RECT 1525.885 917.495 1526.215 917.510 ;
        RECT 1526.805 917.495 1527.135 917.510 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2112.005 1594.005 2112.175 1642.115 ;
        RECT 2112.465 1499.485 2112.635 1545.555 ;
        RECT 2112.005 786.505 2112.175 821.015 ;
        RECT 2112.005 689.605 2112.175 724.455 ;
        RECT 2112.005 593.045 2112.175 627.895 ;
        RECT 2112.005 496.485 2112.175 531.335 ;
        RECT 2112.005 386.325 2112.175 434.775 ;
        RECT 2112.465 138.125 2112.635 193.035 ;
      LAYER mcon ;
        RECT 2112.005 1641.945 2112.175 1642.115 ;
        RECT 2112.465 1545.385 2112.635 1545.555 ;
        RECT 2112.005 820.845 2112.175 821.015 ;
        RECT 2112.005 724.285 2112.175 724.455 ;
        RECT 2112.005 627.725 2112.175 627.895 ;
        RECT 2112.005 531.165 2112.175 531.335 ;
        RECT 2112.005 434.605 2112.175 434.775 ;
        RECT 2112.465 192.865 2112.635 193.035 ;
      LAYER met1 ;
        RECT 2111.470 1678.140 2111.790 1678.200 ;
        RECT 2116.070 1678.140 2116.390 1678.200 ;
        RECT 2111.470 1678.000 2116.390 1678.140 ;
        RECT 2111.470 1677.940 2111.790 1678.000 ;
        RECT 2116.070 1677.940 2116.390 1678.000 ;
        RECT 2111.470 1656.040 2111.790 1656.100 ;
        RECT 2112.390 1656.040 2112.710 1656.100 ;
        RECT 2111.470 1655.900 2112.710 1656.040 ;
        RECT 2111.470 1655.840 2111.790 1655.900 ;
        RECT 2112.390 1655.840 2112.710 1655.900 ;
        RECT 2111.945 1642.100 2112.235 1642.145 ;
        RECT 2112.390 1642.100 2112.710 1642.160 ;
        RECT 2111.945 1641.960 2112.710 1642.100 ;
        RECT 2111.945 1641.915 2112.235 1641.960 ;
        RECT 2112.390 1641.900 2112.710 1641.960 ;
        RECT 2111.930 1594.160 2112.250 1594.220 ;
        RECT 2111.735 1594.020 2112.250 1594.160 ;
        RECT 2111.930 1593.960 2112.250 1594.020 ;
        RECT 2111.470 1559.140 2111.790 1559.200 ;
        RECT 2112.390 1559.140 2112.710 1559.200 ;
        RECT 2111.470 1559.000 2112.710 1559.140 ;
        RECT 2111.470 1558.940 2111.790 1559.000 ;
        RECT 2112.390 1558.940 2112.710 1559.000 ;
        RECT 2112.390 1545.540 2112.710 1545.600 ;
        RECT 2112.195 1545.400 2112.710 1545.540 ;
        RECT 2112.390 1545.340 2112.710 1545.400 ;
        RECT 2112.390 1499.640 2112.710 1499.700 ;
        RECT 2112.195 1499.500 2112.710 1499.640 ;
        RECT 2112.390 1499.440 2112.710 1499.500 ;
        RECT 2111.470 1414.640 2111.790 1414.700 ;
        RECT 2112.390 1414.640 2112.710 1414.700 ;
        RECT 2111.470 1414.500 2112.710 1414.640 ;
        RECT 2111.470 1414.440 2111.790 1414.500 ;
        RECT 2112.390 1414.440 2112.710 1414.500 ;
        RECT 2111.470 1318.080 2111.790 1318.140 ;
        RECT 2112.390 1318.080 2112.710 1318.140 ;
        RECT 2111.470 1317.940 2112.710 1318.080 ;
        RECT 2111.470 1317.880 2111.790 1317.940 ;
        RECT 2112.390 1317.880 2112.710 1317.940 ;
        RECT 2111.470 1221.520 2111.790 1221.580 ;
        RECT 2112.390 1221.520 2112.710 1221.580 ;
        RECT 2111.470 1221.380 2112.710 1221.520 ;
        RECT 2111.470 1221.320 2111.790 1221.380 ;
        RECT 2112.390 1221.320 2112.710 1221.380 ;
        RECT 2111.470 1124.960 2111.790 1125.020 ;
        RECT 2112.390 1124.960 2112.710 1125.020 ;
        RECT 2111.470 1124.820 2112.710 1124.960 ;
        RECT 2111.470 1124.760 2111.790 1124.820 ;
        RECT 2112.390 1124.760 2112.710 1124.820 ;
        RECT 2111.470 1028.400 2111.790 1028.460 ;
        RECT 2112.390 1028.400 2112.710 1028.460 ;
        RECT 2111.470 1028.260 2112.710 1028.400 ;
        RECT 2111.470 1028.200 2111.790 1028.260 ;
        RECT 2112.390 1028.200 2112.710 1028.260 ;
        RECT 2111.470 931.840 2111.790 931.900 ;
        RECT 2112.390 931.840 2112.710 931.900 ;
        RECT 2111.470 931.700 2112.710 931.840 ;
        RECT 2111.470 931.640 2111.790 931.700 ;
        RECT 2112.390 931.640 2112.710 931.700 ;
        RECT 2112.390 869.620 2112.710 869.680 ;
        RECT 2113.310 869.620 2113.630 869.680 ;
        RECT 2112.390 869.480 2113.630 869.620 ;
        RECT 2112.390 869.420 2112.710 869.480 ;
        RECT 2113.310 869.420 2113.630 869.480 ;
        RECT 2111.470 835.280 2111.790 835.340 ;
        RECT 2112.390 835.280 2112.710 835.340 ;
        RECT 2111.470 835.140 2112.710 835.280 ;
        RECT 2111.470 835.080 2111.790 835.140 ;
        RECT 2112.390 835.080 2112.710 835.140 ;
        RECT 2111.930 821.000 2112.250 821.060 ;
        RECT 2111.735 820.860 2112.250 821.000 ;
        RECT 2111.930 820.800 2112.250 820.860 ;
        RECT 2111.930 786.660 2112.250 786.720 ;
        RECT 2111.735 786.520 2112.250 786.660 ;
        RECT 2111.930 786.460 2112.250 786.520 ;
        RECT 2111.470 738.380 2111.790 738.440 ;
        RECT 2112.390 738.380 2112.710 738.440 ;
        RECT 2111.470 738.240 2112.710 738.380 ;
        RECT 2111.470 738.180 2111.790 738.240 ;
        RECT 2112.390 738.180 2112.710 738.240 ;
        RECT 2111.930 724.440 2112.250 724.500 ;
        RECT 2111.735 724.300 2112.250 724.440 ;
        RECT 2111.930 724.240 2112.250 724.300 ;
        RECT 2111.930 689.760 2112.250 689.820 ;
        RECT 2111.735 689.620 2112.250 689.760 ;
        RECT 2111.930 689.560 2112.250 689.620 ;
        RECT 2111.470 641.820 2111.790 641.880 ;
        RECT 2112.390 641.820 2112.710 641.880 ;
        RECT 2111.470 641.680 2112.710 641.820 ;
        RECT 2111.470 641.620 2111.790 641.680 ;
        RECT 2112.390 641.620 2112.710 641.680 ;
        RECT 2111.930 627.880 2112.250 627.940 ;
        RECT 2111.735 627.740 2112.250 627.880 ;
        RECT 2111.930 627.680 2112.250 627.740 ;
        RECT 2111.930 593.200 2112.250 593.260 ;
        RECT 2111.735 593.060 2112.250 593.200 ;
        RECT 2111.930 593.000 2112.250 593.060 ;
        RECT 2111.470 545.260 2111.790 545.320 ;
        RECT 2112.390 545.260 2112.710 545.320 ;
        RECT 2111.470 545.120 2112.710 545.260 ;
        RECT 2111.470 545.060 2111.790 545.120 ;
        RECT 2112.390 545.060 2112.710 545.120 ;
        RECT 2111.930 531.320 2112.250 531.380 ;
        RECT 2111.735 531.180 2112.250 531.320 ;
        RECT 2111.930 531.120 2112.250 531.180 ;
        RECT 2111.930 496.640 2112.250 496.700 ;
        RECT 2111.735 496.500 2112.250 496.640 ;
        RECT 2111.930 496.440 2112.250 496.500 ;
        RECT 2111.470 448.700 2111.790 448.760 ;
        RECT 2112.390 448.700 2112.710 448.760 ;
        RECT 2111.470 448.560 2112.710 448.700 ;
        RECT 2111.470 448.500 2111.790 448.560 ;
        RECT 2112.390 448.500 2112.710 448.560 ;
        RECT 2111.930 434.760 2112.250 434.820 ;
        RECT 2111.735 434.620 2112.250 434.760 ;
        RECT 2111.930 434.560 2112.250 434.620 ;
        RECT 2111.945 386.480 2112.235 386.525 ;
        RECT 2112.390 386.480 2112.710 386.540 ;
        RECT 2111.945 386.340 2112.710 386.480 ;
        RECT 2111.945 386.295 2112.235 386.340 ;
        RECT 2112.390 386.280 2112.710 386.340 ;
        RECT 2111.930 241.640 2112.250 241.700 ;
        RECT 2112.390 241.640 2112.710 241.700 ;
        RECT 2111.930 241.500 2112.710 241.640 ;
        RECT 2111.930 241.440 2112.250 241.500 ;
        RECT 2112.390 241.440 2112.710 241.500 ;
        RECT 2112.390 193.020 2112.710 193.080 ;
        RECT 2112.195 192.880 2112.710 193.020 ;
        RECT 2112.390 192.820 2112.710 192.880 ;
        RECT 2111.930 138.280 2112.250 138.340 ;
        RECT 2112.405 138.280 2112.695 138.325 ;
        RECT 2111.930 138.140 2112.695 138.280 ;
        RECT 2111.930 138.080 2112.250 138.140 ;
        RECT 2112.405 138.095 2112.695 138.140 ;
        RECT 2110.550 96.120 2110.870 96.180 ;
        RECT 2112.390 96.120 2112.710 96.180 ;
        RECT 2110.550 95.980 2112.710 96.120 ;
        RECT 2110.550 95.920 2110.870 95.980 ;
        RECT 2112.390 95.920 2112.710 95.980 ;
        RECT 2111.470 48.520 2111.790 48.580 ;
        RECT 2112.390 48.520 2112.710 48.580 ;
        RECT 2111.470 48.380 2112.710 48.520 ;
        RECT 2111.470 48.320 2111.790 48.380 ;
        RECT 2112.390 48.320 2112.710 48.380 ;
        RECT 1881.930 25.400 1882.250 25.460 ;
        RECT 2111.470 25.400 2111.790 25.460 ;
        RECT 1881.930 25.260 2111.790 25.400 ;
        RECT 1881.930 25.200 1882.250 25.260 ;
        RECT 2111.470 25.200 2111.790 25.260 ;
      LAYER via ;
        RECT 2111.500 1677.940 2111.760 1678.200 ;
        RECT 2116.100 1677.940 2116.360 1678.200 ;
        RECT 2111.500 1655.840 2111.760 1656.100 ;
        RECT 2112.420 1655.840 2112.680 1656.100 ;
        RECT 2112.420 1641.900 2112.680 1642.160 ;
        RECT 2111.960 1593.960 2112.220 1594.220 ;
        RECT 2111.500 1558.940 2111.760 1559.200 ;
        RECT 2112.420 1558.940 2112.680 1559.200 ;
        RECT 2112.420 1545.340 2112.680 1545.600 ;
        RECT 2112.420 1499.440 2112.680 1499.700 ;
        RECT 2111.500 1414.440 2111.760 1414.700 ;
        RECT 2112.420 1414.440 2112.680 1414.700 ;
        RECT 2111.500 1317.880 2111.760 1318.140 ;
        RECT 2112.420 1317.880 2112.680 1318.140 ;
        RECT 2111.500 1221.320 2111.760 1221.580 ;
        RECT 2112.420 1221.320 2112.680 1221.580 ;
        RECT 2111.500 1124.760 2111.760 1125.020 ;
        RECT 2112.420 1124.760 2112.680 1125.020 ;
        RECT 2111.500 1028.200 2111.760 1028.460 ;
        RECT 2112.420 1028.200 2112.680 1028.460 ;
        RECT 2111.500 931.640 2111.760 931.900 ;
        RECT 2112.420 931.640 2112.680 931.900 ;
        RECT 2112.420 869.420 2112.680 869.680 ;
        RECT 2113.340 869.420 2113.600 869.680 ;
        RECT 2111.500 835.080 2111.760 835.340 ;
        RECT 2112.420 835.080 2112.680 835.340 ;
        RECT 2111.960 820.800 2112.220 821.060 ;
        RECT 2111.960 786.460 2112.220 786.720 ;
        RECT 2111.500 738.180 2111.760 738.440 ;
        RECT 2112.420 738.180 2112.680 738.440 ;
        RECT 2111.960 724.240 2112.220 724.500 ;
        RECT 2111.960 689.560 2112.220 689.820 ;
        RECT 2111.500 641.620 2111.760 641.880 ;
        RECT 2112.420 641.620 2112.680 641.880 ;
        RECT 2111.960 627.680 2112.220 627.940 ;
        RECT 2111.960 593.000 2112.220 593.260 ;
        RECT 2111.500 545.060 2111.760 545.320 ;
        RECT 2112.420 545.060 2112.680 545.320 ;
        RECT 2111.960 531.120 2112.220 531.380 ;
        RECT 2111.960 496.440 2112.220 496.700 ;
        RECT 2111.500 448.500 2111.760 448.760 ;
        RECT 2112.420 448.500 2112.680 448.760 ;
        RECT 2111.960 434.560 2112.220 434.820 ;
        RECT 2112.420 386.280 2112.680 386.540 ;
        RECT 2111.960 241.440 2112.220 241.700 ;
        RECT 2112.420 241.440 2112.680 241.700 ;
        RECT 2112.420 192.820 2112.680 193.080 ;
        RECT 2111.960 138.080 2112.220 138.340 ;
        RECT 2110.580 95.920 2110.840 96.180 ;
        RECT 2112.420 95.920 2112.680 96.180 ;
        RECT 2111.500 48.320 2111.760 48.580 ;
        RECT 2112.420 48.320 2112.680 48.580 ;
        RECT 1881.960 25.200 1882.220 25.460 ;
        RECT 2111.500 25.200 2111.760 25.460 ;
      LAYER met2 ;
        RECT 2117.400 1700.410 2117.680 1702.400 ;
        RECT 2116.160 1700.270 2117.680 1700.410 ;
        RECT 2116.160 1678.230 2116.300 1700.270 ;
        RECT 2117.400 1700.000 2117.680 1700.270 ;
        RECT 2111.500 1677.910 2111.760 1678.230 ;
        RECT 2116.100 1677.910 2116.360 1678.230 ;
        RECT 2111.560 1656.130 2111.700 1677.910 ;
        RECT 2111.500 1655.810 2111.760 1656.130 ;
        RECT 2112.420 1655.810 2112.680 1656.130 ;
        RECT 2112.480 1642.190 2112.620 1655.810 ;
        RECT 2112.420 1641.870 2112.680 1642.190 ;
        RECT 2111.960 1593.930 2112.220 1594.250 ;
        RECT 2112.020 1559.650 2112.160 1593.930 ;
        RECT 2111.560 1559.510 2112.160 1559.650 ;
        RECT 2111.560 1559.230 2111.700 1559.510 ;
        RECT 2111.500 1558.910 2111.760 1559.230 ;
        RECT 2112.420 1558.910 2112.680 1559.230 ;
        RECT 2112.480 1545.630 2112.620 1558.910 ;
        RECT 2112.420 1545.310 2112.680 1545.630 ;
        RECT 2112.420 1499.410 2112.680 1499.730 ;
        RECT 2112.480 1414.730 2112.620 1499.410 ;
        RECT 2111.500 1414.410 2111.760 1414.730 ;
        RECT 2112.420 1414.410 2112.680 1414.730 ;
        RECT 2111.560 1414.130 2111.700 1414.410 ;
        RECT 2111.560 1413.990 2112.160 1414.130 ;
        RECT 2112.020 1366.530 2112.160 1413.990 ;
        RECT 2112.020 1366.390 2112.620 1366.530 ;
        RECT 2112.480 1318.170 2112.620 1366.390 ;
        RECT 2111.500 1317.850 2111.760 1318.170 ;
        RECT 2112.420 1317.850 2112.680 1318.170 ;
        RECT 2111.560 1317.570 2111.700 1317.850 ;
        RECT 2111.560 1317.430 2112.160 1317.570 ;
        RECT 2112.020 1269.970 2112.160 1317.430 ;
        RECT 2112.020 1269.830 2112.620 1269.970 ;
        RECT 2112.480 1221.610 2112.620 1269.830 ;
        RECT 2111.500 1221.290 2111.760 1221.610 ;
        RECT 2112.420 1221.290 2112.680 1221.610 ;
        RECT 2111.560 1221.010 2111.700 1221.290 ;
        RECT 2111.560 1220.870 2112.160 1221.010 ;
        RECT 2112.020 1173.410 2112.160 1220.870 ;
        RECT 2112.020 1173.270 2112.620 1173.410 ;
        RECT 2112.480 1125.050 2112.620 1173.270 ;
        RECT 2111.500 1124.730 2111.760 1125.050 ;
        RECT 2112.420 1124.730 2112.680 1125.050 ;
        RECT 2111.560 1124.450 2111.700 1124.730 ;
        RECT 2111.560 1124.310 2112.160 1124.450 ;
        RECT 2112.020 1076.850 2112.160 1124.310 ;
        RECT 2112.020 1076.710 2112.620 1076.850 ;
        RECT 2112.480 1028.490 2112.620 1076.710 ;
        RECT 2111.500 1028.170 2111.760 1028.490 ;
        RECT 2112.420 1028.170 2112.680 1028.490 ;
        RECT 2111.560 1027.890 2111.700 1028.170 ;
        RECT 2111.560 1027.750 2112.160 1027.890 ;
        RECT 2112.020 980.290 2112.160 1027.750 ;
        RECT 2112.020 980.150 2112.620 980.290 ;
        RECT 2112.480 931.930 2112.620 980.150 ;
        RECT 2111.500 931.610 2111.760 931.930 ;
        RECT 2112.420 931.610 2112.680 931.930 ;
        RECT 2111.560 931.330 2111.700 931.610 ;
        RECT 2111.560 931.190 2112.160 931.330 ;
        RECT 2112.020 917.845 2112.160 931.190 ;
        RECT 2111.950 917.475 2112.230 917.845 ;
        RECT 2113.330 917.475 2113.610 917.845 ;
        RECT 2113.400 869.710 2113.540 917.475 ;
        RECT 2112.420 869.390 2112.680 869.710 ;
        RECT 2113.340 869.390 2113.600 869.710 ;
        RECT 2112.480 835.370 2112.620 869.390 ;
        RECT 2111.500 835.050 2111.760 835.370 ;
        RECT 2112.420 835.050 2112.680 835.370 ;
        RECT 2111.560 834.770 2111.700 835.050 ;
        RECT 2111.560 834.630 2112.160 834.770 ;
        RECT 2112.020 821.090 2112.160 834.630 ;
        RECT 2111.960 820.770 2112.220 821.090 ;
        RECT 2111.960 786.430 2112.220 786.750 ;
        RECT 2112.020 772.890 2112.160 786.430 ;
        RECT 2112.020 772.750 2112.620 772.890 ;
        RECT 2112.480 738.470 2112.620 772.750 ;
        RECT 2111.500 738.210 2111.760 738.470 ;
        RECT 2111.500 738.150 2112.160 738.210 ;
        RECT 2112.420 738.150 2112.680 738.470 ;
        RECT 2111.560 738.070 2112.160 738.150 ;
        RECT 2112.020 724.530 2112.160 738.070 ;
        RECT 2111.960 724.210 2112.220 724.530 ;
        RECT 2111.960 689.530 2112.220 689.850 ;
        RECT 2112.020 676.330 2112.160 689.530 ;
        RECT 2112.020 676.190 2112.620 676.330 ;
        RECT 2112.480 641.910 2112.620 676.190 ;
        RECT 2111.500 641.650 2111.760 641.910 ;
        RECT 2111.500 641.590 2112.160 641.650 ;
        RECT 2112.420 641.590 2112.680 641.910 ;
        RECT 2111.560 641.510 2112.160 641.590 ;
        RECT 2112.020 627.970 2112.160 641.510 ;
        RECT 2111.960 627.650 2112.220 627.970 ;
        RECT 2111.960 592.970 2112.220 593.290 ;
        RECT 2112.020 579.770 2112.160 592.970 ;
        RECT 2112.020 579.630 2112.620 579.770 ;
        RECT 2112.480 545.350 2112.620 579.630 ;
        RECT 2111.500 545.090 2111.760 545.350 ;
        RECT 2111.500 545.030 2112.160 545.090 ;
        RECT 2112.420 545.030 2112.680 545.350 ;
        RECT 2111.560 544.950 2112.160 545.030 ;
        RECT 2112.020 531.410 2112.160 544.950 ;
        RECT 2111.960 531.090 2112.220 531.410 ;
        RECT 2111.960 496.410 2112.220 496.730 ;
        RECT 2112.020 483.210 2112.160 496.410 ;
        RECT 2112.020 483.070 2112.620 483.210 ;
        RECT 2112.480 448.790 2112.620 483.070 ;
        RECT 2111.500 448.530 2111.760 448.790 ;
        RECT 2111.500 448.470 2112.160 448.530 ;
        RECT 2112.420 448.470 2112.680 448.790 ;
        RECT 2111.560 448.390 2112.160 448.470 ;
        RECT 2112.020 434.850 2112.160 448.390 ;
        RECT 2111.960 434.530 2112.220 434.850 ;
        RECT 2112.420 386.250 2112.680 386.570 ;
        RECT 2112.480 351.290 2112.620 386.250 ;
        RECT 2112.020 351.150 2112.620 351.290 ;
        RECT 2112.020 303.690 2112.160 351.150 ;
        RECT 2112.020 303.550 2112.620 303.690 ;
        RECT 2112.480 241.730 2112.620 303.550 ;
        RECT 2111.960 241.410 2112.220 241.730 ;
        RECT 2112.420 241.410 2112.680 241.730 ;
        RECT 2112.020 207.130 2112.160 241.410 ;
        RECT 2112.020 206.990 2112.620 207.130 ;
        RECT 2112.480 193.110 2112.620 206.990 ;
        RECT 2112.420 192.790 2112.680 193.110 ;
        RECT 2111.960 138.050 2112.220 138.370 ;
        RECT 2110.570 137.515 2110.850 137.885 ;
        RECT 2111.490 137.770 2111.770 137.885 ;
        RECT 2112.020 137.770 2112.160 138.050 ;
        RECT 2111.490 137.630 2112.160 137.770 ;
        RECT 2111.490 137.515 2111.770 137.630 ;
        RECT 2110.640 96.210 2110.780 137.515 ;
        RECT 2110.580 95.890 2110.840 96.210 ;
        RECT 2112.420 95.890 2112.680 96.210 ;
        RECT 2112.480 48.610 2112.620 95.890 ;
        RECT 2111.500 48.290 2111.760 48.610 ;
        RECT 2112.420 48.290 2112.680 48.610 ;
        RECT 2111.560 25.490 2111.700 48.290 ;
        RECT 1881.960 25.170 1882.220 25.490 ;
        RECT 2111.500 25.170 2111.760 25.490 ;
        RECT 1882.020 2.400 1882.160 25.170 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
      LAYER via2 ;
        RECT 2111.950 917.520 2112.230 917.800 ;
        RECT 2113.330 917.520 2113.610 917.800 ;
        RECT 2110.570 137.560 2110.850 137.840 ;
        RECT 2111.490 137.560 2111.770 137.840 ;
      LAYER met3 ;
        RECT 2111.925 917.810 2112.255 917.825 ;
        RECT 2113.305 917.810 2113.635 917.825 ;
        RECT 2111.925 917.510 2113.635 917.810 ;
        RECT 2111.925 917.495 2112.255 917.510 ;
        RECT 2113.305 917.495 2113.635 917.510 ;
        RECT 2110.545 137.850 2110.875 137.865 ;
        RECT 2111.465 137.850 2111.795 137.865 ;
        RECT 2110.545 137.550 2111.795 137.850 ;
        RECT 2110.545 137.535 2110.875 137.550 ;
        RECT 2111.465 137.535 2111.795 137.550 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1899.870 31.180 1900.190 31.240 ;
        RECT 2125.730 31.180 2126.050 31.240 ;
        RECT 1899.870 31.040 2126.050 31.180 ;
        RECT 1899.870 30.980 1900.190 31.040 ;
        RECT 2125.730 30.980 2126.050 31.040 ;
      LAYER via ;
        RECT 1899.900 30.980 1900.160 31.240 ;
        RECT 2125.760 30.980 2126.020 31.240 ;
      LAYER met2 ;
        RECT 2126.140 1700.410 2126.420 1702.400 ;
        RECT 2125.820 1700.270 2126.420 1700.410 ;
        RECT 2125.820 31.270 2125.960 1700.270 ;
        RECT 2126.140 1700.000 2126.420 1700.270 ;
        RECT 1899.900 30.950 1900.160 31.270 ;
        RECT 2125.760 30.950 2126.020 31.270 ;
        RECT 1899.960 2.400 1900.100 30.950 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1917.810 25.740 1918.130 25.800 ;
        RECT 2133.550 25.740 2133.870 25.800 ;
        RECT 1917.810 25.600 2133.870 25.740 ;
        RECT 1917.810 25.540 1918.130 25.600 ;
        RECT 2133.550 25.540 2133.870 25.600 ;
      LAYER via ;
        RECT 1917.840 25.540 1918.100 25.800 ;
        RECT 2133.580 25.540 2133.840 25.800 ;
      LAYER met2 ;
        RECT 2135.340 1700.410 2135.620 1702.400 ;
        RECT 2133.640 1700.270 2135.620 1700.410 ;
        RECT 2133.640 25.830 2133.780 1700.270 ;
        RECT 2135.340 1700.000 2135.620 1700.270 ;
        RECT 1917.840 25.510 1918.100 25.830 ;
        RECT 2133.580 25.510 2133.840 25.830 ;
        RECT 1917.900 2.400 1918.040 25.510 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2139.605 1594.005 2139.775 1642.115 ;
        RECT 2140.065 1497.445 2140.235 1545.555 ;
        RECT 2139.605 869.465 2139.775 883.575 ;
        RECT 2139.605 786.505 2139.775 821.015 ;
        RECT 2139.605 676.345 2139.775 690.455 ;
        RECT 2139.605 593.045 2139.775 627.895 ;
        RECT 2139.605 496.485 2139.775 531.335 ;
        RECT 2139.605 386.325 2139.775 434.775 ;
      LAYER mcon ;
        RECT 2139.605 1641.945 2139.775 1642.115 ;
        RECT 2140.065 1545.385 2140.235 1545.555 ;
        RECT 2139.605 883.405 2139.775 883.575 ;
        RECT 2139.605 820.845 2139.775 821.015 ;
        RECT 2139.605 690.285 2139.775 690.455 ;
        RECT 2139.605 627.725 2139.775 627.895 ;
        RECT 2139.605 531.165 2139.775 531.335 ;
        RECT 2139.605 434.605 2139.775 434.775 ;
      LAYER met1 ;
        RECT 2139.545 1642.100 2139.835 1642.145 ;
        RECT 2139.990 1642.100 2140.310 1642.160 ;
        RECT 2139.545 1641.960 2140.310 1642.100 ;
        RECT 2139.545 1641.915 2139.835 1641.960 ;
        RECT 2139.990 1641.900 2140.310 1641.960 ;
        RECT 2139.530 1594.160 2139.850 1594.220 ;
        RECT 2139.335 1594.020 2139.850 1594.160 ;
        RECT 2139.530 1593.960 2139.850 1594.020 ;
        RECT 2139.070 1559.140 2139.390 1559.200 ;
        RECT 2139.990 1559.140 2140.310 1559.200 ;
        RECT 2139.070 1559.000 2140.310 1559.140 ;
        RECT 2139.070 1558.940 2139.390 1559.000 ;
        RECT 2139.990 1558.940 2140.310 1559.000 ;
        RECT 2139.990 1545.540 2140.310 1545.600 ;
        RECT 2139.795 1545.400 2140.310 1545.540 ;
        RECT 2139.990 1545.340 2140.310 1545.400 ;
        RECT 2139.990 1497.600 2140.310 1497.660 ;
        RECT 2139.795 1497.460 2140.310 1497.600 ;
        RECT 2139.990 1497.400 2140.310 1497.460 ;
        RECT 2139.070 1414.640 2139.390 1414.700 ;
        RECT 2139.990 1414.640 2140.310 1414.700 ;
        RECT 2139.070 1414.500 2140.310 1414.640 ;
        RECT 2139.070 1414.440 2139.390 1414.500 ;
        RECT 2139.990 1414.440 2140.310 1414.500 ;
        RECT 2139.070 1318.080 2139.390 1318.140 ;
        RECT 2139.990 1318.080 2140.310 1318.140 ;
        RECT 2139.070 1317.940 2140.310 1318.080 ;
        RECT 2139.070 1317.880 2139.390 1317.940 ;
        RECT 2139.990 1317.880 2140.310 1317.940 ;
        RECT 2139.070 1221.520 2139.390 1221.580 ;
        RECT 2139.990 1221.520 2140.310 1221.580 ;
        RECT 2139.070 1221.380 2140.310 1221.520 ;
        RECT 2139.070 1221.320 2139.390 1221.380 ;
        RECT 2139.990 1221.320 2140.310 1221.380 ;
        RECT 2139.070 1124.960 2139.390 1125.020 ;
        RECT 2139.990 1124.960 2140.310 1125.020 ;
        RECT 2139.070 1124.820 2140.310 1124.960 ;
        RECT 2139.070 1124.760 2139.390 1124.820 ;
        RECT 2139.990 1124.760 2140.310 1124.820 ;
        RECT 2139.070 1028.400 2139.390 1028.460 ;
        RECT 2139.990 1028.400 2140.310 1028.460 ;
        RECT 2139.070 1028.260 2140.310 1028.400 ;
        RECT 2139.070 1028.200 2139.390 1028.260 ;
        RECT 2139.990 1028.200 2140.310 1028.260 ;
        RECT 2139.530 883.560 2139.850 883.620 ;
        RECT 2139.335 883.420 2139.850 883.560 ;
        RECT 2139.530 883.360 2139.850 883.420 ;
        RECT 2139.530 869.620 2139.850 869.680 ;
        RECT 2139.335 869.480 2139.850 869.620 ;
        RECT 2139.530 869.420 2139.850 869.480 ;
        RECT 2139.530 821.000 2139.850 821.060 ;
        RECT 2139.335 820.860 2139.850 821.000 ;
        RECT 2139.530 820.800 2139.850 820.860 ;
        RECT 2139.530 786.660 2139.850 786.720 ;
        RECT 2139.335 786.520 2139.850 786.660 ;
        RECT 2139.530 786.460 2139.850 786.520 ;
        RECT 2139.070 738.380 2139.390 738.440 ;
        RECT 2139.990 738.380 2140.310 738.440 ;
        RECT 2139.070 738.240 2140.310 738.380 ;
        RECT 2139.070 738.180 2139.390 738.240 ;
        RECT 2139.990 738.180 2140.310 738.240 ;
        RECT 2139.545 690.440 2139.835 690.485 ;
        RECT 2139.990 690.440 2140.310 690.500 ;
        RECT 2139.545 690.300 2140.310 690.440 ;
        RECT 2139.545 690.255 2139.835 690.300 ;
        RECT 2139.990 690.240 2140.310 690.300 ;
        RECT 2139.530 676.500 2139.850 676.560 ;
        RECT 2139.335 676.360 2139.850 676.500 ;
        RECT 2139.530 676.300 2139.850 676.360 ;
        RECT 2139.530 627.880 2139.850 627.940 ;
        RECT 2139.335 627.740 2139.850 627.880 ;
        RECT 2139.530 627.680 2139.850 627.740 ;
        RECT 2139.530 593.200 2139.850 593.260 ;
        RECT 2139.335 593.060 2139.850 593.200 ;
        RECT 2139.530 593.000 2139.850 593.060 ;
        RECT 2139.070 545.260 2139.390 545.320 ;
        RECT 2139.990 545.260 2140.310 545.320 ;
        RECT 2139.070 545.120 2140.310 545.260 ;
        RECT 2139.070 545.060 2139.390 545.120 ;
        RECT 2139.990 545.060 2140.310 545.120 ;
        RECT 2139.530 531.320 2139.850 531.380 ;
        RECT 2139.335 531.180 2139.850 531.320 ;
        RECT 2139.530 531.120 2139.850 531.180 ;
        RECT 2139.530 496.640 2139.850 496.700 ;
        RECT 2139.335 496.500 2139.850 496.640 ;
        RECT 2139.530 496.440 2139.850 496.500 ;
        RECT 2139.070 448.700 2139.390 448.760 ;
        RECT 2139.990 448.700 2140.310 448.760 ;
        RECT 2139.070 448.560 2140.310 448.700 ;
        RECT 2139.070 448.500 2139.390 448.560 ;
        RECT 2139.990 448.500 2140.310 448.560 ;
        RECT 2139.530 434.760 2139.850 434.820 ;
        RECT 2139.335 434.620 2139.850 434.760 ;
        RECT 2139.530 434.560 2139.850 434.620 ;
        RECT 2139.545 386.480 2139.835 386.525 ;
        RECT 2139.990 386.480 2140.310 386.540 ;
        RECT 2139.545 386.340 2140.310 386.480 ;
        RECT 2139.545 386.295 2139.835 386.340 ;
        RECT 2139.990 386.280 2140.310 386.340 ;
        RECT 2139.530 159.020 2139.850 159.080 ;
        RECT 2139.160 158.880 2139.850 159.020 ;
        RECT 2139.160 158.740 2139.300 158.880 ;
        RECT 2139.530 158.820 2139.850 158.880 ;
        RECT 2139.070 158.480 2139.390 158.740 ;
        RECT 2139.530 61.780 2139.850 61.840 ;
        RECT 2140.450 61.780 2140.770 61.840 ;
        RECT 2139.530 61.640 2140.770 61.780 ;
        RECT 2139.530 61.580 2139.850 61.640 ;
        RECT 2140.450 61.580 2140.770 61.640 ;
        RECT 1935.290 26.080 1935.610 26.140 ;
        RECT 2139.530 26.080 2139.850 26.140 ;
        RECT 1935.290 25.940 2139.850 26.080 ;
        RECT 1935.290 25.880 1935.610 25.940 ;
        RECT 2139.530 25.880 2139.850 25.940 ;
      LAYER via ;
        RECT 2140.020 1641.900 2140.280 1642.160 ;
        RECT 2139.560 1593.960 2139.820 1594.220 ;
        RECT 2139.100 1558.940 2139.360 1559.200 ;
        RECT 2140.020 1558.940 2140.280 1559.200 ;
        RECT 2140.020 1545.340 2140.280 1545.600 ;
        RECT 2140.020 1497.400 2140.280 1497.660 ;
        RECT 2139.100 1414.440 2139.360 1414.700 ;
        RECT 2140.020 1414.440 2140.280 1414.700 ;
        RECT 2139.100 1317.880 2139.360 1318.140 ;
        RECT 2140.020 1317.880 2140.280 1318.140 ;
        RECT 2139.100 1221.320 2139.360 1221.580 ;
        RECT 2140.020 1221.320 2140.280 1221.580 ;
        RECT 2139.100 1124.760 2139.360 1125.020 ;
        RECT 2140.020 1124.760 2140.280 1125.020 ;
        RECT 2139.100 1028.200 2139.360 1028.460 ;
        RECT 2140.020 1028.200 2140.280 1028.460 ;
        RECT 2139.560 883.360 2139.820 883.620 ;
        RECT 2139.560 869.420 2139.820 869.680 ;
        RECT 2139.560 820.800 2139.820 821.060 ;
        RECT 2139.560 786.460 2139.820 786.720 ;
        RECT 2139.100 738.180 2139.360 738.440 ;
        RECT 2140.020 738.180 2140.280 738.440 ;
        RECT 2140.020 690.240 2140.280 690.500 ;
        RECT 2139.560 676.300 2139.820 676.560 ;
        RECT 2139.560 627.680 2139.820 627.940 ;
        RECT 2139.560 593.000 2139.820 593.260 ;
        RECT 2139.100 545.060 2139.360 545.320 ;
        RECT 2140.020 545.060 2140.280 545.320 ;
        RECT 2139.560 531.120 2139.820 531.380 ;
        RECT 2139.560 496.440 2139.820 496.700 ;
        RECT 2139.100 448.500 2139.360 448.760 ;
        RECT 2140.020 448.500 2140.280 448.760 ;
        RECT 2139.560 434.560 2139.820 434.820 ;
        RECT 2140.020 386.280 2140.280 386.540 ;
        RECT 2139.560 158.820 2139.820 159.080 ;
        RECT 2139.100 158.480 2139.360 158.740 ;
        RECT 2139.560 61.580 2139.820 61.840 ;
        RECT 2140.480 61.580 2140.740 61.840 ;
        RECT 1935.320 25.880 1935.580 26.140 ;
        RECT 2139.560 25.880 2139.820 26.140 ;
      LAYER met2 ;
        RECT 2144.540 1700.410 2144.820 1702.400 ;
        RECT 2142.380 1700.270 2144.820 1700.410 ;
        RECT 2142.380 1656.890 2142.520 1700.270 ;
        RECT 2144.540 1700.000 2144.820 1700.270 ;
        RECT 2141.920 1656.750 2142.520 1656.890 ;
        RECT 2141.920 1643.405 2142.060 1656.750 ;
        RECT 2141.850 1643.035 2142.130 1643.405 ;
        RECT 2140.010 1642.355 2140.290 1642.725 ;
        RECT 2140.080 1642.190 2140.220 1642.355 ;
        RECT 2140.020 1641.870 2140.280 1642.190 ;
        RECT 2139.560 1593.930 2139.820 1594.250 ;
        RECT 2139.620 1559.650 2139.760 1593.930 ;
        RECT 2139.160 1559.510 2139.760 1559.650 ;
        RECT 2139.160 1559.230 2139.300 1559.510 ;
        RECT 2139.100 1558.910 2139.360 1559.230 ;
        RECT 2140.020 1558.910 2140.280 1559.230 ;
        RECT 2140.080 1545.630 2140.220 1558.910 ;
        RECT 2140.020 1545.310 2140.280 1545.630 ;
        RECT 2140.020 1497.370 2140.280 1497.690 ;
        RECT 2140.080 1414.730 2140.220 1497.370 ;
        RECT 2139.100 1414.410 2139.360 1414.730 ;
        RECT 2140.020 1414.410 2140.280 1414.730 ;
        RECT 2139.160 1414.130 2139.300 1414.410 ;
        RECT 2139.160 1413.990 2139.760 1414.130 ;
        RECT 2139.620 1366.530 2139.760 1413.990 ;
        RECT 2139.620 1366.390 2140.220 1366.530 ;
        RECT 2140.080 1318.170 2140.220 1366.390 ;
        RECT 2139.100 1317.850 2139.360 1318.170 ;
        RECT 2140.020 1317.850 2140.280 1318.170 ;
        RECT 2139.160 1317.570 2139.300 1317.850 ;
        RECT 2139.160 1317.430 2139.760 1317.570 ;
        RECT 2139.620 1269.970 2139.760 1317.430 ;
        RECT 2139.620 1269.830 2140.220 1269.970 ;
        RECT 2140.080 1221.610 2140.220 1269.830 ;
        RECT 2139.100 1221.290 2139.360 1221.610 ;
        RECT 2140.020 1221.290 2140.280 1221.610 ;
        RECT 2139.160 1221.010 2139.300 1221.290 ;
        RECT 2139.160 1220.870 2139.760 1221.010 ;
        RECT 2139.620 1173.410 2139.760 1220.870 ;
        RECT 2139.620 1173.270 2140.220 1173.410 ;
        RECT 2140.080 1125.050 2140.220 1173.270 ;
        RECT 2139.100 1124.730 2139.360 1125.050 ;
        RECT 2140.020 1124.730 2140.280 1125.050 ;
        RECT 2139.160 1124.450 2139.300 1124.730 ;
        RECT 2139.160 1124.310 2139.760 1124.450 ;
        RECT 2139.620 1076.850 2139.760 1124.310 ;
        RECT 2139.620 1076.710 2140.220 1076.850 ;
        RECT 2140.080 1028.490 2140.220 1076.710 ;
        RECT 2139.100 1028.170 2139.360 1028.490 ;
        RECT 2140.020 1028.170 2140.280 1028.490 ;
        RECT 2139.160 1027.890 2139.300 1028.170 ;
        RECT 2139.160 1027.750 2139.760 1027.890 ;
        RECT 2139.620 980.290 2139.760 1027.750 ;
        RECT 2139.620 980.150 2140.220 980.290 ;
        RECT 2140.080 917.730 2140.220 980.150 ;
        RECT 2139.620 917.590 2140.220 917.730 ;
        RECT 2139.620 883.650 2139.760 917.590 ;
        RECT 2139.560 883.330 2139.820 883.650 ;
        RECT 2139.560 869.390 2139.820 869.710 ;
        RECT 2139.620 835.450 2139.760 869.390 ;
        RECT 2139.160 835.310 2139.760 835.450 ;
        RECT 2139.160 834.770 2139.300 835.310 ;
        RECT 2139.160 834.630 2139.760 834.770 ;
        RECT 2139.620 821.090 2139.760 834.630 ;
        RECT 2139.560 820.770 2139.820 821.090 ;
        RECT 2139.560 786.430 2139.820 786.750 ;
        RECT 2139.620 772.890 2139.760 786.430 ;
        RECT 2139.620 772.750 2140.220 772.890 ;
        RECT 2140.080 738.470 2140.220 772.750 ;
        RECT 2139.100 738.210 2139.360 738.470 ;
        RECT 2140.020 738.210 2140.280 738.470 ;
        RECT 2139.100 738.150 2140.280 738.210 ;
        RECT 2139.160 738.070 2140.220 738.150 ;
        RECT 2140.080 690.530 2140.220 738.070 ;
        RECT 2140.020 690.210 2140.280 690.530 ;
        RECT 2139.560 676.270 2139.820 676.590 ;
        RECT 2139.620 642.330 2139.760 676.270 ;
        RECT 2139.160 642.190 2139.760 642.330 ;
        RECT 2139.160 641.650 2139.300 642.190 ;
        RECT 2139.160 641.510 2139.760 641.650 ;
        RECT 2139.620 627.970 2139.760 641.510 ;
        RECT 2139.560 627.650 2139.820 627.970 ;
        RECT 2139.560 592.970 2139.820 593.290 ;
        RECT 2139.620 579.770 2139.760 592.970 ;
        RECT 2139.620 579.630 2140.220 579.770 ;
        RECT 2140.080 545.350 2140.220 579.630 ;
        RECT 2139.100 545.090 2139.360 545.350 ;
        RECT 2139.100 545.030 2139.760 545.090 ;
        RECT 2140.020 545.030 2140.280 545.350 ;
        RECT 2139.160 544.950 2139.760 545.030 ;
        RECT 2139.620 531.410 2139.760 544.950 ;
        RECT 2139.560 531.090 2139.820 531.410 ;
        RECT 2139.560 496.410 2139.820 496.730 ;
        RECT 2139.620 483.210 2139.760 496.410 ;
        RECT 2139.620 483.070 2140.220 483.210 ;
        RECT 2140.080 448.790 2140.220 483.070 ;
        RECT 2139.100 448.530 2139.360 448.790 ;
        RECT 2139.100 448.470 2139.760 448.530 ;
        RECT 2140.020 448.470 2140.280 448.790 ;
        RECT 2139.160 448.390 2139.760 448.470 ;
        RECT 2139.620 434.850 2139.760 448.390 ;
        RECT 2139.560 434.530 2139.820 434.850 ;
        RECT 2140.020 386.250 2140.280 386.570 ;
        RECT 2140.080 351.290 2140.220 386.250 ;
        RECT 2139.620 351.150 2140.220 351.290 ;
        RECT 2139.620 303.690 2139.760 351.150 ;
        RECT 2139.620 303.550 2140.220 303.690 ;
        RECT 2140.080 255.410 2140.220 303.550 ;
        RECT 2139.160 255.270 2140.220 255.410 ;
        RECT 2139.160 254.730 2139.300 255.270 ;
        RECT 2139.160 254.590 2139.760 254.730 ;
        RECT 2139.620 159.110 2139.760 254.590 ;
        RECT 2139.560 158.790 2139.820 159.110 ;
        RECT 2139.100 158.450 2139.360 158.770 ;
        RECT 2139.160 131.650 2139.300 158.450 ;
        RECT 2139.160 131.510 2139.760 131.650 ;
        RECT 2139.620 124.285 2139.760 131.510 ;
        RECT 2139.550 123.915 2139.830 124.285 ;
        RECT 2140.470 123.915 2140.750 124.285 ;
        RECT 2140.540 61.870 2140.680 123.915 ;
        RECT 2139.560 61.550 2139.820 61.870 ;
        RECT 2140.480 61.550 2140.740 61.870 ;
        RECT 2139.620 26.170 2139.760 61.550 ;
        RECT 1935.320 25.850 1935.580 26.170 ;
        RECT 2139.560 25.850 2139.820 26.170 ;
        RECT 1935.380 2.400 1935.520 25.850 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
      LAYER via2 ;
        RECT 2141.850 1643.080 2142.130 1643.360 ;
        RECT 2140.010 1642.400 2140.290 1642.680 ;
        RECT 2139.550 123.960 2139.830 124.240 ;
        RECT 2140.470 123.960 2140.750 124.240 ;
      LAYER met3 ;
        RECT 2141.825 1643.370 2142.155 1643.385 ;
        RECT 2139.310 1643.070 2142.155 1643.370 ;
        RECT 2139.310 1642.690 2139.610 1643.070 ;
        RECT 2141.825 1643.055 2142.155 1643.070 ;
        RECT 2139.985 1642.690 2140.315 1642.705 ;
        RECT 2139.310 1642.390 2140.315 1642.690 ;
        RECT 2139.985 1642.375 2140.315 1642.390 ;
        RECT 2139.525 124.250 2139.855 124.265 ;
        RECT 2140.445 124.250 2140.775 124.265 ;
        RECT 2139.525 123.950 2140.775 124.250 ;
        RECT 2139.525 123.935 2139.855 123.950 ;
        RECT 2140.445 123.935 2140.775 123.950 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1953.230 26.420 1953.550 26.480 ;
        RECT 2153.330 26.420 2153.650 26.480 ;
        RECT 1953.230 26.280 2153.650 26.420 ;
        RECT 1953.230 26.220 1953.550 26.280 ;
        RECT 2153.330 26.220 2153.650 26.280 ;
      LAYER via ;
        RECT 1953.260 26.220 1953.520 26.480 ;
        RECT 2153.360 26.220 2153.620 26.480 ;
      LAYER met2 ;
        RECT 2153.740 1700.410 2154.020 1702.400 ;
        RECT 2153.420 1700.270 2154.020 1700.410 ;
        RECT 2153.420 26.510 2153.560 1700.270 ;
        RECT 2153.740 1700.000 2154.020 1700.270 ;
        RECT 1953.260 26.190 1953.520 26.510 ;
        RECT 2153.360 26.190 2153.620 26.510 ;
        RECT 1953.320 2.400 1953.460 26.190 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1971.170 26.760 1971.490 26.820 ;
        RECT 2160.690 26.760 2161.010 26.820 ;
        RECT 1971.170 26.620 2161.010 26.760 ;
        RECT 1971.170 26.560 1971.490 26.620 ;
        RECT 2160.690 26.560 2161.010 26.620 ;
      LAYER via ;
        RECT 1971.200 26.560 1971.460 26.820 ;
        RECT 2160.720 26.560 2160.980 26.820 ;
      LAYER met2 ;
        RECT 2162.940 1700.410 2163.220 1702.400 ;
        RECT 2160.780 1700.270 2163.220 1700.410 ;
        RECT 2160.780 26.850 2160.920 1700.270 ;
        RECT 2162.940 1700.000 2163.220 1700.270 ;
        RECT 1971.200 26.530 1971.460 26.850 ;
        RECT 2160.720 26.530 2160.980 26.850 ;
        RECT 1971.260 2.400 1971.400 26.530 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2168.585 1594.005 2168.755 1642.115 ;
        RECT 2167.205 1497.445 2167.375 1545.555 ;
        RECT 2168.125 1352.605 2168.295 1400.715 ;
        RECT 2168.125 1256.045 2168.295 1304.155 ;
        RECT 2168.125 869.465 2168.295 883.235 ;
        RECT 2168.125 593.045 2168.295 627.895 ;
        RECT 2167.205 386.325 2167.375 434.775 ;
        RECT 2168.125 241.485 2168.295 289.595 ;
        RECT 2168.125 186.745 2168.295 206.635 ;
        RECT 2168.125 138.125 2168.295 186.235 ;
      LAYER mcon ;
        RECT 2168.585 1641.945 2168.755 1642.115 ;
        RECT 2167.205 1545.385 2167.375 1545.555 ;
        RECT 2168.125 1400.545 2168.295 1400.715 ;
        RECT 2168.125 1303.985 2168.295 1304.155 ;
        RECT 2168.125 883.065 2168.295 883.235 ;
        RECT 2168.125 627.725 2168.295 627.895 ;
        RECT 2167.205 434.605 2167.375 434.775 ;
        RECT 2168.125 289.425 2168.295 289.595 ;
        RECT 2168.125 206.465 2168.295 206.635 ;
        RECT 2168.125 186.065 2168.295 186.235 ;
      LAYER met1 ;
        RECT 2168.510 1666.580 2168.830 1666.640 ;
        RECT 2170.810 1666.580 2171.130 1666.640 ;
        RECT 2168.510 1666.440 2171.130 1666.580 ;
        RECT 2168.510 1666.380 2168.830 1666.440 ;
        RECT 2170.810 1666.380 2171.130 1666.440 ;
        RECT 2168.510 1642.100 2168.830 1642.160 ;
        RECT 2168.315 1641.960 2168.830 1642.100 ;
        RECT 2168.510 1641.900 2168.830 1641.960 ;
        RECT 2168.525 1594.160 2168.815 1594.205 ;
        RECT 2168.970 1594.160 2169.290 1594.220 ;
        RECT 2168.525 1594.020 2169.290 1594.160 ;
        RECT 2168.525 1593.975 2168.815 1594.020 ;
        RECT 2168.970 1593.960 2169.290 1594.020 ;
        RECT 2167.130 1559.480 2167.450 1559.540 ;
        RECT 2168.970 1559.480 2169.290 1559.540 ;
        RECT 2167.130 1559.340 2169.290 1559.480 ;
        RECT 2167.130 1559.280 2167.450 1559.340 ;
        RECT 2168.970 1559.280 2169.290 1559.340 ;
        RECT 2167.130 1545.540 2167.450 1545.600 ;
        RECT 2166.935 1545.400 2167.450 1545.540 ;
        RECT 2167.130 1545.340 2167.450 1545.400 ;
        RECT 2167.145 1497.600 2167.435 1497.645 ;
        RECT 2168.510 1497.600 2168.830 1497.660 ;
        RECT 2167.145 1497.460 2168.830 1497.600 ;
        RECT 2167.145 1497.415 2167.435 1497.460 ;
        RECT 2168.510 1497.400 2168.830 1497.460 ;
        RECT 2168.050 1400.700 2168.370 1400.760 ;
        RECT 2167.855 1400.560 2168.370 1400.700 ;
        RECT 2168.050 1400.500 2168.370 1400.560 ;
        RECT 2168.065 1352.760 2168.355 1352.805 ;
        RECT 2168.510 1352.760 2168.830 1352.820 ;
        RECT 2168.065 1352.620 2168.830 1352.760 ;
        RECT 2168.065 1352.575 2168.355 1352.620 ;
        RECT 2168.510 1352.560 2168.830 1352.620 ;
        RECT 2168.050 1304.140 2168.370 1304.200 ;
        RECT 2167.855 1304.000 2168.370 1304.140 ;
        RECT 2168.050 1303.940 2168.370 1304.000 ;
        RECT 2168.065 1256.200 2168.355 1256.245 ;
        RECT 2168.510 1256.200 2168.830 1256.260 ;
        RECT 2168.065 1256.060 2168.830 1256.200 ;
        RECT 2168.065 1256.015 2168.355 1256.060 ;
        RECT 2168.510 1256.000 2168.830 1256.060 ;
        RECT 2167.130 1159.300 2167.450 1159.360 ;
        RECT 2168.510 1159.300 2168.830 1159.360 ;
        RECT 2167.130 1159.160 2168.830 1159.300 ;
        RECT 2167.130 1159.100 2167.450 1159.160 ;
        RECT 2168.510 1159.100 2168.830 1159.160 ;
        RECT 2167.130 1062.740 2167.450 1062.800 ;
        RECT 2168.510 1062.740 2168.830 1062.800 ;
        RECT 2167.130 1062.600 2168.830 1062.740 ;
        RECT 2167.130 1062.540 2167.450 1062.600 ;
        RECT 2168.510 1062.540 2168.830 1062.600 ;
        RECT 2167.130 966.180 2167.450 966.240 ;
        RECT 2168.510 966.180 2168.830 966.240 ;
        RECT 2167.130 966.040 2168.830 966.180 ;
        RECT 2167.130 965.980 2167.450 966.040 ;
        RECT 2168.510 965.980 2168.830 966.040 ;
        RECT 2168.050 883.220 2168.370 883.280 ;
        RECT 2167.855 883.080 2168.370 883.220 ;
        RECT 2168.050 883.020 2168.370 883.080 ;
        RECT 2168.050 869.620 2168.370 869.680 ;
        RECT 2167.855 869.480 2168.370 869.620 ;
        RECT 2168.050 869.420 2168.370 869.480 ;
        RECT 2166.210 821.000 2166.530 821.060 ;
        RECT 2167.130 821.000 2167.450 821.060 ;
        RECT 2166.210 820.860 2167.450 821.000 ;
        RECT 2166.210 820.800 2166.530 820.860 ;
        RECT 2167.130 820.800 2167.450 820.860 ;
        RECT 2168.050 724.440 2168.370 724.500 ;
        RECT 2168.970 724.440 2169.290 724.500 ;
        RECT 2168.050 724.300 2169.290 724.440 ;
        RECT 2168.050 724.240 2168.370 724.300 ;
        RECT 2168.970 724.240 2169.290 724.300 ;
        RECT 2168.050 627.880 2168.370 627.940 ;
        RECT 2167.855 627.740 2168.370 627.880 ;
        RECT 2168.050 627.680 2168.370 627.740 ;
        RECT 2168.050 593.200 2168.370 593.260 ;
        RECT 2167.855 593.060 2168.370 593.200 ;
        RECT 2168.050 593.000 2168.370 593.060 ;
        RECT 2167.145 434.760 2167.435 434.805 ;
        RECT 2167.590 434.760 2167.910 434.820 ;
        RECT 2167.145 434.620 2167.910 434.760 ;
        RECT 2167.145 434.575 2167.435 434.620 ;
        RECT 2167.590 434.560 2167.910 434.620 ;
        RECT 2167.130 386.480 2167.450 386.540 ;
        RECT 2166.935 386.340 2167.450 386.480 ;
        RECT 2167.130 386.280 2167.450 386.340 ;
        RECT 2167.130 338.200 2167.450 338.260 ;
        RECT 2167.590 338.200 2167.910 338.260 ;
        RECT 2167.130 338.060 2167.910 338.200 ;
        RECT 2167.130 338.000 2167.450 338.060 ;
        RECT 2167.590 338.000 2167.910 338.060 ;
        RECT 2167.590 303.520 2167.910 303.580 ;
        RECT 2168.510 303.520 2168.830 303.580 ;
        RECT 2167.590 303.380 2168.830 303.520 ;
        RECT 2167.590 303.320 2167.910 303.380 ;
        RECT 2168.510 303.320 2168.830 303.380 ;
        RECT 2168.065 289.580 2168.355 289.625 ;
        RECT 2168.510 289.580 2168.830 289.640 ;
        RECT 2168.065 289.440 2168.830 289.580 ;
        RECT 2168.065 289.395 2168.355 289.440 ;
        RECT 2168.510 289.380 2168.830 289.440 ;
        RECT 2168.050 241.640 2168.370 241.700 ;
        RECT 2167.855 241.500 2168.370 241.640 ;
        RECT 2168.050 241.440 2168.370 241.500 ;
        RECT 2168.050 206.620 2168.370 206.680 ;
        RECT 2167.855 206.480 2168.370 206.620 ;
        RECT 2168.050 206.420 2168.370 206.480 ;
        RECT 2167.590 186.900 2167.910 186.960 ;
        RECT 2168.065 186.900 2168.355 186.945 ;
        RECT 2167.590 186.760 2168.355 186.900 ;
        RECT 2167.590 186.700 2167.910 186.760 ;
        RECT 2168.065 186.715 2168.355 186.760 ;
        RECT 2168.050 186.220 2168.370 186.280 ;
        RECT 2167.855 186.080 2168.370 186.220 ;
        RECT 2168.050 186.020 2168.370 186.080 ;
        RECT 2168.065 138.280 2168.355 138.325 ;
        RECT 2168.510 138.280 2168.830 138.340 ;
        RECT 2168.065 138.140 2168.830 138.280 ;
        RECT 2168.065 138.095 2168.355 138.140 ;
        RECT 2168.510 138.080 2168.830 138.140 ;
        RECT 1989.110 27.100 1989.430 27.160 ;
        RECT 2168.050 27.100 2168.370 27.160 ;
        RECT 1989.110 26.960 2168.370 27.100 ;
        RECT 1989.110 26.900 1989.430 26.960 ;
        RECT 2168.050 26.900 2168.370 26.960 ;
      LAYER via ;
        RECT 2168.540 1666.380 2168.800 1666.640 ;
        RECT 2170.840 1666.380 2171.100 1666.640 ;
        RECT 2168.540 1641.900 2168.800 1642.160 ;
        RECT 2169.000 1593.960 2169.260 1594.220 ;
        RECT 2167.160 1559.280 2167.420 1559.540 ;
        RECT 2169.000 1559.280 2169.260 1559.540 ;
        RECT 2167.160 1545.340 2167.420 1545.600 ;
        RECT 2168.540 1497.400 2168.800 1497.660 ;
        RECT 2168.080 1400.500 2168.340 1400.760 ;
        RECT 2168.540 1352.560 2168.800 1352.820 ;
        RECT 2168.080 1303.940 2168.340 1304.200 ;
        RECT 2168.540 1256.000 2168.800 1256.260 ;
        RECT 2167.160 1159.100 2167.420 1159.360 ;
        RECT 2168.540 1159.100 2168.800 1159.360 ;
        RECT 2167.160 1062.540 2167.420 1062.800 ;
        RECT 2168.540 1062.540 2168.800 1062.800 ;
        RECT 2167.160 965.980 2167.420 966.240 ;
        RECT 2168.540 965.980 2168.800 966.240 ;
        RECT 2168.080 883.020 2168.340 883.280 ;
        RECT 2168.080 869.420 2168.340 869.680 ;
        RECT 2166.240 820.800 2166.500 821.060 ;
        RECT 2167.160 820.800 2167.420 821.060 ;
        RECT 2168.080 724.240 2168.340 724.500 ;
        RECT 2169.000 724.240 2169.260 724.500 ;
        RECT 2168.080 627.680 2168.340 627.940 ;
        RECT 2168.080 593.000 2168.340 593.260 ;
        RECT 2167.620 434.560 2167.880 434.820 ;
        RECT 2167.160 386.280 2167.420 386.540 ;
        RECT 2167.160 338.000 2167.420 338.260 ;
        RECT 2167.620 338.000 2167.880 338.260 ;
        RECT 2167.620 303.320 2167.880 303.580 ;
        RECT 2168.540 303.320 2168.800 303.580 ;
        RECT 2168.540 289.380 2168.800 289.640 ;
        RECT 2168.080 241.440 2168.340 241.700 ;
        RECT 2168.080 206.420 2168.340 206.680 ;
        RECT 2167.620 186.700 2167.880 186.960 ;
        RECT 2168.080 186.020 2168.340 186.280 ;
        RECT 2168.540 138.080 2168.800 138.340 ;
        RECT 1989.140 26.900 1989.400 27.160 ;
        RECT 2168.080 26.900 2168.340 27.160 ;
      LAYER met2 ;
        RECT 2172.140 1700.410 2172.420 1702.400 ;
        RECT 2170.900 1700.270 2172.420 1700.410 ;
        RECT 2170.900 1666.670 2171.040 1700.270 ;
        RECT 2172.140 1700.000 2172.420 1700.270 ;
        RECT 2168.540 1666.350 2168.800 1666.670 ;
        RECT 2170.840 1666.350 2171.100 1666.670 ;
        RECT 2168.600 1642.190 2168.740 1666.350 ;
        RECT 2168.540 1641.870 2168.800 1642.190 ;
        RECT 2169.000 1593.930 2169.260 1594.250 ;
        RECT 2169.060 1559.570 2169.200 1593.930 ;
        RECT 2167.160 1559.250 2167.420 1559.570 ;
        RECT 2169.000 1559.250 2169.260 1559.570 ;
        RECT 2167.220 1545.630 2167.360 1559.250 ;
        RECT 2167.160 1545.310 2167.420 1545.630 ;
        RECT 2168.540 1497.370 2168.800 1497.690 ;
        RECT 2168.600 1425.010 2168.740 1497.370 ;
        RECT 2168.140 1424.870 2168.740 1425.010 ;
        RECT 2168.140 1400.790 2168.280 1424.870 ;
        RECT 2168.080 1400.470 2168.340 1400.790 ;
        RECT 2168.540 1352.530 2168.800 1352.850 ;
        RECT 2168.600 1317.570 2168.740 1352.530 ;
        RECT 2168.140 1317.430 2168.740 1317.570 ;
        RECT 2168.140 1304.230 2168.280 1317.430 ;
        RECT 2168.080 1303.910 2168.340 1304.230 ;
        RECT 2168.540 1255.970 2168.800 1256.290 ;
        RECT 2168.600 1221.010 2168.740 1255.970 ;
        RECT 2168.140 1220.870 2168.740 1221.010 ;
        RECT 2168.140 1207.525 2168.280 1220.870 ;
        RECT 2167.150 1207.155 2167.430 1207.525 ;
        RECT 2168.070 1207.155 2168.350 1207.525 ;
        RECT 2167.220 1159.390 2167.360 1207.155 ;
        RECT 2167.160 1159.070 2167.420 1159.390 ;
        RECT 2168.540 1159.070 2168.800 1159.390 ;
        RECT 2168.600 1124.450 2168.740 1159.070 ;
        RECT 2168.140 1124.310 2168.740 1124.450 ;
        RECT 2168.140 1110.965 2168.280 1124.310 ;
        RECT 2167.150 1110.595 2167.430 1110.965 ;
        RECT 2168.070 1110.595 2168.350 1110.965 ;
        RECT 2167.220 1062.830 2167.360 1110.595 ;
        RECT 2167.160 1062.510 2167.420 1062.830 ;
        RECT 2168.540 1062.510 2168.800 1062.830 ;
        RECT 2168.600 1027.890 2168.740 1062.510 ;
        RECT 2168.140 1027.750 2168.740 1027.890 ;
        RECT 2168.140 1014.405 2168.280 1027.750 ;
        RECT 2167.150 1014.035 2167.430 1014.405 ;
        RECT 2168.070 1014.035 2168.350 1014.405 ;
        RECT 2167.220 966.270 2167.360 1014.035 ;
        RECT 2167.160 965.950 2167.420 966.270 ;
        RECT 2168.540 965.950 2168.800 966.270 ;
        RECT 2168.600 931.330 2168.740 965.950 ;
        RECT 2168.140 931.190 2168.740 931.330 ;
        RECT 2168.140 883.310 2168.280 931.190 ;
        RECT 2168.080 882.990 2168.340 883.310 ;
        RECT 2168.080 869.390 2168.340 869.710 ;
        RECT 2168.140 834.770 2168.280 869.390 ;
        RECT 2167.220 834.630 2168.280 834.770 ;
        RECT 2167.220 821.090 2167.360 834.630 ;
        RECT 2166.240 820.770 2166.500 821.090 ;
        RECT 2167.160 820.770 2167.420 821.090 ;
        RECT 2166.300 773.005 2166.440 820.770 ;
        RECT 2166.230 772.635 2166.510 773.005 ;
        RECT 2168.530 772.635 2168.810 773.005 ;
        RECT 2168.600 738.210 2168.740 772.635 ;
        RECT 2168.140 738.070 2168.740 738.210 ;
        RECT 2168.140 724.530 2168.280 738.070 ;
        RECT 2168.080 724.210 2168.340 724.530 ;
        RECT 2169.000 724.210 2169.260 724.530 ;
        RECT 2169.060 676.445 2169.200 724.210 ;
        RECT 2168.070 676.075 2168.350 676.445 ;
        RECT 2168.990 676.075 2169.270 676.445 ;
        RECT 2168.140 627.970 2168.280 676.075 ;
        RECT 2168.080 627.650 2168.340 627.970 ;
        RECT 2168.080 592.970 2168.340 593.290 ;
        RECT 2168.140 579.770 2168.280 592.970 ;
        RECT 2168.140 579.630 2168.740 579.770 ;
        RECT 2168.600 545.090 2168.740 579.630 ;
        RECT 2168.140 544.950 2168.740 545.090 ;
        RECT 2168.140 507.010 2168.280 544.950 ;
        RECT 2167.220 506.870 2168.280 507.010 ;
        RECT 2167.220 483.325 2167.360 506.870 ;
        RECT 2167.150 482.955 2167.430 483.325 ;
        RECT 2168.530 482.955 2168.810 483.325 ;
        RECT 2168.600 448.530 2168.740 482.955 ;
        RECT 2167.680 448.390 2168.740 448.530 ;
        RECT 2167.680 434.850 2167.820 448.390 ;
        RECT 2167.620 434.530 2167.880 434.850 ;
        RECT 2167.160 386.250 2167.420 386.570 ;
        RECT 2167.220 338.290 2167.360 386.250 ;
        RECT 2167.160 337.970 2167.420 338.290 ;
        RECT 2167.620 337.970 2167.880 338.290 ;
        RECT 2167.680 303.610 2167.820 337.970 ;
        RECT 2167.620 303.290 2167.880 303.610 ;
        RECT 2168.540 303.290 2168.800 303.610 ;
        RECT 2168.600 289.670 2168.740 303.290 ;
        RECT 2168.540 289.350 2168.800 289.670 ;
        RECT 2168.080 241.410 2168.340 241.730 ;
        RECT 2168.140 206.710 2168.280 241.410 ;
        RECT 2168.080 206.390 2168.340 206.710 ;
        RECT 2167.620 186.730 2167.880 186.990 ;
        RECT 2167.620 186.670 2168.280 186.730 ;
        RECT 2167.680 186.590 2168.280 186.670 ;
        RECT 2168.140 186.310 2168.280 186.590 ;
        RECT 2168.080 185.990 2168.340 186.310 ;
        RECT 2168.540 138.050 2168.800 138.370 ;
        RECT 2168.600 113.970 2168.740 138.050 ;
        RECT 2168.140 113.830 2168.740 113.970 ;
        RECT 2168.140 27.190 2168.280 113.830 ;
        RECT 1989.140 26.870 1989.400 27.190 ;
        RECT 2168.080 26.870 2168.340 27.190 ;
        RECT 1989.200 2.400 1989.340 26.870 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
      LAYER via2 ;
        RECT 2167.150 1207.200 2167.430 1207.480 ;
        RECT 2168.070 1207.200 2168.350 1207.480 ;
        RECT 2167.150 1110.640 2167.430 1110.920 ;
        RECT 2168.070 1110.640 2168.350 1110.920 ;
        RECT 2167.150 1014.080 2167.430 1014.360 ;
        RECT 2168.070 1014.080 2168.350 1014.360 ;
        RECT 2166.230 772.680 2166.510 772.960 ;
        RECT 2168.530 772.680 2168.810 772.960 ;
        RECT 2168.070 676.120 2168.350 676.400 ;
        RECT 2168.990 676.120 2169.270 676.400 ;
        RECT 2167.150 483.000 2167.430 483.280 ;
        RECT 2168.530 483.000 2168.810 483.280 ;
      LAYER met3 ;
        RECT 2167.125 1207.490 2167.455 1207.505 ;
        RECT 2168.045 1207.490 2168.375 1207.505 ;
        RECT 2167.125 1207.190 2168.375 1207.490 ;
        RECT 2167.125 1207.175 2167.455 1207.190 ;
        RECT 2168.045 1207.175 2168.375 1207.190 ;
        RECT 2167.125 1110.930 2167.455 1110.945 ;
        RECT 2168.045 1110.930 2168.375 1110.945 ;
        RECT 2167.125 1110.630 2168.375 1110.930 ;
        RECT 2167.125 1110.615 2167.455 1110.630 ;
        RECT 2168.045 1110.615 2168.375 1110.630 ;
        RECT 2167.125 1014.370 2167.455 1014.385 ;
        RECT 2168.045 1014.370 2168.375 1014.385 ;
        RECT 2167.125 1014.070 2168.375 1014.370 ;
        RECT 2167.125 1014.055 2167.455 1014.070 ;
        RECT 2168.045 1014.055 2168.375 1014.070 ;
        RECT 2166.205 772.970 2166.535 772.985 ;
        RECT 2168.505 772.970 2168.835 772.985 ;
        RECT 2166.205 772.670 2168.835 772.970 ;
        RECT 2166.205 772.655 2166.535 772.670 ;
        RECT 2168.505 772.655 2168.835 772.670 ;
        RECT 2168.045 676.410 2168.375 676.425 ;
        RECT 2168.965 676.410 2169.295 676.425 ;
        RECT 2168.045 676.110 2169.295 676.410 ;
        RECT 2168.045 676.095 2168.375 676.110 ;
        RECT 2168.965 676.095 2169.295 676.110 ;
        RECT 2167.125 483.290 2167.455 483.305 ;
        RECT 2168.505 483.290 2168.835 483.305 ;
        RECT 2167.125 482.990 2168.835 483.290 ;
        RECT 2167.125 482.975 2167.455 482.990 ;
        RECT 2168.505 482.975 2168.835 482.990 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2006.590 27.440 2006.910 27.500 ;
        RECT 2180.930 27.440 2181.250 27.500 ;
        RECT 2006.590 27.300 2181.250 27.440 ;
        RECT 2006.590 27.240 2006.910 27.300 ;
        RECT 2180.930 27.240 2181.250 27.300 ;
      LAYER via ;
        RECT 2006.620 27.240 2006.880 27.500 ;
        RECT 2180.960 27.240 2181.220 27.500 ;
      LAYER met2 ;
        RECT 2181.340 1700.410 2181.620 1702.400 ;
        RECT 2181.020 1700.270 2181.620 1700.410 ;
        RECT 2181.020 27.530 2181.160 1700.270 ;
        RECT 2181.340 1700.000 2181.620 1700.270 ;
        RECT 2006.620 27.210 2006.880 27.530 ;
        RECT 2180.960 27.210 2181.220 27.530 ;
        RECT 2006.680 2.400 2006.820 27.210 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2024.530 23.700 2024.850 23.760 ;
        RECT 2188.750 23.700 2189.070 23.760 ;
        RECT 2024.530 23.560 2189.070 23.700 ;
        RECT 2024.530 23.500 2024.850 23.560 ;
        RECT 2188.750 23.500 2189.070 23.560 ;
      LAYER via ;
        RECT 2024.560 23.500 2024.820 23.760 ;
        RECT 2188.780 23.500 2189.040 23.760 ;
      LAYER met2 ;
        RECT 2190.540 1700.410 2190.820 1702.400 ;
        RECT 2188.840 1700.270 2190.820 1700.410 ;
        RECT 2188.840 23.790 2188.980 1700.270 ;
        RECT 2190.540 1700.000 2190.820 1700.270 ;
        RECT 2024.560 23.470 2024.820 23.790 ;
        RECT 2188.780 23.470 2189.040 23.790 ;
        RECT 2024.620 2.400 2024.760 23.470 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2048.910 1689.020 2049.230 1689.080 ;
        RECT 2199.790 1689.020 2200.110 1689.080 ;
        RECT 2048.910 1688.880 2200.110 1689.020 ;
        RECT 2048.910 1688.820 2049.230 1688.880 ;
        RECT 2199.790 1688.820 2200.110 1688.880 ;
        RECT 2042.470 17.240 2042.790 17.300 ;
        RECT 2048.910 17.240 2049.230 17.300 ;
        RECT 2042.470 17.100 2049.230 17.240 ;
        RECT 2042.470 17.040 2042.790 17.100 ;
        RECT 2048.910 17.040 2049.230 17.100 ;
      LAYER via ;
        RECT 2048.940 1688.820 2049.200 1689.080 ;
        RECT 2199.820 1688.820 2200.080 1689.080 ;
        RECT 2042.500 17.040 2042.760 17.300 ;
        RECT 2048.940 17.040 2049.200 17.300 ;
      LAYER met2 ;
        RECT 2199.740 1700.000 2200.020 1702.400 ;
        RECT 2199.880 1689.110 2200.020 1700.000 ;
        RECT 2048.940 1688.790 2049.200 1689.110 ;
        RECT 2199.820 1688.790 2200.080 1689.110 ;
        RECT 2049.000 17.330 2049.140 1688.790 ;
        RECT 2042.500 17.010 2042.760 17.330 ;
        RECT 2048.940 17.010 2049.200 17.330 ;
        RECT 2042.560 2.400 2042.700 17.010 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.610 66.880 758.930 66.940 ;
        RECT 1539.690 66.880 1540.010 66.940 ;
        RECT 758.610 66.740 1540.010 66.880 ;
        RECT 758.610 66.680 758.930 66.740 ;
        RECT 1539.690 66.680 1540.010 66.740 ;
      LAYER via ;
        RECT 758.640 66.680 758.900 66.940 ;
        RECT 1539.720 66.680 1539.980 66.940 ;
      LAYER met2 ;
        RECT 1538.720 1700.410 1539.000 1702.400 ;
        RECT 1538.720 1700.270 1539.920 1700.410 ;
        RECT 1538.720 1700.000 1539.000 1700.270 ;
        RECT 1539.780 66.970 1539.920 1700.270 ;
        RECT 758.640 66.650 758.900 66.970 ;
        RECT 1539.720 66.650 1539.980 66.970 ;
        RECT 758.700 17.410 758.840 66.650 ;
        RECT 757.780 17.270 758.840 17.410 ;
        RECT 757.780 2.400 757.920 17.270 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2062.710 1688.680 2063.030 1688.740 ;
        RECT 2208.990 1688.680 2209.310 1688.740 ;
        RECT 2062.710 1688.540 2209.310 1688.680 ;
        RECT 2062.710 1688.480 2063.030 1688.540 ;
        RECT 2208.990 1688.480 2209.310 1688.540 ;
        RECT 2060.410 20.640 2060.730 20.700 ;
        RECT 2062.710 20.640 2063.030 20.700 ;
        RECT 2060.410 20.500 2063.030 20.640 ;
        RECT 2060.410 20.440 2060.730 20.500 ;
        RECT 2062.710 20.440 2063.030 20.500 ;
      LAYER via ;
        RECT 2062.740 1688.480 2063.000 1688.740 ;
        RECT 2209.020 1688.480 2209.280 1688.740 ;
        RECT 2060.440 20.440 2060.700 20.700 ;
        RECT 2062.740 20.440 2063.000 20.700 ;
      LAYER met2 ;
        RECT 2208.940 1700.000 2209.220 1702.400 ;
        RECT 2209.080 1688.770 2209.220 1700.000 ;
        RECT 2062.740 1688.450 2063.000 1688.770 ;
        RECT 2209.020 1688.450 2209.280 1688.770 ;
        RECT 2062.800 20.730 2062.940 1688.450 ;
        RECT 2060.440 20.410 2060.700 20.730 ;
        RECT 2062.740 20.410 2063.000 20.730 ;
        RECT 2060.500 2.400 2060.640 20.410 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2083.410 1690.040 2083.730 1690.100 ;
        RECT 2218.190 1690.040 2218.510 1690.100 ;
        RECT 2083.410 1689.900 2218.510 1690.040 ;
        RECT 2083.410 1689.840 2083.730 1689.900 ;
        RECT 2218.190 1689.840 2218.510 1689.900 ;
        RECT 2078.350 15.540 2078.670 15.600 ;
        RECT 2083.410 15.540 2083.730 15.600 ;
        RECT 2078.350 15.400 2083.730 15.540 ;
        RECT 2078.350 15.340 2078.670 15.400 ;
        RECT 2083.410 15.340 2083.730 15.400 ;
      LAYER via ;
        RECT 2083.440 1689.840 2083.700 1690.100 ;
        RECT 2218.220 1689.840 2218.480 1690.100 ;
        RECT 2078.380 15.340 2078.640 15.600 ;
        RECT 2083.440 15.340 2083.700 15.600 ;
      LAYER met2 ;
        RECT 2218.140 1700.000 2218.420 1702.400 ;
        RECT 2218.280 1690.130 2218.420 1700.000 ;
        RECT 2083.440 1689.810 2083.700 1690.130 ;
        RECT 2218.220 1689.810 2218.480 1690.130 ;
        RECT 2083.500 15.630 2083.640 1689.810 ;
        RECT 2078.380 15.310 2078.640 15.630 ;
        RECT 2083.440 15.310 2083.700 15.630 ;
        RECT 2078.440 2.400 2078.580 15.310 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2137.765 1684.105 2137.935 1690.395 ;
      LAYER mcon ;
        RECT 2137.765 1690.225 2137.935 1690.395 ;
      LAYER met1 ;
        RECT 2137.705 1690.380 2137.995 1690.425 ;
        RECT 2227.390 1690.380 2227.710 1690.440 ;
        RECT 2137.705 1690.240 2227.710 1690.380 ;
        RECT 2137.705 1690.195 2137.995 1690.240 ;
        RECT 2227.390 1690.180 2227.710 1690.240 ;
        RECT 2100.890 1684.940 2101.210 1685.000 ;
        RECT 2100.890 1684.800 2110.320 1684.940 ;
        RECT 2100.890 1684.740 2101.210 1684.800 ;
        RECT 2110.180 1684.600 2110.320 1684.800 ;
        RECT 2110.180 1684.460 2124.120 1684.600 ;
        RECT 2123.980 1684.260 2124.120 1684.460 ;
        RECT 2137.705 1684.260 2137.995 1684.305 ;
        RECT 2123.980 1684.120 2137.995 1684.260 ;
        RECT 2137.705 1684.075 2137.995 1684.120 ;
        RECT 2095.830 20.640 2096.150 20.700 ;
        RECT 2100.890 20.640 2101.210 20.700 ;
        RECT 2095.830 20.500 2101.210 20.640 ;
        RECT 2095.830 20.440 2096.150 20.500 ;
        RECT 2100.890 20.440 2101.210 20.500 ;
      LAYER via ;
        RECT 2227.420 1690.180 2227.680 1690.440 ;
        RECT 2100.920 1684.740 2101.180 1685.000 ;
        RECT 2095.860 20.440 2096.120 20.700 ;
        RECT 2100.920 20.440 2101.180 20.700 ;
      LAYER met2 ;
        RECT 2227.340 1700.000 2227.620 1702.400 ;
        RECT 2227.480 1690.470 2227.620 1700.000 ;
        RECT 2227.420 1690.150 2227.680 1690.470 ;
        RECT 2100.920 1684.710 2101.180 1685.030 ;
        RECT 2100.980 20.730 2101.120 1684.710 ;
        RECT 2095.860 20.410 2096.120 20.730 ;
        RECT 2100.920 20.410 2101.180 20.730 ;
        RECT 2095.920 2.400 2096.060 20.410 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2163.065 1685.465 2163.235 1686.995 ;
      LAYER mcon ;
        RECT 2163.065 1686.825 2163.235 1686.995 ;
      LAYER met1 ;
        RECT 2163.005 1686.980 2163.295 1687.025 ;
        RECT 2236.590 1686.980 2236.910 1687.040 ;
        RECT 2163.005 1686.840 2236.910 1686.980 ;
        RECT 2163.005 1686.795 2163.295 1686.840 ;
        RECT 2236.590 1686.780 2236.910 1686.840 ;
        RECT 2117.910 1685.620 2118.230 1685.680 ;
        RECT 2163.005 1685.620 2163.295 1685.665 ;
        RECT 2117.910 1685.480 2163.295 1685.620 ;
        RECT 2117.910 1685.420 2118.230 1685.480 ;
        RECT 2163.005 1685.435 2163.295 1685.480 ;
        RECT 2113.770 20.640 2114.090 20.700 ;
        RECT 2117.910 20.640 2118.230 20.700 ;
        RECT 2113.770 20.500 2118.230 20.640 ;
        RECT 2113.770 20.440 2114.090 20.500 ;
        RECT 2117.910 20.440 2118.230 20.500 ;
      LAYER via ;
        RECT 2236.620 1686.780 2236.880 1687.040 ;
        RECT 2117.940 1685.420 2118.200 1685.680 ;
        RECT 2113.800 20.440 2114.060 20.700 ;
        RECT 2117.940 20.440 2118.200 20.700 ;
      LAYER met2 ;
        RECT 2236.540 1700.000 2236.820 1702.400 ;
        RECT 2236.680 1687.070 2236.820 1700.000 ;
        RECT 2236.620 1686.750 2236.880 1687.070 ;
        RECT 2117.940 1685.390 2118.200 1685.710 ;
        RECT 2118.000 20.730 2118.140 1685.390 ;
        RECT 2113.800 20.410 2114.060 20.730 ;
        RECT 2117.940 20.410 2118.200 20.730 ;
        RECT 2113.860 2.400 2114.000 20.410 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2166.745 1685.805 2166.915 1686.655 ;
      LAYER mcon ;
        RECT 2166.745 1686.485 2166.915 1686.655 ;
      LAYER met1 ;
        RECT 2142.750 1686.640 2143.070 1686.700 ;
        RECT 2166.685 1686.640 2166.975 1686.685 ;
        RECT 2142.750 1686.500 2166.975 1686.640 ;
        RECT 2142.750 1686.440 2143.070 1686.500 ;
        RECT 2166.685 1686.455 2166.975 1686.500 ;
        RECT 2166.685 1685.960 2166.975 1686.005 ;
        RECT 2245.790 1685.960 2246.110 1686.020 ;
        RECT 2166.685 1685.820 2246.110 1685.960 ;
        RECT 2166.685 1685.775 2166.975 1685.820 ;
        RECT 2245.790 1685.760 2246.110 1685.820 ;
        RECT 2131.710 17.580 2132.030 17.640 ;
        RECT 2142.290 17.580 2142.610 17.640 ;
        RECT 2131.710 17.440 2142.610 17.580 ;
        RECT 2131.710 17.380 2132.030 17.440 ;
        RECT 2142.290 17.380 2142.610 17.440 ;
      LAYER via ;
        RECT 2142.780 1686.440 2143.040 1686.700 ;
        RECT 2245.820 1685.760 2246.080 1686.020 ;
        RECT 2131.740 17.380 2132.000 17.640 ;
        RECT 2142.320 17.380 2142.580 17.640 ;
      LAYER met2 ;
        RECT 2245.740 1700.000 2246.020 1702.400 ;
        RECT 2142.780 1686.410 2143.040 1686.730 ;
        RECT 2142.840 1656.210 2142.980 1686.410 ;
        RECT 2245.880 1686.050 2246.020 1700.000 ;
        RECT 2245.820 1685.730 2246.080 1686.050 ;
        RECT 2142.380 1656.070 2142.980 1656.210 ;
        RECT 2142.380 17.670 2142.520 1656.070 ;
        RECT 2131.740 17.350 2132.000 17.670 ;
        RECT 2142.320 17.350 2142.580 17.670 ;
        RECT 2131.800 2.400 2131.940 17.350 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2160.765 1686.825 2160.935 1688.015 ;
        RECT 2220.105 1687.505 2220.275 1689.375 ;
      LAYER mcon ;
        RECT 2220.105 1689.205 2220.275 1689.375 ;
        RECT 2160.765 1687.845 2160.935 1688.015 ;
      LAYER met1 ;
        RECT 2220.045 1689.360 2220.335 1689.405 ;
        RECT 2254.990 1689.360 2255.310 1689.420 ;
        RECT 2220.045 1689.220 2255.310 1689.360 ;
        RECT 2220.045 1689.175 2220.335 1689.220 ;
        RECT 2254.990 1689.160 2255.310 1689.220 ;
        RECT 2160.705 1688.000 2160.995 1688.045 ;
        RECT 2160.705 1687.860 2167.820 1688.000 ;
        RECT 2160.705 1687.815 2160.995 1687.860 ;
        RECT 2167.680 1687.660 2167.820 1687.860 ;
        RECT 2220.045 1687.660 2220.335 1687.705 ;
        RECT 2167.680 1687.520 2220.335 1687.660 ;
        RECT 2220.045 1687.475 2220.335 1687.520 ;
        RECT 2152.410 1686.980 2152.730 1687.040 ;
        RECT 2160.705 1686.980 2160.995 1687.025 ;
        RECT 2152.410 1686.840 2160.995 1686.980 ;
        RECT 2152.410 1686.780 2152.730 1686.840 ;
        RECT 2160.705 1686.795 2160.995 1686.840 ;
        RECT 2149.650 20.640 2149.970 20.700 ;
        RECT 2152.410 20.640 2152.730 20.700 ;
        RECT 2149.650 20.500 2152.730 20.640 ;
        RECT 2149.650 20.440 2149.970 20.500 ;
        RECT 2152.410 20.440 2152.730 20.500 ;
      LAYER via ;
        RECT 2255.020 1689.160 2255.280 1689.420 ;
        RECT 2152.440 1686.780 2152.700 1687.040 ;
        RECT 2149.680 20.440 2149.940 20.700 ;
        RECT 2152.440 20.440 2152.700 20.700 ;
      LAYER met2 ;
        RECT 2254.940 1700.000 2255.220 1702.400 ;
        RECT 2255.080 1689.450 2255.220 1700.000 ;
        RECT 2255.020 1689.130 2255.280 1689.450 ;
        RECT 2152.440 1686.750 2152.700 1687.070 ;
        RECT 2152.500 20.730 2152.640 1686.750 ;
        RECT 2149.680 20.410 2149.940 20.730 ;
        RECT 2152.440 20.410 2152.700 20.730 ;
        RECT 2149.740 2.400 2149.880 20.410 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2173.110 1688.000 2173.430 1688.060 ;
        RECT 2264.190 1688.000 2264.510 1688.060 ;
        RECT 2173.110 1687.860 2264.510 1688.000 ;
        RECT 2173.110 1687.800 2173.430 1687.860 ;
        RECT 2264.190 1687.800 2264.510 1687.860 ;
        RECT 2167.590 20.640 2167.910 20.700 ;
        RECT 2173.110 20.640 2173.430 20.700 ;
        RECT 2167.590 20.500 2173.430 20.640 ;
        RECT 2167.590 20.440 2167.910 20.500 ;
        RECT 2173.110 20.440 2173.430 20.500 ;
      LAYER via ;
        RECT 2173.140 1687.800 2173.400 1688.060 ;
        RECT 2264.220 1687.800 2264.480 1688.060 ;
        RECT 2167.620 20.440 2167.880 20.700 ;
        RECT 2173.140 20.440 2173.400 20.700 ;
      LAYER met2 ;
        RECT 2264.140 1700.000 2264.420 1702.400 ;
        RECT 2264.280 1688.090 2264.420 1700.000 ;
        RECT 2173.140 1687.770 2173.400 1688.090 ;
        RECT 2264.220 1687.770 2264.480 1688.090 ;
        RECT 2173.200 20.730 2173.340 1687.770 ;
        RECT 2167.620 20.410 2167.880 20.730 ;
        RECT 2173.140 20.410 2173.400 20.730 ;
        RECT 2167.680 2.400 2167.820 20.410 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2211.750 1688.680 2212.070 1688.740 ;
        RECT 2273.390 1688.680 2273.710 1688.740 ;
        RECT 2211.750 1688.540 2273.710 1688.680 ;
        RECT 2211.750 1688.480 2212.070 1688.540 ;
        RECT 2273.390 1688.480 2273.710 1688.540 ;
        RECT 2185.070 20.640 2185.390 20.700 ;
        RECT 2211.750 20.640 2212.070 20.700 ;
        RECT 2185.070 20.500 2212.070 20.640 ;
        RECT 2185.070 20.440 2185.390 20.500 ;
        RECT 2211.750 20.440 2212.070 20.500 ;
      LAYER via ;
        RECT 2211.780 1688.480 2212.040 1688.740 ;
        RECT 2273.420 1688.480 2273.680 1688.740 ;
        RECT 2185.100 20.440 2185.360 20.700 ;
        RECT 2211.780 20.440 2212.040 20.700 ;
      LAYER met2 ;
        RECT 2273.340 1700.000 2273.620 1702.400 ;
        RECT 2273.480 1688.770 2273.620 1700.000 ;
        RECT 2211.780 1688.450 2212.040 1688.770 ;
        RECT 2273.420 1688.450 2273.680 1688.770 ;
        RECT 2211.840 20.730 2211.980 1688.450 ;
        RECT 2185.100 20.410 2185.360 20.730 ;
        RECT 2211.780 20.410 2212.040 20.730 ;
        RECT 2185.160 2.400 2185.300 20.410 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2225.090 1689.020 2225.410 1689.080 ;
        RECT 2282.590 1689.020 2282.910 1689.080 ;
        RECT 2225.090 1688.880 2282.910 1689.020 ;
        RECT 2225.090 1688.820 2225.410 1688.880 ;
        RECT 2282.590 1688.820 2282.910 1688.880 ;
        RECT 2203.010 20.300 2203.330 20.360 ;
        RECT 2225.090 20.300 2225.410 20.360 ;
        RECT 2203.010 20.160 2225.410 20.300 ;
        RECT 2203.010 20.100 2203.330 20.160 ;
        RECT 2225.090 20.100 2225.410 20.160 ;
      LAYER via ;
        RECT 2225.120 1688.820 2225.380 1689.080 ;
        RECT 2282.620 1688.820 2282.880 1689.080 ;
        RECT 2203.040 20.100 2203.300 20.360 ;
        RECT 2225.120 20.100 2225.380 20.360 ;
      LAYER met2 ;
        RECT 2282.540 1700.000 2282.820 1702.400 ;
        RECT 2282.680 1689.110 2282.820 1700.000 ;
        RECT 2225.120 1688.790 2225.380 1689.110 ;
        RECT 2282.620 1688.790 2282.880 1689.110 ;
        RECT 2225.180 20.390 2225.320 1688.790 ;
        RECT 2203.040 20.070 2203.300 20.390 ;
        RECT 2225.120 20.070 2225.380 20.390 ;
        RECT 2203.100 2.400 2203.240 20.070 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2231.990 1687.320 2232.310 1687.380 ;
        RECT 2291.790 1687.320 2292.110 1687.380 ;
        RECT 2231.990 1687.180 2292.110 1687.320 ;
        RECT 2231.990 1687.120 2232.310 1687.180 ;
        RECT 2291.790 1687.120 2292.110 1687.180 ;
        RECT 2220.950 17.240 2221.270 17.300 ;
        RECT 2231.990 17.240 2232.310 17.300 ;
        RECT 2220.950 17.100 2232.310 17.240 ;
        RECT 2220.950 17.040 2221.270 17.100 ;
        RECT 2231.990 17.040 2232.310 17.100 ;
      LAYER via ;
        RECT 2232.020 1687.120 2232.280 1687.380 ;
        RECT 2291.820 1687.120 2292.080 1687.380 ;
        RECT 2220.980 17.040 2221.240 17.300 ;
        RECT 2232.020 17.040 2232.280 17.300 ;
      LAYER met2 ;
        RECT 2291.740 1700.000 2292.020 1702.400 ;
        RECT 2291.880 1687.410 2292.020 1700.000 ;
        RECT 2232.020 1687.090 2232.280 1687.410 ;
        RECT 2291.820 1687.090 2292.080 1687.410 ;
        RECT 2232.080 17.330 2232.220 1687.090 ;
        RECT 2220.980 17.010 2221.240 17.330 ;
        RECT 2232.020 17.010 2232.280 17.330 ;
        RECT 2221.040 2.400 2221.180 17.010 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.310 68.240 779.630 68.300 ;
        RECT 1545.670 68.240 1545.990 68.300 ;
        RECT 779.310 68.100 1545.990 68.240 ;
        RECT 779.310 68.040 779.630 68.100 ;
        RECT 1545.670 68.040 1545.990 68.100 ;
      LAYER via ;
        RECT 779.340 68.040 779.600 68.300 ;
        RECT 1545.700 68.040 1545.960 68.300 ;
      LAYER met2 ;
        RECT 1547.920 1700.410 1548.200 1702.400 ;
        RECT 1545.760 1700.270 1548.200 1700.410 ;
        RECT 1545.760 68.330 1545.900 1700.270 ;
        RECT 1547.920 1700.000 1548.200 1700.270 ;
        RECT 779.340 68.010 779.600 68.330 ;
        RECT 1545.700 68.010 1545.960 68.330 ;
        RECT 779.400 16.730 779.540 68.010 ;
        RECT 775.720 16.590 779.540 16.730 ;
        RECT 775.720 2.400 775.860 16.590 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2242.110 1686.980 2242.430 1687.040 ;
        RECT 2300.990 1686.980 2301.310 1687.040 ;
        RECT 2242.110 1686.840 2301.310 1686.980 ;
        RECT 2242.110 1686.780 2242.430 1686.840 ;
        RECT 2300.990 1686.780 2301.310 1686.840 ;
        RECT 2238.890 17.920 2239.210 17.980 ;
        RECT 2242.110 17.920 2242.430 17.980 ;
        RECT 2238.890 17.780 2242.430 17.920 ;
        RECT 2238.890 17.720 2239.210 17.780 ;
        RECT 2242.110 17.720 2242.430 17.780 ;
      LAYER via ;
        RECT 2242.140 1686.780 2242.400 1687.040 ;
        RECT 2301.020 1686.780 2301.280 1687.040 ;
        RECT 2238.920 17.720 2239.180 17.980 ;
        RECT 2242.140 17.720 2242.400 17.980 ;
      LAYER met2 ;
        RECT 2300.940 1700.000 2301.220 1702.400 ;
        RECT 2301.080 1687.070 2301.220 1700.000 ;
        RECT 2242.140 1686.750 2242.400 1687.070 ;
        RECT 2301.020 1686.750 2301.280 1687.070 ;
        RECT 2242.200 18.010 2242.340 1686.750 ;
        RECT 2238.920 17.690 2239.180 18.010 ;
        RECT 2242.140 17.690 2242.400 18.010 ;
        RECT 2238.980 2.400 2239.120 17.690 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2266.490 1689.360 2266.810 1689.420 ;
        RECT 2310.190 1689.360 2310.510 1689.420 ;
        RECT 2266.490 1689.220 2310.510 1689.360 ;
        RECT 2266.490 1689.160 2266.810 1689.220 ;
        RECT 2310.190 1689.160 2310.510 1689.220 ;
        RECT 2256.370 20.640 2256.690 20.700 ;
        RECT 2266.490 20.640 2266.810 20.700 ;
        RECT 2256.370 20.500 2266.810 20.640 ;
        RECT 2256.370 20.440 2256.690 20.500 ;
        RECT 2266.490 20.440 2266.810 20.500 ;
      LAYER via ;
        RECT 2266.520 1689.160 2266.780 1689.420 ;
        RECT 2310.220 1689.160 2310.480 1689.420 ;
        RECT 2256.400 20.440 2256.660 20.700 ;
        RECT 2266.520 20.440 2266.780 20.700 ;
      LAYER met2 ;
        RECT 2310.140 1700.000 2310.420 1702.400 ;
        RECT 2310.280 1689.450 2310.420 1700.000 ;
        RECT 2266.520 1689.130 2266.780 1689.450 ;
        RECT 2310.220 1689.130 2310.480 1689.450 ;
        RECT 2266.580 20.730 2266.720 1689.130 ;
        RECT 2256.400 20.410 2256.660 20.730 ;
        RECT 2266.520 20.410 2266.780 20.730 ;
        RECT 2256.460 2.400 2256.600 20.410 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2280.290 1688.680 2280.610 1688.740 ;
        RECT 2319.390 1688.680 2319.710 1688.740 ;
        RECT 2280.290 1688.540 2319.710 1688.680 ;
        RECT 2280.290 1688.480 2280.610 1688.540 ;
        RECT 2319.390 1688.480 2319.710 1688.540 ;
        RECT 2274.310 20.640 2274.630 20.700 ;
        RECT 2280.290 20.640 2280.610 20.700 ;
        RECT 2274.310 20.500 2280.610 20.640 ;
        RECT 2274.310 20.440 2274.630 20.500 ;
        RECT 2280.290 20.440 2280.610 20.500 ;
      LAYER via ;
        RECT 2280.320 1688.480 2280.580 1688.740 ;
        RECT 2319.420 1688.480 2319.680 1688.740 ;
        RECT 2274.340 20.440 2274.600 20.700 ;
        RECT 2280.320 20.440 2280.580 20.700 ;
      LAYER met2 ;
        RECT 2319.340 1700.000 2319.620 1702.400 ;
        RECT 2319.480 1688.770 2319.620 1700.000 ;
        RECT 2280.320 1688.450 2280.580 1688.770 ;
        RECT 2319.420 1688.450 2319.680 1688.770 ;
        RECT 2280.380 20.730 2280.520 1688.450 ;
        RECT 2274.340 20.410 2274.600 20.730 ;
        RECT 2280.320 20.410 2280.580 20.730 ;
        RECT 2274.400 2.400 2274.540 20.410 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2322.150 1683.920 2322.470 1683.980 ;
        RECT 2328.590 1683.920 2328.910 1683.980 ;
        RECT 2322.150 1683.780 2328.910 1683.920 ;
        RECT 2322.150 1683.720 2322.470 1683.780 ;
        RECT 2328.590 1683.720 2328.910 1683.780 ;
        RECT 2292.250 19.960 2292.570 20.020 ;
        RECT 2322.150 19.960 2322.470 20.020 ;
        RECT 2292.250 19.820 2322.470 19.960 ;
        RECT 2292.250 19.760 2292.570 19.820 ;
        RECT 2322.150 19.760 2322.470 19.820 ;
      LAYER via ;
        RECT 2322.180 1683.720 2322.440 1683.980 ;
        RECT 2328.620 1683.720 2328.880 1683.980 ;
        RECT 2292.280 19.760 2292.540 20.020 ;
        RECT 2322.180 19.760 2322.440 20.020 ;
      LAYER met2 ;
        RECT 2328.540 1700.000 2328.820 1702.400 ;
        RECT 2328.680 1684.010 2328.820 1700.000 ;
        RECT 2322.180 1683.690 2322.440 1684.010 ;
        RECT 2328.620 1683.690 2328.880 1684.010 ;
        RECT 2322.240 20.050 2322.380 1683.690 ;
        RECT 2292.280 19.730 2292.540 20.050 ;
        RECT 2322.180 19.730 2322.440 20.050 ;
        RECT 2292.340 2.400 2292.480 19.730 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2332.805 1594.005 2332.975 1608.115 ;
        RECT 2332.805 1497.445 2332.975 1545.555 ;
        RECT 2332.805 1352.605 2332.975 1400.715 ;
        RECT 2332.805 1256.045 2332.975 1304.155 ;
        RECT 2332.805 737.885 2332.975 772.395 ;
        RECT 2333.265 572.645 2333.435 620.755 ;
        RECT 2332.805 379.525 2332.975 427.635 ;
        RECT 2332.345 282.965 2332.515 331.075 ;
      LAYER mcon ;
        RECT 2332.805 1607.945 2332.975 1608.115 ;
        RECT 2332.805 1545.385 2332.975 1545.555 ;
        RECT 2332.805 1400.545 2332.975 1400.715 ;
        RECT 2332.805 1303.985 2332.975 1304.155 ;
        RECT 2332.805 772.225 2332.975 772.395 ;
        RECT 2333.265 620.585 2333.435 620.755 ;
        RECT 2332.805 427.465 2332.975 427.635 ;
        RECT 2332.345 330.905 2332.515 331.075 ;
      LAYER met1 ;
        RECT 2332.730 1666.580 2333.050 1666.640 ;
        RECT 2335.490 1666.580 2335.810 1666.640 ;
        RECT 2332.730 1666.440 2335.810 1666.580 ;
        RECT 2332.730 1666.380 2333.050 1666.440 ;
        RECT 2335.490 1666.380 2335.810 1666.440 ;
        RECT 2332.730 1608.100 2333.050 1608.160 ;
        RECT 2332.535 1607.960 2333.050 1608.100 ;
        RECT 2332.730 1607.900 2333.050 1607.960 ;
        RECT 2332.730 1594.160 2333.050 1594.220 ;
        RECT 2332.535 1594.020 2333.050 1594.160 ;
        RECT 2332.730 1593.960 2333.050 1594.020 ;
        RECT 2332.270 1559.140 2332.590 1559.200 ;
        RECT 2333.190 1559.140 2333.510 1559.200 ;
        RECT 2332.270 1559.000 2333.510 1559.140 ;
        RECT 2332.270 1558.940 2332.590 1559.000 ;
        RECT 2333.190 1558.940 2333.510 1559.000 ;
        RECT 2332.745 1545.540 2333.035 1545.585 ;
        RECT 2333.190 1545.540 2333.510 1545.600 ;
        RECT 2332.745 1545.400 2333.510 1545.540 ;
        RECT 2332.745 1545.355 2333.035 1545.400 ;
        RECT 2333.190 1545.340 2333.510 1545.400 ;
        RECT 2332.730 1497.600 2333.050 1497.660 ;
        RECT 2332.535 1497.460 2333.050 1497.600 ;
        RECT 2332.730 1497.400 2333.050 1497.460 ;
        RECT 2332.270 1462.580 2332.590 1462.640 ;
        RECT 2333.190 1462.580 2333.510 1462.640 ;
        RECT 2332.270 1462.440 2333.510 1462.580 ;
        RECT 2332.270 1462.380 2332.590 1462.440 ;
        RECT 2333.190 1462.380 2333.510 1462.440 ;
        RECT 2332.730 1400.700 2333.050 1400.760 ;
        RECT 2332.535 1400.560 2333.050 1400.700 ;
        RECT 2332.730 1400.500 2333.050 1400.560 ;
        RECT 2332.745 1352.760 2333.035 1352.805 ;
        RECT 2333.190 1352.760 2333.510 1352.820 ;
        RECT 2332.745 1352.620 2333.510 1352.760 ;
        RECT 2332.745 1352.575 2333.035 1352.620 ;
        RECT 2333.190 1352.560 2333.510 1352.620 ;
        RECT 2332.730 1304.140 2333.050 1304.200 ;
        RECT 2332.535 1304.000 2333.050 1304.140 ;
        RECT 2332.730 1303.940 2333.050 1304.000 ;
        RECT 2332.745 1256.200 2333.035 1256.245 ;
        RECT 2333.190 1256.200 2333.510 1256.260 ;
        RECT 2332.745 1256.060 2333.510 1256.200 ;
        RECT 2332.745 1256.015 2333.035 1256.060 ;
        RECT 2333.190 1256.000 2333.510 1256.060 ;
        RECT 2332.730 1207.240 2333.050 1207.300 ;
        RECT 2333.190 1207.240 2333.510 1207.300 ;
        RECT 2332.730 1207.100 2333.510 1207.240 ;
        RECT 2332.730 1207.040 2333.050 1207.100 ;
        RECT 2333.190 1207.040 2333.510 1207.100 ;
        RECT 2332.730 1110.680 2333.050 1110.740 ;
        RECT 2333.190 1110.680 2333.510 1110.740 ;
        RECT 2332.730 1110.540 2333.510 1110.680 ;
        RECT 2332.730 1110.480 2333.050 1110.540 ;
        RECT 2333.190 1110.480 2333.510 1110.540 ;
        RECT 2332.730 1014.120 2333.050 1014.180 ;
        RECT 2333.190 1014.120 2333.510 1014.180 ;
        RECT 2332.730 1013.980 2333.510 1014.120 ;
        RECT 2332.730 1013.920 2333.050 1013.980 ;
        RECT 2333.190 1013.920 2333.510 1013.980 ;
        RECT 2332.730 917.560 2333.050 917.620 ;
        RECT 2333.190 917.560 2333.510 917.620 ;
        RECT 2332.730 917.420 2333.510 917.560 ;
        RECT 2332.730 917.360 2333.050 917.420 ;
        RECT 2333.190 917.360 2333.510 917.420 ;
        RECT 2332.730 773.060 2333.050 773.120 ;
        RECT 2333.190 773.060 2333.510 773.120 ;
        RECT 2332.730 772.920 2333.510 773.060 ;
        RECT 2332.730 772.860 2333.050 772.920 ;
        RECT 2333.190 772.860 2333.510 772.920 ;
        RECT 2332.730 772.380 2333.050 772.440 ;
        RECT 2332.535 772.240 2333.050 772.380 ;
        RECT 2332.730 772.180 2333.050 772.240 ;
        RECT 2332.730 738.040 2333.050 738.100 ;
        RECT 2332.535 737.900 2333.050 738.040 ;
        RECT 2332.730 737.840 2333.050 737.900 ;
        RECT 2332.270 690.100 2332.590 690.160 ;
        RECT 2333.190 690.100 2333.510 690.160 ;
        RECT 2332.270 689.960 2333.510 690.100 ;
        RECT 2332.270 689.900 2332.590 689.960 ;
        RECT 2333.190 689.900 2333.510 689.960 ;
        RECT 2332.270 641.620 2332.590 641.880 ;
        RECT 2332.360 641.480 2332.500 641.620 ;
        RECT 2332.730 641.480 2333.050 641.540 ;
        RECT 2332.360 641.340 2333.050 641.480 ;
        RECT 2332.730 641.280 2333.050 641.340 ;
        RECT 2333.190 627.880 2333.510 627.940 ;
        RECT 2333.650 627.880 2333.970 627.940 ;
        RECT 2333.190 627.740 2333.970 627.880 ;
        RECT 2333.190 627.680 2333.510 627.740 ;
        RECT 2333.650 627.680 2333.970 627.740 ;
        RECT 2333.205 620.740 2333.495 620.785 ;
        RECT 2333.650 620.740 2333.970 620.800 ;
        RECT 2333.205 620.600 2333.970 620.740 ;
        RECT 2333.205 620.555 2333.495 620.600 ;
        RECT 2333.650 620.540 2333.970 620.600 ;
        RECT 2333.190 572.800 2333.510 572.860 ;
        RECT 2332.995 572.660 2333.510 572.800 ;
        RECT 2333.190 572.600 2333.510 572.660 ;
        RECT 2333.190 545.260 2333.510 545.320 ;
        RECT 2332.820 545.120 2333.510 545.260 ;
        RECT 2332.820 544.980 2332.960 545.120 ;
        RECT 2333.190 545.060 2333.510 545.120 ;
        RECT 2332.730 544.720 2333.050 544.980 ;
        RECT 2332.730 496.780 2333.050 497.040 ;
        RECT 2332.270 496.640 2332.590 496.700 ;
        RECT 2332.820 496.640 2332.960 496.780 ;
        RECT 2332.270 496.500 2332.960 496.640 ;
        RECT 2332.270 496.440 2332.590 496.500 ;
        RECT 2332.730 427.620 2333.050 427.680 ;
        RECT 2332.535 427.480 2333.050 427.620 ;
        RECT 2332.730 427.420 2333.050 427.480 ;
        RECT 2332.745 379.680 2333.035 379.725 ;
        RECT 2333.190 379.680 2333.510 379.740 ;
        RECT 2332.745 379.540 2333.510 379.680 ;
        RECT 2332.745 379.495 2333.035 379.540 ;
        RECT 2333.190 379.480 2333.510 379.540 ;
        RECT 2332.270 331.060 2332.590 331.120 ;
        RECT 2332.075 330.920 2332.590 331.060 ;
        RECT 2332.270 330.860 2332.590 330.920 ;
        RECT 2332.285 283.120 2332.575 283.165 ;
        RECT 2334.110 283.120 2334.430 283.180 ;
        RECT 2332.285 282.980 2334.430 283.120 ;
        RECT 2332.285 282.935 2332.575 282.980 ;
        RECT 2334.110 282.920 2334.430 282.980 ;
        RECT 2333.190 241.640 2333.510 241.700 ;
        RECT 2334.110 241.640 2334.430 241.700 ;
        RECT 2333.190 241.500 2334.430 241.640 ;
        RECT 2333.190 241.440 2333.510 241.500 ;
        RECT 2334.110 241.440 2334.430 241.500 ;
        RECT 2332.730 145.080 2333.050 145.140 ;
        RECT 2333.190 145.080 2333.510 145.140 ;
        RECT 2332.730 144.940 2333.510 145.080 ;
        RECT 2332.730 144.880 2333.050 144.940 ;
        RECT 2333.190 144.880 2333.510 144.940 ;
        RECT 2310.190 17.240 2310.510 17.300 ;
        RECT 2332.270 17.240 2332.590 17.300 ;
        RECT 2310.190 17.100 2332.590 17.240 ;
        RECT 2310.190 17.040 2310.510 17.100 ;
        RECT 2332.270 17.040 2332.590 17.100 ;
      LAYER via ;
        RECT 2332.760 1666.380 2333.020 1666.640 ;
        RECT 2335.520 1666.380 2335.780 1666.640 ;
        RECT 2332.760 1607.900 2333.020 1608.160 ;
        RECT 2332.760 1593.960 2333.020 1594.220 ;
        RECT 2332.300 1558.940 2332.560 1559.200 ;
        RECT 2333.220 1558.940 2333.480 1559.200 ;
        RECT 2333.220 1545.340 2333.480 1545.600 ;
        RECT 2332.760 1497.400 2333.020 1497.660 ;
        RECT 2332.300 1462.380 2332.560 1462.640 ;
        RECT 2333.220 1462.380 2333.480 1462.640 ;
        RECT 2332.760 1400.500 2333.020 1400.760 ;
        RECT 2333.220 1352.560 2333.480 1352.820 ;
        RECT 2332.760 1303.940 2333.020 1304.200 ;
        RECT 2333.220 1256.000 2333.480 1256.260 ;
        RECT 2332.760 1207.040 2333.020 1207.300 ;
        RECT 2333.220 1207.040 2333.480 1207.300 ;
        RECT 2332.760 1110.480 2333.020 1110.740 ;
        RECT 2333.220 1110.480 2333.480 1110.740 ;
        RECT 2332.760 1013.920 2333.020 1014.180 ;
        RECT 2333.220 1013.920 2333.480 1014.180 ;
        RECT 2332.760 917.360 2333.020 917.620 ;
        RECT 2333.220 917.360 2333.480 917.620 ;
        RECT 2332.760 772.860 2333.020 773.120 ;
        RECT 2333.220 772.860 2333.480 773.120 ;
        RECT 2332.760 772.180 2333.020 772.440 ;
        RECT 2332.760 737.840 2333.020 738.100 ;
        RECT 2332.300 689.900 2332.560 690.160 ;
        RECT 2333.220 689.900 2333.480 690.160 ;
        RECT 2332.300 641.620 2332.560 641.880 ;
        RECT 2332.760 641.280 2333.020 641.540 ;
        RECT 2333.220 627.680 2333.480 627.940 ;
        RECT 2333.680 627.680 2333.940 627.940 ;
        RECT 2333.680 620.540 2333.940 620.800 ;
        RECT 2333.220 572.600 2333.480 572.860 ;
        RECT 2333.220 545.060 2333.480 545.320 ;
        RECT 2332.760 544.720 2333.020 544.980 ;
        RECT 2332.760 496.780 2333.020 497.040 ;
        RECT 2332.300 496.440 2332.560 496.700 ;
        RECT 2332.760 427.420 2333.020 427.680 ;
        RECT 2333.220 379.480 2333.480 379.740 ;
        RECT 2332.300 330.860 2332.560 331.120 ;
        RECT 2334.140 282.920 2334.400 283.180 ;
        RECT 2333.220 241.440 2333.480 241.700 ;
        RECT 2334.140 241.440 2334.400 241.700 ;
        RECT 2332.760 144.880 2333.020 145.140 ;
        RECT 2333.220 144.880 2333.480 145.140 ;
        RECT 2310.220 17.040 2310.480 17.300 ;
        RECT 2332.300 17.040 2332.560 17.300 ;
      LAYER met2 ;
        RECT 2337.740 1700.410 2338.020 1702.400 ;
        RECT 2335.580 1700.270 2338.020 1700.410 ;
        RECT 2335.580 1666.670 2335.720 1700.270 ;
        RECT 2337.740 1700.000 2338.020 1700.270 ;
        RECT 2332.760 1666.350 2333.020 1666.670 ;
        RECT 2335.520 1666.350 2335.780 1666.670 ;
        RECT 2332.820 1608.190 2332.960 1666.350 ;
        RECT 2332.760 1607.870 2333.020 1608.190 ;
        RECT 2332.760 1593.930 2333.020 1594.250 ;
        RECT 2332.820 1559.650 2332.960 1593.930 ;
        RECT 2332.360 1559.510 2332.960 1559.650 ;
        RECT 2332.360 1559.230 2332.500 1559.510 ;
        RECT 2332.300 1558.910 2332.560 1559.230 ;
        RECT 2333.220 1558.910 2333.480 1559.230 ;
        RECT 2333.280 1545.630 2333.420 1558.910 ;
        RECT 2333.220 1545.310 2333.480 1545.630 ;
        RECT 2332.760 1497.370 2333.020 1497.690 ;
        RECT 2332.820 1463.090 2332.960 1497.370 ;
        RECT 2332.360 1462.950 2332.960 1463.090 ;
        RECT 2332.360 1462.670 2332.500 1462.950 ;
        RECT 2332.300 1462.350 2332.560 1462.670 ;
        RECT 2333.220 1462.350 2333.480 1462.670 ;
        RECT 2333.280 1401.210 2333.420 1462.350 ;
        RECT 2332.820 1401.070 2333.420 1401.210 ;
        RECT 2332.820 1400.790 2332.960 1401.070 ;
        RECT 2332.760 1400.470 2333.020 1400.790 ;
        RECT 2333.220 1352.530 2333.480 1352.850 ;
        RECT 2333.280 1317.570 2333.420 1352.530 ;
        RECT 2332.820 1317.430 2333.420 1317.570 ;
        RECT 2332.820 1304.230 2332.960 1317.430 ;
        RECT 2332.760 1303.910 2333.020 1304.230 ;
        RECT 2333.220 1255.970 2333.480 1256.290 ;
        RECT 2333.280 1221.010 2333.420 1255.970 ;
        RECT 2332.820 1220.870 2333.420 1221.010 ;
        RECT 2332.820 1207.330 2332.960 1220.870 ;
        RECT 2332.760 1207.010 2333.020 1207.330 ;
        RECT 2333.220 1207.010 2333.480 1207.330 ;
        RECT 2333.280 1124.450 2333.420 1207.010 ;
        RECT 2332.820 1124.310 2333.420 1124.450 ;
        RECT 2332.820 1110.770 2332.960 1124.310 ;
        RECT 2332.760 1110.450 2333.020 1110.770 ;
        RECT 2333.220 1110.450 2333.480 1110.770 ;
        RECT 2333.280 1027.890 2333.420 1110.450 ;
        RECT 2332.820 1027.750 2333.420 1027.890 ;
        RECT 2332.820 1014.210 2332.960 1027.750 ;
        RECT 2332.760 1013.890 2333.020 1014.210 ;
        RECT 2333.220 1013.890 2333.480 1014.210 ;
        RECT 2333.280 931.330 2333.420 1013.890 ;
        RECT 2332.820 931.190 2333.420 931.330 ;
        RECT 2332.820 917.650 2332.960 931.190 ;
        RECT 2332.760 917.330 2333.020 917.650 ;
        RECT 2333.220 917.330 2333.480 917.650 ;
        RECT 2333.280 834.770 2333.420 917.330 ;
        RECT 2332.820 834.630 2333.420 834.770 ;
        RECT 2332.820 786.490 2332.960 834.630 ;
        RECT 2332.820 786.350 2333.420 786.490 ;
        RECT 2333.280 773.150 2333.420 786.350 ;
        RECT 2332.760 772.830 2333.020 773.150 ;
        RECT 2333.220 772.830 2333.480 773.150 ;
        RECT 2332.820 772.470 2332.960 772.830 ;
        RECT 2332.760 772.150 2333.020 772.470 ;
        RECT 2332.760 737.810 2333.020 738.130 ;
        RECT 2332.820 724.610 2332.960 737.810 ;
        RECT 2332.820 724.470 2333.420 724.610 ;
        RECT 2333.280 690.190 2333.420 724.470 ;
        RECT 2332.300 689.870 2332.560 690.190 ;
        RECT 2333.220 689.870 2333.480 690.190 ;
        RECT 2332.360 641.910 2332.500 689.870 ;
        RECT 2332.300 641.590 2332.560 641.910 ;
        RECT 2332.760 641.250 2333.020 641.570 ;
        RECT 2332.820 628.050 2332.960 641.250 ;
        RECT 2332.820 627.970 2333.420 628.050 ;
        RECT 2332.820 627.910 2333.480 627.970 ;
        RECT 2333.220 627.650 2333.480 627.910 ;
        RECT 2333.680 627.650 2333.940 627.970 ;
        RECT 2333.740 620.830 2333.880 627.650 ;
        RECT 2333.680 620.510 2333.940 620.830 ;
        RECT 2333.220 572.570 2333.480 572.890 ;
        RECT 2333.280 545.350 2333.420 572.570 ;
        RECT 2333.220 545.030 2333.480 545.350 ;
        RECT 2332.760 544.690 2333.020 545.010 ;
        RECT 2332.820 497.070 2332.960 544.690 ;
        RECT 2332.760 496.750 2333.020 497.070 ;
        RECT 2332.300 496.410 2332.560 496.730 ;
        RECT 2332.360 483.325 2332.500 496.410 ;
        RECT 2332.290 482.955 2332.570 483.325 ;
        RECT 2333.210 482.955 2333.490 483.325 ;
        RECT 2333.280 448.530 2333.420 482.955 ;
        RECT 2332.820 448.390 2333.420 448.530 ;
        RECT 2332.820 427.710 2332.960 448.390 ;
        RECT 2332.760 427.390 2333.020 427.710 ;
        RECT 2333.220 379.450 2333.480 379.770 ;
        RECT 2333.280 338.370 2333.420 379.450 ;
        RECT 2332.360 338.230 2333.420 338.370 ;
        RECT 2332.360 331.150 2332.500 338.230 ;
        RECT 2332.300 330.830 2332.560 331.150 ;
        RECT 2334.140 282.890 2334.400 283.210 ;
        RECT 2334.200 241.730 2334.340 282.890 ;
        RECT 2333.220 241.410 2333.480 241.730 ;
        RECT 2334.140 241.410 2334.400 241.730 ;
        RECT 2333.280 145.170 2333.420 241.410 ;
        RECT 2332.760 144.850 2333.020 145.170 ;
        RECT 2333.220 144.850 2333.480 145.170 ;
        RECT 2332.820 110.570 2332.960 144.850 ;
        RECT 2332.820 110.430 2333.420 110.570 ;
        RECT 2333.280 62.290 2333.420 110.430 ;
        RECT 2332.360 62.150 2333.420 62.290 ;
        RECT 2332.360 17.330 2332.500 62.150 ;
        RECT 2310.220 17.010 2310.480 17.330 ;
        RECT 2332.300 17.010 2332.560 17.330 ;
        RECT 2310.280 2.400 2310.420 17.010 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
      LAYER via2 ;
        RECT 2332.290 483.000 2332.570 483.280 ;
        RECT 2333.210 483.000 2333.490 483.280 ;
      LAYER met3 ;
        RECT 2332.265 483.290 2332.595 483.305 ;
        RECT 2333.185 483.290 2333.515 483.305 ;
        RECT 2332.265 482.990 2333.515 483.290 ;
        RECT 2332.265 482.975 2332.595 482.990 ;
        RECT 2333.185 482.975 2333.515 482.990 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2331.810 1688.340 2332.130 1688.400 ;
        RECT 2346.990 1688.340 2347.310 1688.400 ;
        RECT 2331.810 1688.200 2347.310 1688.340 ;
        RECT 2331.810 1688.140 2332.130 1688.200 ;
        RECT 2346.990 1688.140 2347.310 1688.200 ;
        RECT 2328.130 14.520 2328.450 14.580 ;
        RECT 2331.810 14.520 2332.130 14.580 ;
        RECT 2328.130 14.380 2332.130 14.520 ;
        RECT 2328.130 14.320 2328.450 14.380 ;
        RECT 2331.810 14.320 2332.130 14.380 ;
      LAYER via ;
        RECT 2331.840 1688.140 2332.100 1688.400 ;
        RECT 2347.020 1688.140 2347.280 1688.400 ;
        RECT 2328.160 14.320 2328.420 14.580 ;
        RECT 2331.840 14.320 2332.100 14.580 ;
      LAYER met2 ;
        RECT 2346.940 1700.000 2347.220 1702.400 ;
        RECT 2347.080 1688.430 2347.220 1700.000 ;
        RECT 2331.840 1688.110 2332.100 1688.430 ;
        RECT 2347.020 1688.110 2347.280 1688.430 ;
        RECT 2331.900 14.610 2332.040 1688.110 ;
        RECT 2328.160 14.290 2328.420 14.610 ;
        RECT 2331.840 14.290 2332.100 14.610 ;
        RECT 2328.220 2.400 2328.360 14.290 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2349.290 1683.920 2349.610 1683.980 ;
        RECT 2356.190 1683.920 2356.510 1683.980 ;
        RECT 2349.290 1683.780 2356.510 1683.920 ;
        RECT 2349.290 1683.720 2349.610 1683.780 ;
        RECT 2356.190 1683.720 2356.510 1683.780 ;
        RECT 2345.610 20.640 2345.930 20.700 ;
        RECT 2349.290 20.640 2349.610 20.700 ;
        RECT 2345.610 20.500 2349.610 20.640 ;
        RECT 2345.610 20.440 2345.930 20.500 ;
        RECT 2349.290 20.440 2349.610 20.500 ;
      LAYER via ;
        RECT 2349.320 1683.720 2349.580 1683.980 ;
        RECT 2356.220 1683.720 2356.480 1683.980 ;
        RECT 2345.640 20.440 2345.900 20.700 ;
        RECT 2349.320 20.440 2349.580 20.700 ;
      LAYER met2 ;
        RECT 2356.140 1700.000 2356.420 1702.400 ;
        RECT 2356.280 1684.010 2356.420 1700.000 ;
        RECT 2349.320 1683.690 2349.580 1684.010 ;
        RECT 2356.220 1683.690 2356.480 1684.010 ;
        RECT 2349.380 20.730 2349.520 1683.690 ;
        RECT 2345.640 20.410 2345.900 20.730 ;
        RECT 2349.320 20.410 2349.580 20.730 ;
        RECT 2345.700 2.400 2345.840 20.410 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2360.405 1594.005 2360.575 1642.115 ;
        RECT 2360.405 1497.445 2360.575 1545.555 ;
        RECT 2360.405 1352.605 2360.575 1400.715 ;
        RECT 2360.405 1256.045 2360.575 1304.155 ;
        RECT 2360.405 641.325 2360.575 717.655 ;
        RECT 2360.405 338.045 2360.575 403.835 ;
        RECT 2360.405 241.485 2360.575 289.595 ;
        RECT 2360.405 144.925 2360.575 193.035 ;
      LAYER mcon ;
        RECT 2360.405 1641.945 2360.575 1642.115 ;
        RECT 2360.405 1545.385 2360.575 1545.555 ;
        RECT 2360.405 1400.545 2360.575 1400.715 ;
        RECT 2360.405 1303.985 2360.575 1304.155 ;
        RECT 2360.405 717.485 2360.575 717.655 ;
        RECT 2360.405 403.665 2360.575 403.835 ;
        RECT 2360.405 289.425 2360.575 289.595 ;
        RECT 2360.405 192.865 2360.575 193.035 ;
      LAYER met1 ;
        RECT 2360.345 1642.100 2360.635 1642.145 ;
        RECT 2360.790 1642.100 2361.110 1642.160 ;
        RECT 2360.345 1641.960 2361.110 1642.100 ;
        RECT 2360.345 1641.915 2360.635 1641.960 ;
        RECT 2360.790 1641.900 2361.110 1641.960 ;
        RECT 2360.330 1594.160 2360.650 1594.220 ;
        RECT 2360.135 1594.020 2360.650 1594.160 ;
        RECT 2360.330 1593.960 2360.650 1594.020 ;
        RECT 2359.870 1559.140 2360.190 1559.200 ;
        RECT 2360.790 1559.140 2361.110 1559.200 ;
        RECT 2359.870 1559.000 2361.110 1559.140 ;
        RECT 2359.870 1558.940 2360.190 1559.000 ;
        RECT 2360.790 1558.940 2361.110 1559.000 ;
        RECT 2360.345 1545.540 2360.635 1545.585 ;
        RECT 2360.790 1545.540 2361.110 1545.600 ;
        RECT 2360.345 1545.400 2361.110 1545.540 ;
        RECT 2360.345 1545.355 2360.635 1545.400 ;
        RECT 2360.790 1545.340 2361.110 1545.400 ;
        RECT 2360.330 1497.600 2360.650 1497.660 ;
        RECT 2360.135 1497.460 2360.650 1497.600 ;
        RECT 2360.330 1497.400 2360.650 1497.460 ;
        RECT 2359.870 1462.580 2360.190 1462.640 ;
        RECT 2360.790 1462.580 2361.110 1462.640 ;
        RECT 2359.870 1462.440 2361.110 1462.580 ;
        RECT 2359.870 1462.380 2360.190 1462.440 ;
        RECT 2360.790 1462.380 2361.110 1462.440 ;
        RECT 2360.330 1400.700 2360.650 1400.760 ;
        RECT 2360.135 1400.560 2360.650 1400.700 ;
        RECT 2360.330 1400.500 2360.650 1400.560 ;
        RECT 2360.345 1352.760 2360.635 1352.805 ;
        RECT 2360.790 1352.760 2361.110 1352.820 ;
        RECT 2360.345 1352.620 2361.110 1352.760 ;
        RECT 2360.345 1352.575 2360.635 1352.620 ;
        RECT 2360.790 1352.560 2361.110 1352.620 ;
        RECT 2360.330 1304.140 2360.650 1304.200 ;
        RECT 2360.135 1304.000 2360.650 1304.140 ;
        RECT 2360.330 1303.940 2360.650 1304.000 ;
        RECT 2360.345 1256.200 2360.635 1256.245 ;
        RECT 2360.790 1256.200 2361.110 1256.260 ;
        RECT 2360.345 1256.060 2361.110 1256.200 ;
        RECT 2360.345 1256.015 2360.635 1256.060 ;
        RECT 2360.790 1256.000 2361.110 1256.060 ;
        RECT 2360.790 1159.300 2361.110 1159.360 ;
        RECT 2361.710 1159.300 2362.030 1159.360 ;
        RECT 2360.790 1159.160 2362.030 1159.300 ;
        RECT 2360.790 1159.100 2361.110 1159.160 ;
        RECT 2361.710 1159.100 2362.030 1159.160 ;
        RECT 2360.790 1062.740 2361.110 1062.800 ;
        RECT 2361.710 1062.740 2362.030 1062.800 ;
        RECT 2360.790 1062.600 2362.030 1062.740 ;
        RECT 2360.790 1062.540 2361.110 1062.600 ;
        RECT 2361.710 1062.540 2362.030 1062.600 ;
        RECT 2360.790 966.180 2361.110 966.240 ;
        RECT 2361.710 966.180 2362.030 966.240 ;
        RECT 2360.790 966.040 2362.030 966.180 ;
        RECT 2360.790 965.980 2361.110 966.040 ;
        RECT 2361.710 965.980 2362.030 966.040 ;
        RECT 2360.790 869.620 2361.110 869.680 ;
        RECT 2361.710 869.620 2362.030 869.680 ;
        RECT 2360.790 869.480 2362.030 869.620 ;
        RECT 2360.790 869.420 2361.110 869.480 ;
        RECT 2361.710 869.420 2362.030 869.480 ;
        RECT 2360.330 821.000 2360.650 821.060 ;
        RECT 2361.710 821.000 2362.030 821.060 ;
        RECT 2360.330 820.860 2362.030 821.000 ;
        RECT 2360.330 820.800 2360.650 820.860 ;
        RECT 2361.710 820.800 2362.030 820.860 ;
        RECT 2360.330 717.640 2360.650 717.700 ;
        RECT 2360.135 717.500 2360.650 717.640 ;
        RECT 2360.330 717.440 2360.650 717.500 ;
        RECT 2360.330 641.480 2360.650 641.540 ;
        RECT 2360.135 641.340 2360.650 641.480 ;
        RECT 2360.330 641.280 2360.650 641.340 ;
        RECT 2360.330 593.340 2360.650 593.600 ;
        RECT 2359.870 593.200 2360.190 593.260 ;
        RECT 2360.420 593.200 2360.560 593.340 ;
        RECT 2359.870 593.060 2360.560 593.200 ;
        RECT 2359.870 593.000 2360.190 593.060 ;
        RECT 2360.330 496.780 2360.650 497.040 ;
        RECT 2359.870 496.640 2360.190 496.700 ;
        RECT 2360.420 496.640 2360.560 496.780 ;
        RECT 2359.870 496.500 2360.560 496.640 ;
        RECT 2359.870 496.440 2360.190 496.500 ;
        RECT 2360.330 403.820 2360.650 403.880 ;
        RECT 2360.135 403.680 2360.650 403.820 ;
        RECT 2360.330 403.620 2360.650 403.680 ;
        RECT 2360.330 338.200 2360.650 338.260 ;
        RECT 2360.135 338.060 2360.650 338.200 ;
        RECT 2360.330 338.000 2360.650 338.060 ;
        RECT 2359.870 303.520 2360.190 303.580 ;
        RECT 2360.790 303.520 2361.110 303.580 ;
        RECT 2359.870 303.380 2361.110 303.520 ;
        RECT 2359.870 303.320 2360.190 303.380 ;
        RECT 2360.790 303.320 2361.110 303.380 ;
        RECT 2360.345 289.580 2360.635 289.625 ;
        RECT 2360.790 289.580 2361.110 289.640 ;
        RECT 2360.345 289.440 2361.110 289.580 ;
        RECT 2360.345 289.395 2360.635 289.440 ;
        RECT 2360.790 289.380 2361.110 289.440 ;
        RECT 2360.330 241.640 2360.650 241.700 ;
        RECT 2360.135 241.500 2360.650 241.640 ;
        RECT 2360.330 241.440 2360.650 241.500 ;
        RECT 2359.870 206.960 2360.190 207.020 ;
        RECT 2360.790 206.960 2361.110 207.020 ;
        RECT 2359.870 206.820 2361.110 206.960 ;
        RECT 2359.870 206.760 2360.190 206.820 ;
        RECT 2360.790 206.760 2361.110 206.820 ;
        RECT 2360.345 193.020 2360.635 193.065 ;
        RECT 2360.790 193.020 2361.110 193.080 ;
        RECT 2360.345 192.880 2361.110 193.020 ;
        RECT 2360.345 192.835 2360.635 192.880 ;
        RECT 2360.790 192.820 2361.110 192.880 ;
        RECT 2360.330 145.080 2360.650 145.140 ;
        RECT 2360.135 144.940 2360.650 145.080 ;
        RECT 2360.330 144.880 2360.650 144.940 ;
        RECT 2360.790 20.640 2361.110 20.700 ;
        RECT 2363.550 20.640 2363.870 20.700 ;
        RECT 2360.790 20.500 2363.870 20.640 ;
        RECT 2360.790 20.440 2361.110 20.500 ;
        RECT 2363.550 20.440 2363.870 20.500 ;
      LAYER via ;
        RECT 2360.820 1641.900 2361.080 1642.160 ;
        RECT 2360.360 1593.960 2360.620 1594.220 ;
        RECT 2359.900 1558.940 2360.160 1559.200 ;
        RECT 2360.820 1558.940 2361.080 1559.200 ;
        RECT 2360.820 1545.340 2361.080 1545.600 ;
        RECT 2360.360 1497.400 2360.620 1497.660 ;
        RECT 2359.900 1462.380 2360.160 1462.640 ;
        RECT 2360.820 1462.380 2361.080 1462.640 ;
        RECT 2360.360 1400.500 2360.620 1400.760 ;
        RECT 2360.820 1352.560 2361.080 1352.820 ;
        RECT 2360.360 1303.940 2360.620 1304.200 ;
        RECT 2360.820 1256.000 2361.080 1256.260 ;
        RECT 2360.820 1159.100 2361.080 1159.360 ;
        RECT 2361.740 1159.100 2362.000 1159.360 ;
        RECT 2360.820 1062.540 2361.080 1062.800 ;
        RECT 2361.740 1062.540 2362.000 1062.800 ;
        RECT 2360.820 965.980 2361.080 966.240 ;
        RECT 2361.740 965.980 2362.000 966.240 ;
        RECT 2360.820 869.420 2361.080 869.680 ;
        RECT 2361.740 869.420 2362.000 869.680 ;
        RECT 2360.360 820.800 2360.620 821.060 ;
        RECT 2361.740 820.800 2362.000 821.060 ;
        RECT 2360.360 717.440 2360.620 717.700 ;
        RECT 2360.360 641.280 2360.620 641.540 ;
        RECT 2360.360 593.340 2360.620 593.600 ;
        RECT 2359.900 593.000 2360.160 593.260 ;
        RECT 2360.360 496.780 2360.620 497.040 ;
        RECT 2359.900 496.440 2360.160 496.700 ;
        RECT 2360.360 403.620 2360.620 403.880 ;
        RECT 2360.360 338.000 2360.620 338.260 ;
        RECT 2359.900 303.320 2360.160 303.580 ;
        RECT 2360.820 303.320 2361.080 303.580 ;
        RECT 2360.820 289.380 2361.080 289.640 ;
        RECT 2360.360 241.440 2360.620 241.700 ;
        RECT 2359.900 206.760 2360.160 207.020 ;
        RECT 2360.820 206.760 2361.080 207.020 ;
        RECT 2360.820 192.820 2361.080 193.080 ;
        RECT 2360.360 144.880 2360.620 145.140 ;
        RECT 2360.820 20.440 2361.080 20.700 ;
        RECT 2363.580 20.440 2363.840 20.700 ;
      LAYER met2 ;
        RECT 2365.340 1700.410 2365.620 1702.400 ;
        RECT 2362.720 1700.270 2365.620 1700.410 ;
        RECT 2362.720 1666.410 2362.860 1700.270 ;
        RECT 2365.340 1700.000 2365.620 1700.270 ;
        RECT 2360.880 1666.270 2362.860 1666.410 ;
        RECT 2360.880 1642.190 2361.020 1666.270 ;
        RECT 2360.820 1641.870 2361.080 1642.190 ;
        RECT 2360.360 1593.930 2360.620 1594.250 ;
        RECT 2360.420 1559.650 2360.560 1593.930 ;
        RECT 2359.960 1559.510 2360.560 1559.650 ;
        RECT 2359.960 1559.230 2360.100 1559.510 ;
        RECT 2359.900 1558.910 2360.160 1559.230 ;
        RECT 2360.820 1558.910 2361.080 1559.230 ;
        RECT 2360.880 1545.630 2361.020 1558.910 ;
        RECT 2360.820 1545.310 2361.080 1545.630 ;
        RECT 2360.360 1497.370 2360.620 1497.690 ;
        RECT 2360.420 1463.090 2360.560 1497.370 ;
        RECT 2359.960 1462.950 2360.560 1463.090 ;
        RECT 2359.960 1462.670 2360.100 1462.950 ;
        RECT 2359.900 1462.350 2360.160 1462.670 ;
        RECT 2360.820 1462.350 2361.080 1462.670 ;
        RECT 2360.880 1401.210 2361.020 1462.350 ;
        RECT 2360.420 1401.070 2361.020 1401.210 ;
        RECT 2360.420 1400.790 2360.560 1401.070 ;
        RECT 2360.360 1400.470 2360.620 1400.790 ;
        RECT 2360.820 1352.530 2361.080 1352.850 ;
        RECT 2360.880 1317.570 2361.020 1352.530 ;
        RECT 2360.420 1317.430 2361.020 1317.570 ;
        RECT 2360.420 1304.230 2360.560 1317.430 ;
        RECT 2360.360 1303.910 2360.620 1304.230 ;
        RECT 2360.820 1255.970 2361.080 1256.290 ;
        RECT 2360.880 1221.010 2361.020 1255.970 ;
        RECT 2360.420 1220.870 2361.020 1221.010 ;
        RECT 2360.420 1207.525 2360.560 1220.870 ;
        RECT 2360.350 1207.155 2360.630 1207.525 ;
        RECT 2361.730 1207.155 2362.010 1207.525 ;
        RECT 2361.800 1159.390 2361.940 1207.155 ;
        RECT 2360.820 1159.070 2361.080 1159.390 ;
        RECT 2361.740 1159.070 2362.000 1159.390 ;
        RECT 2360.880 1124.450 2361.020 1159.070 ;
        RECT 2360.420 1124.310 2361.020 1124.450 ;
        RECT 2360.420 1110.965 2360.560 1124.310 ;
        RECT 2360.350 1110.595 2360.630 1110.965 ;
        RECT 2361.730 1110.595 2362.010 1110.965 ;
        RECT 2361.800 1062.830 2361.940 1110.595 ;
        RECT 2360.820 1062.510 2361.080 1062.830 ;
        RECT 2361.740 1062.510 2362.000 1062.830 ;
        RECT 2360.880 1027.890 2361.020 1062.510 ;
        RECT 2360.420 1027.750 2361.020 1027.890 ;
        RECT 2360.420 1014.405 2360.560 1027.750 ;
        RECT 2360.350 1014.035 2360.630 1014.405 ;
        RECT 2361.730 1014.035 2362.010 1014.405 ;
        RECT 2361.800 966.270 2361.940 1014.035 ;
        RECT 2360.820 965.950 2361.080 966.270 ;
        RECT 2361.740 965.950 2362.000 966.270 ;
        RECT 2360.880 931.330 2361.020 965.950 ;
        RECT 2360.420 931.190 2361.020 931.330 ;
        RECT 2360.420 917.845 2360.560 931.190 ;
        RECT 2360.350 917.475 2360.630 917.845 ;
        RECT 2361.730 917.475 2362.010 917.845 ;
        RECT 2361.800 869.710 2361.940 917.475 ;
        RECT 2360.820 869.390 2361.080 869.710 ;
        RECT 2361.740 869.390 2362.000 869.710 ;
        RECT 2360.880 834.770 2361.020 869.390 ;
        RECT 2360.420 834.630 2361.020 834.770 ;
        RECT 2360.420 821.090 2360.560 834.630 ;
        RECT 2360.360 820.770 2360.620 821.090 ;
        RECT 2361.740 820.770 2362.000 821.090 ;
        RECT 2361.800 773.005 2361.940 820.770 ;
        RECT 2360.810 772.635 2361.090 773.005 ;
        RECT 2361.730 772.635 2362.010 773.005 ;
        RECT 2360.880 738.210 2361.020 772.635 ;
        RECT 2360.420 738.070 2361.020 738.210 ;
        RECT 2360.420 717.730 2360.560 738.070 ;
        RECT 2360.360 717.410 2360.620 717.730 ;
        RECT 2360.360 641.250 2360.620 641.570 ;
        RECT 2360.420 593.630 2360.560 641.250 ;
        RECT 2360.360 593.310 2360.620 593.630 ;
        RECT 2359.900 592.970 2360.160 593.290 ;
        RECT 2359.960 579.885 2360.100 592.970 ;
        RECT 2359.890 579.515 2360.170 579.885 ;
        RECT 2360.810 579.515 2361.090 579.885 ;
        RECT 2360.880 545.090 2361.020 579.515 ;
        RECT 2360.420 544.950 2361.020 545.090 ;
        RECT 2360.420 497.070 2360.560 544.950 ;
        RECT 2360.360 496.750 2360.620 497.070 ;
        RECT 2359.900 496.410 2360.160 496.730 ;
        RECT 2359.960 483.325 2360.100 496.410 ;
        RECT 2359.890 482.955 2360.170 483.325 ;
        RECT 2360.810 482.955 2361.090 483.325 ;
        RECT 2360.880 448.530 2361.020 482.955 ;
        RECT 2360.420 448.390 2361.020 448.530 ;
        RECT 2360.420 403.910 2360.560 448.390 ;
        RECT 2360.360 403.590 2360.620 403.910 ;
        RECT 2360.360 337.970 2360.620 338.290 ;
        RECT 2360.420 303.690 2360.560 337.970 ;
        RECT 2359.960 303.610 2360.560 303.690 ;
        RECT 2359.900 303.550 2360.560 303.610 ;
        RECT 2359.900 303.290 2360.160 303.550 ;
        RECT 2360.820 303.290 2361.080 303.610 ;
        RECT 2360.880 289.670 2361.020 303.290 ;
        RECT 2360.820 289.350 2361.080 289.670 ;
        RECT 2360.360 241.410 2360.620 241.730 ;
        RECT 2360.420 207.130 2360.560 241.410 ;
        RECT 2359.960 207.050 2360.560 207.130 ;
        RECT 2359.900 206.990 2360.560 207.050 ;
        RECT 2359.900 206.730 2360.160 206.990 ;
        RECT 2360.820 206.730 2361.080 207.050 ;
        RECT 2360.880 193.110 2361.020 206.730 ;
        RECT 2360.820 192.790 2361.080 193.110 ;
        RECT 2360.360 144.850 2360.620 145.170 ;
        RECT 2360.420 120.770 2360.560 144.850 ;
        RECT 2360.420 120.630 2361.020 120.770 ;
        RECT 2360.880 20.730 2361.020 120.630 ;
        RECT 2360.820 20.410 2361.080 20.730 ;
        RECT 2363.580 20.410 2363.840 20.730 ;
        RECT 2363.640 2.400 2363.780 20.410 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
      LAYER via2 ;
        RECT 2360.350 1207.200 2360.630 1207.480 ;
        RECT 2361.730 1207.200 2362.010 1207.480 ;
        RECT 2360.350 1110.640 2360.630 1110.920 ;
        RECT 2361.730 1110.640 2362.010 1110.920 ;
        RECT 2360.350 1014.080 2360.630 1014.360 ;
        RECT 2361.730 1014.080 2362.010 1014.360 ;
        RECT 2360.350 917.520 2360.630 917.800 ;
        RECT 2361.730 917.520 2362.010 917.800 ;
        RECT 2360.810 772.680 2361.090 772.960 ;
        RECT 2361.730 772.680 2362.010 772.960 ;
        RECT 2359.890 579.560 2360.170 579.840 ;
        RECT 2360.810 579.560 2361.090 579.840 ;
        RECT 2359.890 483.000 2360.170 483.280 ;
        RECT 2360.810 483.000 2361.090 483.280 ;
      LAYER met3 ;
        RECT 2360.325 1207.490 2360.655 1207.505 ;
        RECT 2361.705 1207.490 2362.035 1207.505 ;
        RECT 2360.325 1207.190 2362.035 1207.490 ;
        RECT 2360.325 1207.175 2360.655 1207.190 ;
        RECT 2361.705 1207.175 2362.035 1207.190 ;
        RECT 2360.325 1110.930 2360.655 1110.945 ;
        RECT 2361.705 1110.930 2362.035 1110.945 ;
        RECT 2360.325 1110.630 2362.035 1110.930 ;
        RECT 2360.325 1110.615 2360.655 1110.630 ;
        RECT 2361.705 1110.615 2362.035 1110.630 ;
        RECT 2360.325 1014.370 2360.655 1014.385 ;
        RECT 2361.705 1014.370 2362.035 1014.385 ;
        RECT 2360.325 1014.070 2362.035 1014.370 ;
        RECT 2360.325 1014.055 2360.655 1014.070 ;
        RECT 2361.705 1014.055 2362.035 1014.070 ;
        RECT 2360.325 917.810 2360.655 917.825 ;
        RECT 2361.705 917.810 2362.035 917.825 ;
        RECT 2360.325 917.510 2362.035 917.810 ;
        RECT 2360.325 917.495 2360.655 917.510 ;
        RECT 2361.705 917.495 2362.035 917.510 ;
        RECT 2360.785 772.970 2361.115 772.985 ;
        RECT 2361.705 772.970 2362.035 772.985 ;
        RECT 2360.785 772.670 2362.035 772.970 ;
        RECT 2360.785 772.655 2361.115 772.670 ;
        RECT 2361.705 772.655 2362.035 772.670 ;
        RECT 2359.865 579.850 2360.195 579.865 ;
        RECT 2360.785 579.850 2361.115 579.865 ;
        RECT 2359.865 579.550 2361.115 579.850 ;
        RECT 2359.865 579.535 2360.195 579.550 ;
        RECT 2360.785 579.535 2361.115 579.550 ;
        RECT 2359.865 483.290 2360.195 483.305 ;
        RECT 2360.785 483.290 2361.115 483.305 ;
        RECT 2359.865 482.990 2361.115 483.290 ;
        RECT 2359.865 482.975 2360.195 482.990 ;
        RECT 2360.785 482.975 2361.115 482.990 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2374.590 1683.920 2374.910 1683.980 ;
        RECT 2380.110 1683.920 2380.430 1683.980 ;
        RECT 2374.590 1683.780 2380.430 1683.920 ;
        RECT 2374.590 1683.720 2374.910 1683.780 ;
        RECT 2380.110 1683.720 2380.430 1683.780 ;
      LAYER via ;
        RECT 2374.620 1683.720 2374.880 1683.980 ;
        RECT 2380.140 1683.720 2380.400 1683.980 ;
      LAYER met2 ;
        RECT 2374.540 1700.000 2374.820 1702.400 ;
        RECT 2374.680 1684.010 2374.820 1700.000 ;
        RECT 2374.620 1683.690 2374.880 1684.010 ;
        RECT 2380.140 1683.690 2380.400 1684.010 ;
        RECT 2380.200 17.410 2380.340 1683.690 ;
        RECT 2380.200 17.270 2381.720 17.410 ;
        RECT 2381.580 2.400 2381.720 17.270 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2387.010 15.200 2387.330 15.260 ;
        RECT 2399.430 15.200 2399.750 15.260 ;
        RECT 2387.010 15.060 2399.750 15.200 ;
        RECT 2387.010 15.000 2387.330 15.060 ;
        RECT 2399.430 15.000 2399.750 15.060 ;
      LAYER via ;
        RECT 2387.040 15.000 2387.300 15.260 ;
        RECT 2399.460 15.000 2399.720 15.260 ;
      LAYER met2 ;
        RECT 2383.740 1700.410 2384.020 1702.400 ;
        RECT 2383.740 1700.270 2386.320 1700.410 ;
        RECT 2383.740 1700.000 2384.020 1700.270 ;
        RECT 2386.180 1688.680 2386.320 1700.270 ;
        RECT 2386.180 1688.540 2387.240 1688.680 ;
        RECT 2387.100 15.290 2387.240 1688.540 ;
        RECT 2387.040 14.970 2387.300 15.290 ;
        RECT 2399.460 14.970 2399.720 15.290 ;
        RECT 2399.520 2.400 2399.660 14.970 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1553.565 1449.165 1553.735 1497.275 ;
        RECT 1553.565 1352.605 1553.735 1400.715 ;
        RECT 1553.565 1256.045 1553.735 1304.155 ;
        RECT 1553.565 579.785 1553.735 627.895 ;
        RECT 1553.565 483.225 1553.735 531.335 ;
        RECT 1553.565 386.325 1553.735 434.775 ;
        RECT 1552.645 206.805 1552.815 234.515 ;
      LAYER mcon ;
        RECT 1553.565 1497.105 1553.735 1497.275 ;
        RECT 1553.565 1400.545 1553.735 1400.715 ;
        RECT 1553.565 1303.985 1553.735 1304.155 ;
        RECT 1553.565 627.725 1553.735 627.895 ;
        RECT 1553.565 531.165 1553.735 531.335 ;
        RECT 1553.565 434.605 1553.735 434.775 ;
        RECT 1552.645 234.345 1552.815 234.515 ;
      LAYER met1 ;
        RECT 1553.490 1678.140 1553.810 1678.200 ;
        RECT 1555.790 1678.140 1556.110 1678.200 ;
        RECT 1553.490 1678.000 1556.110 1678.140 ;
        RECT 1553.490 1677.940 1553.810 1678.000 ;
        RECT 1555.790 1677.940 1556.110 1678.000 ;
        RECT 1553.490 1497.260 1553.810 1497.320 ;
        RECT 1553.295 1497.120 1553.810 1497.260 ;
        RECT 1553.490 1497.060 1553.810 1497.120 ;
        RECT 1553.490 1449.320 1553.810 1449.380 ;
        RECT 1553.295 1449.180 1553.810 1449.320 ;
        RECT 1553.490 1449.120 1553.810 1449.180 ;
        RECT 1553.490 1400.700 1553.810 1400.760 ;
        RECT 1553.295 1400.560 1553.810 1400.700 ;
        RECT 1553.490 1400.500 1553.810 1400.560 ;
        RECT 1553.490 1352.760 1553.810 1352.820 ;
        RECT 1553.295 1352.620 1553.810 1352.760 ;
        RECT 1553.490 1352.560 1553.810 1352.620 ;
        RECT 1553.490 1304.140 1553.810 1304.200 ;
        RECT 1553.295 1304.000 1553.810 1304.140 ;
        RECT 1553.490 1303.940 1553.810 1304.000 ;
        RECT 1553.490 1256.200 1553.810 1256.260 ;
        RECT 1553.295 1256.060 1553.810 1256.200 ;
        RECT 1553.490 1256.000 1553.810 1256.060 ;
        RECT 1553.490 1159.300 1553.810 1159.360 ;
        RECT 1554.410 1159.300 1554.730 1159.360 ;
        RECT 1553.490 1159.160 1554.730 1159.300 ;
        RECT 1553.490 1159.100 1553.810 1159.160 ;
        RECT 1554.410 1159.100 1554.730 1159.160 ;
        RECT 1553.490 1062.740 1553.810 1062.800 ;
        RECT 1554.410 1062.740 1554.730 1062.800 ;
        RECT 1553.490 1062.600 1554.730 1062.740 ;
        RECT 1553.490 1062.540 1553.810 1062.600 ;
        RECT 1554.410 1062.540 1554.730 1062.600 ;
        RECT 1553.490 966.180 1553.810 966.240 ;
        RECT 1554.410 966.180 1554.730 966.240 ;
        RECT 1553.490 966.040 1554.730 966.180 ;
        RECT 1553.490 965.980 1553.810 966.040 ;
        RECT 1554.410 965.980 1554.730 966.040 ;
        RECT 1553.490 821.000 1553.810 821.060 ;
        RECT 1554.410 821.000 1554.730 821.060 ;
        RECT 1553.490 820.860 1554.730 821.000 ;
        RECT 1553.490 820.800 1553.810 820.860 ;
        RECT 1554.410 820.800 1554.730 820.860 ;
        RECT 1553.490 724.440 1553.810 724.500 ;
        RECT 1554.410 724.440 1554.730 724.500 ;
        RECT 1553.490 724.300 1554.730 724.440 ;
        RECT 1553.490 724.240 1553.810 724.300 ;
        RECT 1554.410 724.240 1554.730 724.300 ;
        RECT 1553.490 627.880 1553.810 627.940 ;
        RECT 1553.295 627.740 1553.810 627.880 ;
        RECT 1553.490 627.680 1553.810 627.740 ;
        RECT 1553.490 579.940 1553.810 580.000 ;
        RECT 1553.295 579.800 1553.810 579.940 ;
        RECT 1553.490 579.740 1553.810 579.800 ;
        RECT 1553.490 531.320 1553.810 531.380 ;
        RECT 1553.295 531.180 1553.810 531.320 ;
        RECT 1553.490 531.120 1553.810 531.180 ;
        RECT 1553.490 483.380 1553.810 483.440 ;
        RECT 1553.295 483.240 1553.810 483.380 ;
        RECT 1553.490 483.180 1553.810 483.240 ;
        RECT 1553.490 434.760 1553.810 434.820 ;
        RECT 1553.295 434.620 1553.810 434.760 ;
        RECT 1553.490 434.560 1553.810 434.620 ;
        RECT 1553.490 386.480 1553.810 386.540 ;
        RECT 1553.295 386.340 1553.810 386.480 ;
        RECT 1553.490 386.280 1553.810 386.340 ;
        RECT 1552.585 234.500 1552.875 234.545 ;
        RECT 1553.030 234.500 1553.350 234.560 ;
        RECT 1552.585 234.360 1553.350 234.500 ;
        RECT 1552.585 234.315 1552.875 234.360 ;
        RECT 1553.030 234.300 1553.350 234.360 ;
        RECT 1552.585 206.960 1552.875 207.005 ;
        RECT 1553.030 206.960 1553.350 207.020 ;
        RECT 1552.585 206.820 1553.350 206.960 ;
        RECT 1552.585 206.775 1552.875 206.820 ;
        RECT 1553.030 206.760 1553.350 206.820 ;
        RECT 1552.110 96.800 1552.430 96.860 ;
        RECT 1553.490 96.800 1553.810 96.860 ;
        RECT 1552.110 96.660 1553.810 96.800 ;
        RECT 1552.110 96.600 1552.430 96.660 ;
        RECT 1553.490 96.600 1553.810 96.660 ;
        RECT 799.550 68.580 799.870 68.640 ;
        RECT 1553.490 68.580 1553.810 68.640 ;
        RECT 799.550 68.440 1553.810 68.580 ;
        RECT 799.550 68.380 799.870 68.440 ;
        RECT 1553.490 68.380 1553.810 68.440 ;
        RECT 793.570 20.980 793.890 21.040 ;
        RECT 799.550 20.980 799.870 21.040 ;
        RECT 793.570 20.840 799.870 20.980 ;
        RECT 793.570 20.780 793.890 20.840 ;
        RECT 799.550 20.780 799.870 20.840 ;
      LAYER via ;
        RECT 1553.520 1677.940 1553.780 1678.200 ;
        RECT 1555.820 1677.940 1556.080 1678.200 ;
        RECT 1553.520 1497.060 1553.780 1497.320 ;
        RECT 1553.520 1449.120 1553.780 1449.380 ;
        RECT 1553.520 1400.500 1553.780 1400.760 ;
        RECT 1553.520 1352.560 1553.780 1352.820 ;
        RECT 1553.520 1303.940 1553.780 1304.200 ;
        RECT 1553.520 1256.000 1553.780 1256.260 ;
        RECT 1553.520 1159.100 1553.780 1159.360 ;
        RECT 1554.440 1159.100 1554.700 1159.360 ;
        RECT 1553.520 1062.540 1553.780 1062.800 ;
        RECT 1554.440 1062.540 1554.700 1062.800 ;
        RECT 1553.520 965.980 1553.780 966.240 ;
        RECT 1554.440 965.980 1554.700 966.240 ;
        RECT 1553.520 820.800 1553.780 821.060 ;
        RECT 1554.440 820.800 1554.700 821.060 ;
        RECT 1553.520 724.240 1553.780 724.500 ;
        RECT 1554.440 724.240 1554.700 724.500 ;
        RECT 1553.520 627.680 1553.780 627.940 ;
        RECT 1553.520 579.740 1553.780 580.000 ;
        RECT 1553.520 531.120 1553.780 531.380 ;
        RECT 1553.520 483.180 1553.780 483.440 ;
        RECT 1553.520 434.560 1553.780 434.820 ;
        RECT 1553.520 386.280 1553.780 386.540 ;
        RECT 1553.060 234.300 1553.320 234.560 ;
        RECT 1553.060 206.760 1553.320 207.020 ;
        RECT 1552.140 96.600 1552.400 96.860 ;
        RECT 1553.520 96.600 1553.780 96.860 ;
        RECT 799.580 68.380 799.840 68.640 ;
        RECT 1553.520 68.380 1553.780 68.640 ;
        RECT 793.600 20.780 793.860 21.040 ;
        RECT 799.580 20.780 799.840 21.040 ;
      LAYER met2 ;
        RECT 1557.120 1700.410 1557.400 1702.400 ;
        RECT 1555.880 1700.270 1557.400 1700.410 ;
        RECT 1555.880 1678.230 1556.020 1700.270 ;
        RECT 1557.120 1700.000 1557.400 1700.270 ;
        RECT 1553.520 1677.910 1553.780 1678.230 ;
        RECT 1555.820 1677.910 1556.080 1678.230 ;
        RECT 1553.580 1559.650 1553.720 1677.910 ;
        RECT 1553.120 1559.510 1553.720 1559.650 ;
        RECT 1553.120 1558.970 1553.260 1559.510 ;
        RECT 1553.120 1558.830 1553.720 1558.970 ;
        RECT 1553.580 1497.350 1553.720 1558.830 ;
        RECT 1553.520 1497.030 1553.780 1497.350 ;
        RECT 1553.520 1449.090 1553.780 1449.410 ;
        RECT 1553.580 1400.790 1553.720 1449.090 ;
        RECT 1553.520 1400.470 1553.780 1400.790 ;
        RECT 1553.520 1352.530 1553.780 1352.850 ;
        RECT 1553.580 1304.230 1553.720 1352.530 ;
        RECT 1553.520 1303.910 1553.780 1304.230 ;
        RECT 1553.520 1255.970 1553.780 1256.290 ;
        RECT 1553.580 1207.525 1553.720 1255.970 ;
        RECT 1553.510 1207.155 1553.790 1207.525 ;
        RECT 1554.430 1207.155 1554.710 1207.525 ;
        RECT 1554.500 1159.390 1554.640 1207.155 ;
        RECT 1553.520 1159.070 1553.780 1159.390 ;
        RECT 1554.440 1159.070 1554.700 1159.390 ;
        RECT 1553.580 1110.965 1553.720 1159.070 ;
        RECT 1553.510 1110.595 1553.790 1110.965 ;
        RECT 1554.430 1110.595 1554.710 1110.965 ;
        RECT 1554.500 1062.830 1554.640 1110.595 ;
        RECT 1553.520 1062.510 1553.780 1062.830 ;
        RECT 1554.440 1062.510 1554.700 1062.830 ;
        RECT 1553.580 1014.405 1553.720 1062.510 ;
        RECT 1553.510 1014.035 1553.790 1014.405 ;
        RECT 1554.430 1014.035 1554.710 1014.405 ;
        RECT 1554.500 966.270 1554.640 1014.035 ;
        RECT 1553.520 965.950 1553.780 966.270 ;
        RECT 1554.440 965.950 1554.700 966.270 ;
        RECT 1553.580 883.730 1553.720 965.950 ;
        RECT 1553.120 883.590 1553.720 883.730 ;
        RECT 1553.120 883.050 1553.260 883.590 ;
        RECT 1553.120 882.910 1553.720 883.050 ;
        RECT 1553.580 821.090 1553.720 882.910 ;
        RECT 1553.520 820.770 1553.780 821.090 ;
        RECT 1554.440 820.770 1554.700 821.090 ;
        RECT 1554.500 773.005 1554.640 820.770 ;
        RECT 1553.510 772.635 1553.790 773.005 ;
        RECT 1554.430 772.635 1554.710 773.005 ;
        RECT 1553.580 724.530 1553.720 772.635 ;
        RECT 1553.520 724.210 1553.780 724.530 ;
        RECT 1554.440 724.210 1554.700 724.530 ;
        RECT 1554.500 676.445 1554.640 724.210 ;
        RECT 1553.510 676.075 1553.790 676.445 ;
        RECT 1554.430 676.075 1554.710 676.445 ;
        RECT 1553.580 627.970 1553.720 676.075 ;
        RECT 1553.520 627.650 1553.780 627.970 ;
        RECT 1553.520 579.710 1553.780 580.030 ;
        RECT 1553.580 531.410 1553.720 579.710 ;
        RECT 1553.520 531.090 1553.780 531.410 ;
        RECT 1553.520 483.150 1553.780 483.470 ;
        RECT 1553.580 434.850 1553.720 483.150 ;
        RECT 1553.520 434.530 1553.780 434.850 ;
        RECT 1553.520 386.250 1553.780 386.570 ;
        RECT 1553.580 303.180 1553.720 386.250 ;
        RECT 1553.120 303.040 1553.720 303.180 ;
        RECT 1553.120 302.330 1553.260 303.040 ;
        RECT 1553.120 302.190 1553.720 302.330 ;
        RECT 1553.580 242.605 1553.720 302.190 ;
        RECT 1553.510 242.235 1553.790 242.605 ;
        RECT 1553.050 241.555 1553.330 241.925 ;
        RECT 1553.120 234.590 1553.260 241.555 ;
        RECT 1553.060 234.270 1553.320 234.590 ;
        RECT 1553.060 206.730 1553.320 207.050 ;
        RECT 1553.120 144.685 1553.260 206.730 ;
        RECT 1552.130 144.315 1552.410 144.685 ;
        RECT 1553.050 144.315 1553.330 144.685 ;
        RECT 1552.200 96.890 1552.340 144.315 ;
        RECT 1552.140 96.570 1552.400 96.890 ;
        RECT 1553.520 96.570 1553.780 96.890 ;
        RECT 1553.580 68.670 1553.720 96.570 ;
        RECT 799.580 68.350 799.840 68.670 ;
        RECT 1553.520 68.350 1553.780 68.670 ;
        RECT 799.640 21.070 799.780 68.350 ;
        RECT 793.600 20.750 793.860 21.070 ;
        RECT 799.580 20.750 799.840 21.070 ;
        RECT 793.660 2.400 793.800 20.750 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 1553.510 1207.200 1553.790 1207.480 ;
        RECT 1554.430 1207.200 1554.710 1207.480 ;
        RECT 1553.510 1110.640 1553.790 1110.920 ;
        RECT 1554.430 1110.640 1554.710 1110.920 ;
        RECT 1553.510 1014.080 1553.790 1014.360 ;
        RECT 1554.430 1014.080 1554.710 1014.360 ;
        RECT 1553.510 772.680 1553.790 772.960 ;
        RECT 1554.430 772.680 1554.710 772.960 ;
        RECT 1553.510 676.120 1553.790 676.400 ;
        RECT 1554.430 676.120 1554.710 676.400 ;
        RECT 1553.510 242.280 1553.790 242.560 ;
        RECT 1553.050 241.600 1553.330 241.880 ;
        RECT 1552.130 144.360 1552.410 144.640 ;
        RECT 1553.050 144.360 1553.330 144.640 ;
      LAYER met3 ;
        RECT 1553.485 1207.490 1553.815 1207.505 ;
        RECT 1554.405 1207.490 1554.735 1207.505 ;
        RECT 1553.485 1207.190 1554.735 1207.490 ;
        RECT 1553.485 1207.175 1553.815 1207.190 ;
        RECT 1554.405 1207.175 1554.735 1207.190 ;
        RECT 1553.485 1110.930 1553.815 1110.945 ;
        RECT 1554.405 1110.930 1554.735 1110.945 ;
        RECT 1553.485 1110.630 1554.735 1110.930 ;
        RECT 1553.485 1110.615 1553.815 1110.630 ;
        RECT 1554.405 1110.615 1554.735 1110.630 ;
        RECT 1553.485 1014.370 1553.815 1014.385 ;
        RECT 1554.405 1014.370 1554.735 1014.385 ;
        RECT 1553.485 1014.070 1554.735 1014.370 ;
        RECT 1553.485 1014.055 1553.815 1014.070 ;
        RECT 1554.405 1014.055 1554.735 1014.070 ;
        RECT 1553.485 772.970 1553.815 772.985 ;
        RECT 1554.405 772.970 1554.735 772.985 ;
        RECT 1553.485 772.670 1554.735 772.970 ;
        RECT 1553.485 772.655 1553.815 772.670 ;
        RECT 1554.405 772.655 1554.735 772.670 ;
        RECT 1553.485 676.410 1553.815 676.425 ;
        RECT 1554.405 676.410 1554.735 676.425 ;
        RECT 1553.485 676.110 1554.735 676.410 ;
        RECT 1553.485 676.095 1553.815 676.110 ;
        RECT 1554.405 676.095 1554.735 676.110 ;
        RECT 1553.485 242.570 1553.815 242.585 ;
        RECT 1552.350 242.270 1553.815 242.570 ;
        RECT 1552.350 241.890 1552.650 242.270 ;
        RECT 1553.485 242.255 1553.815 242.270 ;
        RECT 1553.025 241.890 1553.355 241.905 ;
        RECT 1552.350 241.590 1553.355 241.890 ;
        RECT 1553.025 241.575 1553.355 241.590 ;
        RECT 1552.105 144.650 1552.435 144.665 ;
        RECT 1553.025 144.650 1553.355 144.665 ;
        RECT 1552.105 144.350 1553.355 144.650 ;
        RECT 1552.105 144.335 1552.435 144.350 ;
        RECT 1553.025 144.335 1553.355 144.350 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.310 59.060 641.630 59.120 ;
        RECT 1476.670 59.060 1476.990 59.120 ;
        RECT 641.310 58.920 1476.990 59.060 ;
        RECT 641.310 58.860 641.630 58.920 ;
        RECT 1476.670 58.860 1476.990 58.920 ;
      LAYER via ;
        RECT 641.340 58.860 641.600 59.120 ;
        RECT 1476.700 58.860 1476.960 59.120 ;
      LAYER met2 ;
        RECT 1477.540 1700.410 1477.820 1702.400 ;
        RECT 1476.760 1700.270 1477.820 1700.410 ;
        RECT 1476.760 59.150 1476.900 1700.270 ;
        RECT 1477.540 1700.000 1477.820 1700.270 ;
        RECT 641.340 58.830 641.600 59.150 ;
        RECT 1476.700 58.830 1476.960 59.150 ;
        RECT 641.400 17.410 641.540 58.830 ;
        RECT 639.100 17.270 641.540 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2395.750 1688.680 2396.070 1688.740 ;
        RECT 2395.750 1688.540 2401.500 1688.680 ;
        RECT 2395.750 1688.480 2396.070 1688.540 ;
        RECT 2401.360 1688.340 2401.500 1688.540 ;
        RECT 2401.360 1688.200 2416.680 1688.340 ;
        RECT 2416.540 1688.000 2416.680 1688.200 ;
        RECT 2422.890 1688.000 2423.210 1688.060 ;
        RECT 2416.540 1687.860 2423.210 1688.000 ;
        RECT 2422.890 1687.800 2423.210 1687.860 ;
      LAYER via ;
        RECT 2395.780 1688.480 2396.040 1688.740 ;
        RECT 2422.920 1687.800 2423.180 1688.060 ;
      LAYER met2 ;
        RECT 2395.700 1700.000 2395.980 1702.400 ;
        RECT 2395.840 1688.770 2395.980 1700.000 ;
        RECT 2395.780 1688.450 2396.040 1688.770 ;
        RECT 2422.920 1687.770 2423.180 1688.090 ;
        RECT 2422.980 2.400 2423.120 1687.770 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2404.950 1687.320 2405.270 1687.380 ;
        RECT 2425.190 1687.320 2425.510 1687.380 ;
        RECT 2404.950 1687.180 2425.510 1687.320 ;
        RECT 2404.950 1687.120 2405.270 1687.180 ;
        RECT 2425.190 1687.120 2425.510 1687.180 ;
        RECT 2425.190 16.220 2425.510 16.280 ;
        RECT 2440.830 16.220 2441.150 16.280 ;
        RECT 2425.190 16.080 2441.150 16.220 ;
        RECT 2425.190 16.020 2425.510 16.080 ;
        RECT 2440.830 16.020 2441.150 16.080 ;
      LAYER via ;
        RECT 2404.980 1687.120 2405.240 1687.380 ;
        RECT 2425.220 1687.120 2425.480 1687.380 ;
        RECT 2425.220 16.020 2425.480 16.280 ;
        RECT 2440.860 16.020 2441.120 16.280 ;
      LAYER met2 ;
        RECT 2404.900 1700.000 2405.180 1702.400 ;
        RECT 2405.040 1687.410 2405.180 1700.000 ;
        RECT 2404.980 1687.090 2405.240 1687.410 ;
        RECT 2425.220 1687.090 2425.480 1687.410 ;
        RECT 2425.280 16.310 2425.420 1687.090 ;
        RECT 2425.220 15.990 2425.480 16.310 ;
        RECT 2440.860 15.990 2441.120 16.310 ;
        RECT 2440.920 2.400 2441.060 15.990 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2431.705 1686.825 2431.875 1689.035 ;
      LAYER mcon ;
        RECT 2431.705 1688.865 2431.875 1689.035 ;
      LAYER met1 ;
        RECT 2414.150 1689.020 2414.470 1689.080 ;
        RECT 2431.645 1689.020 2431.935 1689.065 ;
        RECT 2414.150 1688.880 2431.935 1689.020 ;
        RECT 2414.150 1688.820 2414.470 1688.880 ;
        RECT 2431.645 1688.835 2431.935 1688.880 ;
        RECT 2431.645 1686.980 2431.935 1687.025 ;
        RECT 2457.390 1686.980 2457.710 1687.040 ;
        RECT 2431.645 1686.840 2457.710 1686.980 ;
        RECT 2431.645 1686.795 2431.935 1686.840 ;
        RECT 2457.390 1686.780 2457.710 1686.840 ;
      LAYER via ;
        RECT 2414.180 1688.820 2414.440 1689.080 ;
        RECT 2457.420 1686.780 2457.680 1687.040 ;
      LAYER met2 ;
        RECT 2414.100 1700.000 2414.380 1702.400 ;
        RECT 2414.240 1689.110 2414.380 1700.000 ;
        RECT 2414.180 1688.790 2414.440 1689.110 ;
        RECT 2457.420 1686.750 2457.680 1687.070 ;
        RECT 2457.480 3.130 2457.620 1686.750 ;
        RECT 2457.480 2.990 2458.540 3.130 ;
        RECT 2458.400 2.960 2458.540 2.990 ;
        RECT 2458.400 2.820 2459.000 2.960 ;
        RECT 2458.860 2.400 2459.000 2.820 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2423.350 1686.980 2423.670 1687.040 ;
        RECT 2428.410 1686.980 2428.730 1687.040 ;
        RECT 2423.350 1686.840 2428.730 1686.980 ;
        RECT 2423.350 1686.780 2423.670 1686.840 ;
        RECT 2428.410 1686.780 2428.730 1686.840 ;
        RECT 2428.410 18.600 2428.730 18.660 ;
        RECT 2476.710 18.600 2477.030 18.660 ;
        RECT 2428.410 18.460 2477.030 18.600 ;
        RECT 2428.410 18.400 2428.730 18.460 ;
        RECT 2476.710 18.400 2477.030 18.460 ;
      LAYER via ;
        RECT 2423.380 1686.780 2423.640 1687.040 ;
        RECT 2428.440 1686.780 2428.700 1687.040 ;
        RECT 2428.440 18.400 2428.700 18.660 ;
        RECT 2476.740 18.400 2477.000 18.660 ;
      LAYER met2 ;
        RECT 2423.300 1700.000 2423.580 1702.400 ;
        RECT 2423.440 1687.070 2423.580 1700.000 ;
        RECT 2423.380 1686.750 2423.640 1687.070 ;
        RECT 2428.440 1686.750 2428.700 1687.070 ;
        RECT 2428.500 18.690 2428.640 1686.750 ;
        RECT 2428.440 18.370 2428.700 18.690 ;
        RECT 2476.740 18.370 2477.000 18.690 ;
        RECT 2476.800 2.400 2476.940 18.370 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2435.310 17.580 2435.630 17.640 ;
        RECT 2494.650 17.580 2494.970 17.640 ;
        RECT 2435.310 17.440 2494.970 17.580 ;
        RECT 2435.310 17.380 2435.630 17.440 ;
        RECT 2494.650 17.380 2494.970 17.440 ;
      LAYER via ;
        RECT 2435.340 17.380 2435.600 17.640 ;
        RECT 2494.680 17.380 2494.940 17.640 ;
      LAYER met2 ;
        RECT 2432.500 1700.410 2432.780 1702.400 ;
        RECT 2432.500 1700.270 2435.540 1700.410 ;
        RECT 2432.500 1700.000 2432.780 1700.270 ;
        RECT 2435.400 17.670 2435.540 1700.270 ;
        RECT 2435.340 17.350 2435.600 17.670 ;
        RECT 2494.680 17.350 2494.940 17.670 ;
        RECT 2494.740 2.400 2494.880 17.350 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2441.750 16.560 2442.070 16.620 ;
        RECT 2512.130 16.560 2512.450 16.620 ;
        RECT 2441.750 16.420 2512.450 16.560 ;
        RECT 2441.750 16.360 2442.070 16.420 ;
        RECT 2512.130 16.360 2512.450 16.420 ;
      LAYER via ;
        RECT 2441.780 16.360 2442.040 16.620 ;
        RECT 2512.160 16.360 2512.420 16.620 ;
      LAYER met2 ;
        RECT 2441.700 1700.000 2441.980 1702.400 ;
        RECT 2441.840 16.650 2441.980 1700.000 ;
        RECT 2441.780 16.330 2442.040 16.650 ;
        RECT 2512.160 16.330 2512.420 16.650 ;
        RECT 2512.220 2.400 2512.360 16.330 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2450.950 1689.700 2451.270 1689.760 ;
        RECT 2507.990 1689.700 2508.310 1689.760 ;
        RECT 2450.950 1689.560 2508.310 1689.700 ;
        RECT 2450.950 1689.500 2451.270 1689.560 ;
        RECT 2507.990 1689.500 2508.310 1689.560 ;
        RECT 2507.990 15.540 2508.310 15.600 ;
        RECT 2530.070 15.540 2530.390 15.600 ;
        RECT 2507.990 15.400 2530.390 15.540 ;
        RECT 2507.990 15.340 2508.310 15.400 ;
        RECT 2530.070 15.340 2530.390 15.400 ;
      LAYER via ;
        RECT 2450.980 1689.500 2451.240 1689.760 ;
        RECT 2508.020 1689.500 2508.280 1689.760 ;
        RECT 2508.020 15.340 2508.280 15.600 ;
        RECT 2530.100 15.340 2530.360 15.600 ;
      LAYER met2 ;
        RECT 2450.900 1700.000 2451.180 1702.400 ;
        RECT 2451.040 1689.790 2451.180 1700.000 ;
        RECT 2450.980 1689.470 2451.240 1689.790 ;
        RECT 2508.020 1689.470 2508.280 1689.790 ;
        RECT 2508.080 15.630 2508.220 1689.470 ;
        RECT 2508.020 15.310 2508.280 15.630 ;
        RECT 2530.100 15.310 2530.360 15.630 ;
        RECT 2530.160 2.400 2530.300 15.310 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2462.450 20.300 2462.770 20.360 ;
        RECT 2548.010 20.300 2548.330 20.360 ;
        RECT 2462.450 20.160 2548.330 20.300 ;
        RECT 2462.450 20.100 2462.770 20.160 ;
        RECT 2548.010 20.100 2548.330 20.160 ;
      LAYER via ;
        RECT 2462.480 20.100 2462.740 20.360 ;
        RECT 2548.040 20.100 2548.300 20.360 ;
      LAYER met2 ;
        RECT 2460.100 1700.410 2460.380 1702.400 ;
        RECT 2460.100 1700.270 2462.680 1700.410 ;
        RECT 2460.100 1700.000 2460.380 1700.270 ;
        RECT 2462.540 20.390 2462.680 1700.270 ;
        RECT 2462.480 20.070 2462.740 20.390 ;
        RECT 2548.040 20.070 2548.300 20.390 ;
        RECT 2548.100 2.400 2548.240 20.070 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2469.350 19.960 2469.670 20.020 ;
        RECT 2565.950 19.960 2566.270 20.020 ;
        RECT 2469.350 19.820 2566.270 19.960 ;
        RECT 2469.350 19.760 2469.670 19.820 ;
        RECT 2565.950 19.760 2566.270 19.820 ;
      LAYER via ;
        RECT 2469.380 19.760 2469.640 20.020 ;
        RECT 2565.980 19.760 2566.240 20.020 ;
      LAYER met2 ;
        RECT 2469.300 1700.000 2469.580 1702.400 ;
        RECT 2469.440 20.050 2469.580 1700.000 ;
        RECT 2469.380 19.730 2469.640 20.050 ;
        RECT 2565.980 19.730 2566.240 20.050 ;
        RECT 2566.040 2.400 2566.180 19.730 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2548.545 16.745 2548.715 19.295 ;
      LAYER mcon ;
        RECT 2548.545 19.125 2548.715 19.295 ;
      LAYER met1 ;
        RECT 2478.550 1688.000 2478.870 1688.060 ;
        RECT 2483.610 1688.000 2483.930 1688.060 ;
        RECT 2478.550 1687.860 2483.930 1688.000 ;
        RECT 2478.550 1687.800 2478.870 1687.860 ;
        RECT 2483.610 1687.800 2483.930 1687.860 ;
        RECT 2483.610 19.280 2483.930 19.340 ;
        RECT 2548.485 19.280 2548.775 19.325 ;
        RECT 2483.610 19.140 2548.775 19.280 ;
        RECT 2483.610 19.080 2483.930 19.140 ;
        RECT 2548.485 19.095 2548.775 19.140 ;
        RECT 2548.485 16.900 2548.775 16.945 ;
        RECT 2583.890 16.900 2584.210 16.960 ;
        RECT 2548.485 16.760 2584.210 16.900 ;
        RECT 2548.485 16.715 2548.775 16.760 ;
        RECT 2583.890 16.700 2584.210 16.760 ;
      LAYER via ;
        RECT 2478.580 1687.800 2478.840 1688.060 ;
        RECT 2483.640 1687.800 2483.900 1688.060 ;
        RECT 2483.640 19.080 2483.900 19.340 ;
        RECT 2583.920 16.700 2584.180 16.960 ;
      LAYER met2 ;
        RECT 2478.500 1700.000 2478.780 1702.400 ;
        RECT 2478.640 1688.090 2478.780 1700.000 ;
        RECT 2478.580 1687.770 2478.840 1688.090 ;
        RECT 2483.640 1687.770 2483.900 1688.090 ;
        RECT 2483.700 19.370 2483.840 1687.770 ;
        RECT 2483.640 19.050 2483.900 19.370 ;
        RECT 2583.920 16.670 2584.180 16.990 ;
        RECT 2583.980 2.400 2584.120 16.670 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.490 34.240 817.810 34.300 ;
        RECT 1567.750 34.240 1568.070 34.300 ;
        RECT 817.490 34.100 1568.070 34.240 ;
        RECT 817.490 34.040 817.810 34.100 ;
        RECT 1567.750 34.040 1568.070 34.100 ;
      LAYER via ;
        RECT 817.520 34.040 817.780 34.300 ;
        RECT 1567.780 34.040 1568.040 34.300 ;
      LAYER met2 ;
        RECT 1569.080 1700.410 1569.360 1702.400 ;
        RECT 1567.840 1700.270 1569.360 1700.410 ;
        RECT 1567.840 34.330 1567.980 1700.270 ;
        RECT 1569.080 1700.000 1569.360 1700.270 ;
        RECT 817.520 34.010 817.780 34.330 ;
        RECT 1567.780 34.010 1568.040 34.330 ;
        RECT 817.580 2.400 817.720 34.010 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2487.750 1689.020 2488.070 1689.080 ;
        RECT 2549.390 1689.020 2549.710 1689.080 ;
        RECT 2487.750 1688.880 2549.710 1689.020 ;
        RECT 2487.750 1688.820 2488.070 1688.880 ;
        RECT 2549.390 1688.820 2549.710 1688.880 ;
        RECT 2549.390 19.620 2549.710 19.680 ;
        RECT 2601.370 19.620 2601.690 19.680 ;
        RECT 2549.390 19.480 2601.690 19.620 ;
        RECT 2549.390 19.420 2549.710 19.480 ;
        RECT 2601.370 19.420 2601.690 19.480 ;
      LAYER via ;
        RECT 2487.780 1688.820 2488.040 1689.080 ;
        RECT 2549.420 1688.820 2549.680 1689.080 ;
        RECT 2549.420 19.420 2549.680 19.680 ;
        RECT 2601.400 19.420 2601.660 19.680 ;
      LAYER met2 ;
        RECT 2487.700 1700.000 2487.980 1702.400 ;
        RECT 2487.840 1689.110 2487.980 1700.000 ;
        RECT 2487.780 1688.790 2488.040 1689.110 ;
        RECT 2549.420 1688.790 2549.680 1689.110 ;
        RECT 2549.480 19.710 2549.620 1688.790 ;
        RECT 2549.420 19.390 2549.680 19.710 ;
        RECT 2601.400 19.390 2601.660 19.710 ;
        RECT 2601.460 2.400 2601.600 19.390 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2496.950 17.920 2497.270 17.980 ;
        RECT 2619.310 17.920 2619.630 17.980 ;
        RECT 2496.950 17.780 2619.630 17.920 ;
        RECT 2496.950 17.720 2497.270 17.780 ;
        RECT 2619.310 17.720 2619.630 17.780 ;
      LAYER via ;
        RECT 2496.980 17.720 2497.240 17.980 ;
        RECT 2619.340 17.720 2619.600 17.980 ;
      LAYER met2 ;
        RECT 2496.900 1700.000 2497.180 1702.400 ;
        RECT 2497.040 18.010 2497.180 1700.000 ;
        RECT 2496.980 17.690 2497.240 18.010 ;
        RECT 2619.340 17.690 2619.600 18.010 ;
        RECT 2619.400 2.400 2619.540 17.690 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2506.150 1689.360 2506.470 1689.420 ;
        RECT 2506.150 1689.220 2565.260 1689.360 ;
        RECT 2506.150 1689.160 2506.470 1689.220 ;
        RECT 2565.120 1688.340 2565.260 1689.220 ;
        RECT 2583.890 1688.340 2584.210 1688.400 ;
        RECT 2565.120 1688.200 2584.210 1688.340 ;
        RECT 2583.890 1688.140 2584.210 1688.200 ;
        RECT 2583.890 19.280 2584.210 19.340 ;
        RECT 2583.890 19.140 2614.480 19.280 ;
        RECT 2583.890 19.080 2584.210 19.140 ;
        RECT 2614.340 18.600 2614.480 19.140 ;
        RECT 2614.340 18.460 2620.000 18.600 ;
        RECT 2619.860 17.920 2620.000 18.460 ;
        RECT 2637.250 17.920 2637.570 17.980 ;
        RECT 2619.860 17.780 2637.570 17.920 ;
        RECT 2637.250 17.720 2637.570 17.780 ;
      LAYER via ;
        RECT 2506.180 1689.160 2506.440 1689.420 ;
        RECT 2583.920 1688.140 2584.180 1688.400 ;
        RECT 2583.920 19.080 2584.180 19.340 ;
        RECT 2637.280 17.720 2637.540 17.980 ;
      LAYER met2 ;
        RECT 2506.100 1700.000 2506.380 1702.400 ;
        RECT 2506.240 1689.450 2506.380 1700.000 ;
        RECT 2506.180 1689.130 2506.440 1689.450 ;
        RECT 2583.920 1688.110 2584.180 1688.430 ;
        RECT 2583.980 19.370 2584.120 1688.110 ;
        RECT 2583.920 19.050 2584.180 19.370 ;
        RECT 2637.280 17.690 2637.540 18.010 ;
        RECT 2637.340 2.400 2637.480 17.690 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2518.570 14.180 2518.890 14.240 ;
        RECT 2655.190 14.180 2655.510 14.240 ;
        RECT 2518.570 14.040 2655.510 14.180 ;
        RECT 2518.570 13.980 2518.890 14.040 ;
        RECT 2655.190 13.980 2655.510 14.040 ;
      LAYER via ;
        RECT 2518.600 13.980 2518.860 14.240 ;
        RECT 2655.220 13.980 2655.480 14.240 ;
      LAYER met2 ;
        RECT 2515.300 1700.410 2515.580 1702.400 ;
        RECT 2515.300 1700.270 2517.880 1700.410 ;
        RECT 2515.300 1700.000 2515.580 1700.270 ;
        RECT 2517.740 1688.850 2517.880 1700.270 ;
        RECT 2517.740 1688.710 2518.340 1688.850 ;
        RECT 2518.200 17.920 2518.340 1688.710 ;
        RECT 2518.200 17.780 2518.800 17.920 ;
        RECT 2518.660 14.270 2518.800 17.780 ;
        RECT 2518.600 13.950 2518.860 14.270 ;
        RECT 2655.220 13.950 2655.480 14.270 ;
        RECT 2655.280 2.400 2655.420 13.950 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2524.550 1684.600 2524.870 1684.660 ;
        RECT 2670.370 1684.600 2670.690 1684.660 ;
        RECT 2524.550 1684.460 2670.690 1684.600 ;
        RECT 2524.550 1684.400 2524.870 1684.460 ;
        RECT 2670.370 1684.400 2670.690 1684.460 ;
      LAYER via ;
        RECT 2524.580 1684.400 2524.840 1684.660 ;
        RECT 2670.400 1684.400 2670.660 1684.660 ;
      LAYER met2 ;
        RECT 2524.500 1700.000 2524.780 1702.400 ;
        RECT 2524.640 1684.690 2524.780 1700.000 ;
        RECT 2524.580 1684.370 2524.840 1684.690 ;
        RECT 2670.400 1684.370 2670.660 1684.690 ;
        RECT 2670.460 16.730 2670.600 1684.370 ;
        RECT 2670.460 16.590 2672.900 16.730 ;
        RECT 2672.760 2.400 2672.900 16.590 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2533.750 1688.680 2534.070 1688.740 ;
        RECT 2538.810 1688.680 2539.130 1688.740 ;
        RECT 2533.750 1688.540 2539.130 1688.680 ;
        RECT 2533.750 1688.480 2534.070 1688.540 ;
        RECT 2538.810 1688.480 2539.130 1688.540 ;
        RECT 2538.810 15.200 2539.130 15.260 ;
        RECT 2690.610 15.200 2690.930 15.260 ;
        RECT 2538.810 15.060 2690.930 15.200 ;
        RECT 2538.810 15.000 2539.130 15.060 ;
        RECT 2690.610 15.000 2690.930 15.060 ;
      LAYER via ;
        RECT 2533.780 1688.480 2534.040 1688.740 ;
        RECT 2538.840 1688.480 2539.100 1688.740 ;
        RECT 2538.840 15.000 2539.100 15.260 ;
        RECT 2690.640 15.000 2690.900 15.260 ;
      LAYER met2 ;
        RECT 2533.700 1700.000 2533.980 1702.400 ;
        RECT 2533.840 1688.770 2533.980 1700.000 ;
        RECT 2533.780 1688.450 2534.040 1688.770 ;
        RECT 2538.840 1688.450 2539.100 1688.770 ;
        RECT 2538.900 15.290 2539.040 1688.450 ;
        RECT 2538.840 14.970 2539.100 15.290 ;
        RECT 2690.640 14.970 2690.900 15.290 ;
        RECT 2690.700 2.400 2690.840 14.970 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2542.950 1686.300 2543.270 1686.360 ;
        RECT 2701.190 1686.300 2701.510 1686.360 ;
        RECT 2542.950 1686.160 2701.510 1686.300 ;
        RECT 2542.950 1686.100 2543.270 1686.160 ;
        RECT 2701.190 1686.100 2701.510 1686.160 ;
        RECT 2701.190 16.220 2701.510 16.280 ;
        RECT 2708.550 16.220 2708.870 16.280 ;
        RECT 2701.190 16.080 2708.870 16.220 ;
        RECT 2701.190 16.020 2701.510 16.080 ;
        RECT 2708.550 16.020 2708.870 16.080 ;
      LAYER via ;
        RECT 2542.980 1686.100 2543.240 1686.360 ;
        RECT 2701.220 1686.100 2701.480 1686.360 ;
        RECT 2701.220 16.020 2701.480 16.280 ;
        RECT 2708.580 16.020 2708.840 16.280 ;
      LAYER met2 ;
        RECT 2542.900 1700.000 2543.180 1702.400 ;
        RECT 2543.040 1686.390 2543.180 1700.000 ;
        RECT 2542.980 1686.070 2543.240 1686.390 ;
        RECT 2701.220 1686.070 2701.480 1686.390 ;
        RECT 2701.280 16.310 2701.420 1686.070 ;
        RECT 2701.220 15.990 2701.480 16.310 ;
        RECT 2708.580 15.990 2708.840 16.310 ;
        RECT 2708.640 2.400 2708.780 15.990 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2552.610 15.880 2552.930 15.940 ;
        RECT 2552.610 15.740 2701.420 15.880 ;
        RECT 2552.610 15.680 2552.930 15.740 ;
        RECT 2701.280 15.540 2701.420 15.740 ;
        RECT 2726.490 15.540 2726.810 15.600 ;
        RECT 2701.280 15.400 2726.810 15.540 ;
        RECT 2726.490 15.340 2726.810 15.400 ;
      LAYER via ;
        RECT 2552.640 15.680 2552.900 15.940 ;
        RECT 2726.520 15.340 2726.780 15.600 ;
      LAYER met2 ;
        RECT 2552.100 1700.410 2552.380 1702.400 ;
        RECT 2552.100 1700.270 2552.840 1700.410 ;
        RECT 2552.100 1700.000 2552.380 1700.270 ;
        RECT 2552.700 15.970 2552.840 1700.270 ;
        RECT 2552.640 15.650 2552.900 15.970 ;
        RECT 2726.520 15.310 2726.780 15.630 ;
        RECT 2726.580 2.400 2726.720 15.310 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2561.350 1689.700 2561.670 1689.760 ;
        RECT 2736.150 1689.700 2736.470 1689.760 ;
        RECT 2561.350 1689.560 2736.470 1689.700 ;
        RECT 2561.350 1689.500 2561.670 1689.560 ;
        RECT 2736.150 1689.500 2736.470 1689.560 ;
        RECT 2736.150 15.200 2736.470 15.260 ;
        RECT 2744.430 15.200 2744.750 15.260 ;
        RECT 2736.150 15.060 2744.750 15.200 ;
        RECT 2736.150 15.000 2736.470 15.060 ;
        RECT 2744.430 15.000 2744.750 15.060 ;
      LAYER via ;
        RECT 2561.380 1689.500 2561.640 1689.760 ;
        RECT 2736.180 1689.500 2736.440 1689.760 ;
        RECT 2736.180 15.000 2736.440 15.260 ;
        RECT 2744.460 15.000 2744.720 15.260 ;
      LAYER met2 ;
        RECT 2561.300 1700.000 2561.580 1702.400 ;
        RECT 2561.440 1689.790 2561.580 1700.000 ;
        RECT 2561.380 1689.470 2561.640 1689.790 ;
        RECT 2736.180 1689.470 2736.440 1689.790 ;
        RECT 2736.240 15.290 2736.380 1689.470 ;
        RECT 2736.180 14.970 2736.440 15.290 ;
        RECT 2744.460 14.970 2744.720 15.290 ;
        RECT 2744.520 2.400 2744.660 14.970 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2573.310 16.560 2573.630 16.620 ;
        RECT 2761.910 16.560 2762.230 16.620 ;
        RECT 2573.310 16.420 2762.230 16.560 ;
        RECT 2573.310 16.360 2573.630 16.420 ;
        RECT 2761.910 16.360 2762.230 16.420 ;
      LAYER via ;
        RECT 2573.340 16.360 2573.600 16.620 ;
        RECT 2761.940 16.360 2762.200 16.620 ;
      LAYER met2 ;
        RECT 2570.040 1701.090 2570.320 1702.400 ;
        RECT 2570.040 1700.950 2573.080 1701.090 ;
        RECT 2570.040 1700.000 2570.320 1700.950 ;
        RECT 2572.940 1688.680 2573.080 1700.950 ;
        RECT 2572.940 1688.540 2573.540 1688.680 ;
        RECT 2573.400 16.650 2573.540 1688.540 ;
        RECT 2573.340 16.330 2573.600 16.650 ;
        RECT 2761.940 16.330 2762.200 16.650 ;
        RECT 2762.000 2.400 2762.140 16.330 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1573.270 1689.360 1573.590 1689.420 ;
        RECT 1576.950 1689.360 1577.270 1689.420 ;
        RECT 1573.270 1689.220 1577.270 1689.360 ;
        RECT 1573.270 1689.160 1573.590 1689.220 ;
        RECT 1576.950 1689.160 1577.270 1689.220 ;
        RECT 835.430 30.500 835.750 30.560 ;
        RECT 1572.810 30.500 1573.130 30.560 ;
        RECT 835.430 30.360 1573.130 30.500 ;
        RECT 835.430 30.300 835.750 30.360 ;
        RECT 1572.810 30.300 1573.130 30.360 ;
      LAYER via ;
        RECT 1573.300 1689.160 1573.560 1689.420 ;
        RECT 1576.980 1689.160 1577.240 1689.420 ;
        RECT 835.460 30.300 835.720 30.560 ;
        RECT 1572.840 30.300 1573.100 30.560 ;
      LAYER met2 ;
        RECT 1578.280 1700.410 1578.560 1702.400 ;
        RECT 1577.040 1700.270 1578.560 1700.410 ;
        RECT 1577.040 1689.450 1577.180 1700.270 ;
        RECT 1578.280 1700.000 1578.560 1700.270 ;
        RECT 1573.300 1689.130 1573.560 1689.450 ;
        RECT 1576.980 1689.130 1577.240 1689.450 ;
        RECT 1573.360 31.010 1573.500 1689.130 ;
        RECT 1572.900 30.870 1573.500 31.010 ;
        RECT 1572.900 30.590 1573.040 30.870 ;
        RECT 835.460 30.270 835.720 30.590 ;
        RECT 1572.840 30.270 1573.100 30.590 ;
        RECT 835.520 2.400 835.660 30.270 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2579.290 1689.020 2579.610 1689.080 ;
        RECT 2579.290 1688.880 2593.320 1689.020 ;
        RECT 2579.290 1688.820 2579.610 1688.880 ;
        RECT 2593.180 1688.680 2593.320 1688.880 ;
        RECT 2774.330 1688.680 2774.650 1688.740 ;
        RECT 2593.180 1688.540 2774.650 1688.680 ;
        RECT 2774.330 1688.480 2774.650 1688.540 ;
      LAYER via ;
        RECT 2579.320 1688.820 2579.580 1689.080 ;
        RECT 2774.360 1688.480 2774.620 1688.740 ;
      LAYER met2 ;
        RECT 2579.240 1700.000 2579.520 1702.400 ;
        RECT 2579.380 1689.110 2579.520 1700.000 ;
        RECT 2579.320 1688.790 2579.580 1689.110 ;
        RECT 2774.360 1688.450 2774.620 1688.770 ;
        RECT 2774.420 16.730 2774.560 1688.450 ;
        RECT 2774.420 16.590 2780.080 16.730 ;
        RECT 2779.940 2.400 2780.080 16.590 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2588.490 1688.000 2588.810 1688.060 ;
        RECT 2594.010 1688.000 2594.330 1688.060 ;
        RECT 2588.490 1687.860 2594.330 1688.000 ;
        RECT 2588.490 1687.800 2588.810 1687.860 ;
        RECT 2594.010 1687.800 2594.330 1687.860 ;
        RECT 2594.010 20.640 2594.330 20.700 ;
        RECT 2797.790 20.640 2798.110 20.700 ;
        RECT 2594.010 20.500 2798.110 20.640 ;
        RECT 2594.010 20.440 2594.330 20.500 ;
        RECT 2797.790 20.440 2798.110 20.500 ;
      LAYER via ;
        RECT 2588.520 1687.800 2588.780 1688.060 ;
        RECT 2594.040 1687.800 2594.300 1688.060 ;
        RECT 2594.040 20.440 2594.300 20.700 ;
        RECT 2797.820 20.440 2798.080 20.700 ;
      LAYER met2 ;
        RECT 2588.440 1700.000 2588.720 1702.400 ;
        RECT 2588.580 1688.090 2588.720 1700.000 ;
        RECT 2588.520 1687.770 2588.780 1688.090 ;
        RECT 2594.040 1687.770 2594.300 1688.090 ;
        RECT 2594.100 20.730 2594.240 1687.770 ;
        RECT 2594.040 20.410 2594.300 20.730 ;
        RECT 2797.820 20.410 2798.080 20.730 ;
        RECT 2797.880 2.400 2798.020 20.410 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2620.305 1685.805 2620.475 1687.335 ;
        RECT 2633.645 1685.805 2633.815 1688.015 ;
      LAYER mcon ;
        RECT 2633.645 1687.845 2633.815 1688.015 ;
        RECT 2620.305 1687.165 2620.475 1687.335 ;
      LAYER met1 ;
        RECT 2633.585 1688.000 2633.875 1688.045 ;
        RECT 2815.730 1688.000 2816.050 1688.060 ;
        RECT 2633.585 1687.860 2816.050 1688.000 ;
        RECT 2633.585 1687.815 2633.875 1687.860 ;
        RECT 2815.730 1687.800 2816.050 1687.860 ;
        RECT 2597.690 1687.320 2598.010 1687.380 ;
        RECT 2620.245 1687.320 2620.535 1687.365 ;
        RECT 2597.690 1687.180 2620.535 1687.320 ;
        RECT 2597.690 1687.120 2598.010 1687.180 ;
        RECT 2620.245 1687.135 2620.535 1687.180 ;
        RECT 2620.245 1685.960 2620.535 1686.005 ;
        RECT 2633.585 1685.960 2633.875 1686.005 ;
        RECT 2620.245 1685.820 2633.875 1685.960 ;
        RECT 2620.245 1685.775 2620.535 1685.820 ;
        RECT 2633.585 1685.775 2633.875 1685.820 ;
      LAYER via ;
        RECT 2815.760 1687.800 2816.020 1688.060 ;
        RECT 2597.720 1687.120 2597.980 1687.380 ;
      LAYER met2 ;
        RECT 2597.640 1700.000 2597.920 1702.400 ;
        RECT 2597.780 1687.410 2597.920 1700.000 ;
        RECT 2815.760 1687.770 2816.020 1688.090 ;
        RECT 2597.720 1687.090 2597.980 1687.410 ;
        RECT 2815.820 2.400 2815.960 1687.770 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2607.810 19.620 2608.130 19.680 ;
        RECT 2833.670 19.620 2833.990 19.680 ;
        RECT 2607.810 19.480 2833.990 19.620 ;
        RECT 2607.810 19.420 2608.130 19.480 ;
        RECT 2833.670 19.420 2833.990 19.480 ;
      LAYER via ;
        RECT 2607.840 19.420 2608.100 19.680 ;
        RECT 2833.700 19.420 2833.960 19.680 ;
      LAYER met2 ;
        RECT 2606.840 1700.410 2607.120 1702.400 ;
        RECT 2606.840 1700.270 2608.040 1700.410 ;
        RECT 2606.840 1700.000 2607.120 1700.270 ;
        RECT 2607.900 19.710 2608.040 1700.270 ;
        RECT 2607.840 19.390 2608.100 19.710 ;
        RECT 2833.700 19.390 2833.960 19.710 ;
        RECT 2833.760 2.400 2833.900 19.390 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2846.090 1687.320 2846.410 1687.380 ;
        RECT 2634.120 1687.180 2846.410 1687.320 ;
        RECT 2616.090 1686.980 2616.410 1687.040 ;
        RECT 2634.120 1686.980 2634.260 1687.180 ;
        RECT 2846.090 1687.120 2846.410 1687.180 ;
        RECT 2616.090 1686.840 2634.260 1686.980 ;
        RECT 2616.090 1686.780 2616.410 1686.840 ;
        RECT 2846.090 16.900 2846.410 16.960 ;
        RECT 2851.150 16.900 2851.470 16.960 ;
        RECT 2846.090 16.760 2851.470 16.900 ;
        RECT 2846.090 16.700 2846.410 16.760 ;
        RECT 2851.150 16.700 2851.470 16.760 ;
      LAYER via ;
        RECT 2616.120 1686.780 2616.380 1687.040 ;
        RECT 2846.120 1687.120 2846.380 1687.380 ;
        RECT 2846.120 16.700 2846.380 16.960 ;
        RECT 2851.180 16.700 2851.440 16.960 ;
      LAYER met2 ;
        RECT 2616.040 1700.000 2616.320 1702.400 ;
        RECT 2616.180 1687.070 2616.320 1700.000 ;
        RECT 2846.120 1687.090 2846.380 1687.410 ;
        RECT 2616.120 1686.750 2616.380 1687.070 ;
        RECT 2846.180 16.990 2846.320 1687.090 ;
        RECT 2846.120 16.670 2846.380 16.990 ;
        RECT 2851.180 16.670 2851.440 16.990 ;
        RECT 2851.240 2.400 2851.380 16.670 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2627.590 18.260 2627.910 18.320 ;
        RECT 2869.090 18.260 2869.410 18.320 ;
        RECT 2627.590 18.120 2869.410 18.260 ;
        RECT 2627.590 18.060 2627.910 18.120 ;
        RECT 2869.090 18.060 2869.410 18.120 ;
      LAYER via ;
        RECT 2627.620 18.060 2627.880 18.320 ;
        RECT 2869.120 18.060 2869.380 18.320 ;
      LAYER met2 ;
        RECT 2625.240 1700.410 2625.520 1702.400 ;
        RECT 2625.240 1700.270 2627.820 1700.410 ;
        RECT 2625.240 1700.000 2625.520 1700.270 ;
        RECT 2627.680 18.350 2627.820 1700.270 ;
        RECT 2627.620 18.030 2627.880 18.350 ;
        RECT 2869.120 18.030 2869.380 18.350 ;
        RECT 2869.180 2.400 2869.320 18.030 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2634.490 1686.980 2634.810 1687.040 ;
        RECT 2859.890 1686.980 2860.210 1687.040 ;
        RECT 2634.490 1686.840 2860.210 1686.980 ;
        RECT 2634.490 1686.780 2634.810 1686.840 ;
        RECT 2859.890 1686.780 2860.210 1686.840 ;
        RECT 2859.890 15.200 2860.210 15.260 ;
        RECT 2887.030 15.200 2887.350 15.260 ;
        RECT 2859.890 15.060 2887.350 15.200 ;
        RECT 2859.890 15.000 2860.210 15.060 ;
        RECT 2887.030 15.000 2887.350 15.060 ;
      LAYER via ;
        RECT 2634.520 1686.780 2634.780 1687.040 ;
        RECT 2859.920 1686.780 2860.180 1687.040 ;
        RECT 2859.920 15.000 2860.180 15.260 ;
        RECT 2887.060 15.000 2887.320 15.260 ;
      LAYER met2 ;
        RECT 2634.440 1700.000 2634.720 1702.400 ;
        RECT 2634.580 1687.070 2634.720 1700.000 ;
        RECT 2634.520 1686.750 2634.780 1687.070 ;
        RECT 2859.920 1686.750 2860.180 1687.070 ;
        RECT 2859.980 15.290 2860.120 1686.750 ;
        RECT 2859.920 14.970 2860.180 15.290 ;
        RECT 2887.060 14.970 2887.320 15.290 ;
        RECT 2887.120 2.400 2887.260 14.970 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2643.690 1685.960 2644.010 1686.020 ;
        RECT 2648.750 1685.960 2649.070 1686.020 ;
        RECT 2643.690 1685.820 2649.070 1685.960 ;
        RECT 2643.690 1685.760 2644.010 1685.820 ;
        RECT 2648.750 1685.760 2649.070 1685.820 ;
        RECT 2648.750 17.240 2649.070 17.300 ;
        RECT 2904.970 17.240 2905.290 17.300 ;
        RECT 2648.750 17.100 2905.290 17.240 ;
        RECT 2648.750 17.040 2649.070 17.100 ;
        RECT 2904.970 17.040 2905.290 17.100 ;
      LAYER via ;
        RECT 2643.720 1685.760 2643.980 1686.020 ;
        RECT 2648.780 1685.760 2649.040 1686.020 ;
        RECT 2648.780 17.040 2649.040 17.300 ;
        RECT 2905.000 17.040 2905.260 17.300 ;
      LAYER met2 ;
        RECT 2643.640 1700.000 2643.920 1702.400 ;
        RECT 2643.780 1686.050 2643.920 1700.000 ;
        RECT 2643.720 1685.730 2643.980 1686.050 ;
        RECT 2648.780 1685.730 2649.040 1686.050 ;
        RECT 2648.840 17.330 2648.980 1685.730 ;
        RECT 2648.780 17.010 2649.040 17.330 ;
        RECT 2905.000 17.010 2905.260 17.330 ;
        RECT 2905.060 2.400 2905.200 17.010 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 852.910 30.160 853.230 30.220 ;
        RECT 1587.070 30.160 1587.390 30.220 ;
        RECT 852.910 30.020 1587.390 30.160 ;
        RECT 852.910 29.960 853.230 30.020 ;
        RECT 1587.070 29.960 1587.390 30.020 ;
      LAYER via ;
        RECT 852.940 29.960 853.200 30.220 ;
        RECT 1587.100 29.960 1587.360 30.220 ;
      LAYER met2 ;
        RECT 1587.480 1700.410 1587.760 1702.400 ;
        RECT 1587.160 1700.270 1587.760 1700.410 ;
        RECT 1587.160 30.250 1587.300 1700.270 ;
        RECT 1587.480 1700.000 1587.760 1700.270 ;
        RECT 852.940 29.930 853.200 30.250 ;
        RECT 1587.100 29.930 1587.360 30.250 ;
        RECT 853.000 2.400 853.140 29.930 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 29.820 871.170 29.880 ;
        RECT 870.850 29.680 1576.720 29.820 ;
        RECT 870.850 29.620 871.170 29.680 ;
        RECT 1576.580 29.480 1576.720 29.680 ;
        RECT 1594.430 29.480 1594.750 29.540 ;
        RECT 1576.580 29.340 1594.750 29.480 ;
        RECT 1594.430 29.280 1594.750 29.340 ;
      LAYER via ;
        RECT 870.880 29.620 871.140 29.880 ;
        RECT 1594.460 29.280 1594.720 29.540 ;
      LAYER met2 ;
        RECT 1596.680 1700.410 1596.960 1702.400 ;
        RECT 1594.060 1700.270 1596.960 1700.410 ;
        RECT 1594.060 34.410 1594.200 1700.270 ;
        RECT 1596.680 1700.000 1596.960 1700.270 ;
        RECT 1594.060 34.270 1594.660 34.410 ;
        RECT 870.880 29.590 871.140 29.910 ;
        RECT 870.940 2.400 871.080 29.590 ;
        RECT 1594.520 29.570 1594.660 34.270 ;
        RECT 1594.460 29.250 1594.720 29.570 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1576.105 29.325 1576.275 33.915 ;
      LAYER mcon ;
        RECT 1576.105 33.745 1576.275 33.915 ;
      LAYER met1 ;
        RECT 1600.870 1689.700 1601.190 1689.760 ;
        RECT 1604.550 1689.700 1604.870 1689.760 ;
        RECT 1600.870 1689.560 1604.870 1689.700 ;
        RECT 1600.870 1689.500 1601.190 1689.560 ;
        RECT 1604.550 1689.500 1604.870 1689.560 ;
        RECT 1576.045 33.900 1576.335 33.945 ;
        RECT 1600.870 33.900 1601.190 33.960 ;
        RECT 1576.045 33.760 1601.190 33.900 ;
        RECT 1576.045 33.715 1576.335 33.760 ;
        RECT 1600.870 33.700 1601.190 33.760 ;
        RECT 888.790 29.480 889.110 29.540 ;
        RECT 1576.045 29.480 1576.335 29.525 ;
        RECT 888.790 29.340 1576.335 29.480 ;
        RECT 888.790 29.280 889.110 29.340 ;
        RECT 1576.045 29.295 1576.335 29.340 ;
      LAYER via ;
        RECT 1600.900 1689.500 1601.160 1689.760 ;
        RECT 1604.580 1689.500 1604.840 1689.760 ;
        RECT 1600.900 33.700 1601.160 33.960 ;
        RECT 888.820 29.280 889.080 29.540 ;
      LAYER met2 ;
        RECT 1605.880 1700.410 1606.160 1702.400 ;
        RECT 1604.640 1700.270 1606.160 1700.410 ;
        RECT 1604.640 1689.790 1604.780 1700.270 ;
        RECT 1605.880 1700.000 1606.160 1700.270 ;
        RECT 1600.900 1689.470 1601.160 1689.790 ;
        RECT 1604.580 1689.470 1604.840 1689.790 ;
        RECT 1600.960 33.990 1601.100 1689.470 ;
        RECT 1600.900 33.670 1601.160 33.990 ;
        RECT 888.820 29.250 889.080 29.570 ;
        RECT 888.880 2.400 889.020 29.250 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1611.065 28.985 1611.235 30.175 ;
      LAYER mcon ;
        RECT 1611.065 30.005 1611.235 30.175 ;
      LAYER met1 ;
        RECT 1611.005 30.160 1611.295 30.205 ;
        RECT 1614.670 30.160 1614.990 30.220 ;
        RECT 1611.005 30.020 1614.990 30.160 ;
        RECT 1611.005 29.975 1611.295 30.020 ;
        RECT 1614.670 29.960 1614.990 30.020 ;
        RECT 906.730 29.140 907.050 29.200 ;
        RECT 1611.005 29.140 1611.295 29.185 ;
        RECT 906.730 29.000 1611.295 29.140 ;
        RECT 906.730 28.940 907.050 29.000 ;
        RECT 1611.005 28.955 1611.295 29.000 ;
      LAYER via ;
        RECT 1614.700 29.960 1614.960 30.220 ;
        RECT 906.760 28.940 907.020 29.200 ;
      LAYER met2 ;
        RECT 1615.080 1700.410 1615.360 1702.400 ;
        RECT 1614.760 1700.270 1615.360 1700.410 ;
        RECT 1614.760 30.250 1614.900 1700.270 ;
        RECT 1615.080 1700.000 1615.360 1700.270 ;
        RECT 1614.700 29.930 1614.960 30.250 ;
        RECT 906.760 28.910 907.020 29.230 ;
        RECT 906.820 2.400 906.960 28.910 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 28.800 924.530 28.860 ;
        RECT 1621.570 28.800 1621.890 28.860 ;
        RECT 924.210 28.660 1621.890 28.800 ;
        RECT 924.210 28.600 924.530 28.660 ;
        RECT 1621.570 28.600 1621.890 28.660 ;
      LAYER via ;
        RECT 924.240 28.600 924.500 28.860 ;
        RECT 1621.600 28.600 1621.860 28.860 ;
      LAYER met2 ;
        RECT 1624.280 1700.410 1624.560 1702.400 ;
        RECT 1621.660 1700.270 1624.560 1700.410 ;
        RECT 1621.660 28.890 1621.800 1700.270 ;
        RECT 1624.280 1700.000 1624.560 1700.270 ;
        RECT 924.240 28.570 924.500 28.890 ;
        RECT 1621.600 28.570 1621.860 28.890 ;
        RECT 924.300 2.400 924.440 28.570 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1628.470 1663.860 1628.790 1663.920 ;
        RECT 1632.150 1663.860 1632.470 1663.920 ;
        RECT 1628.470 1663.720 1632.470 1663.860 ;
        RECT 1628.470 1663.660 1628.790 1663.720 ;
        RECT 1632.150 1663.660 1632.470 1663.720 ;
        RECT 942.150 28.460 942.470 28.520 ;
        RECT 1628.470 28.460 1628.790 28.520 ;
        RECT 942.150 28.320 1628.790 28.460 ;
        RECT 942.150 28.260 942.470 28.320 ;
        RECT 1628.470 28.260 1628.790 28.320 ;
      LAYER via ;
        RECT 1628.500 1663.660 1628.760 1663.920 ;
        RECT 1632.180 1663.660 1632.440 1663.920 ;
        RECT 942.180 28.260 942.440 28.520 ;
        RECT 1628.500 28.260 1628.760 28.520 ;
      LAYER met2 ;
        RECT 1633.480 1700.410 1633.760 1702.400 ;
        RECT 1632.240 1700.270 1633.760 1700.410 ;
        RECT 1632.240 1663.950 1632.380 1700.270 ;
        RECT 1633.480 1700.000 1633.760 1700.270 ;
        RECT 1628.500 1663.630 1628.760 1663.950 ;
        RECT 1632.180 1663.630 1632.440 1663.950 ;
        RECT 1628.560 28.550 1628.700 1663.630 ;
        RECT 942.180 28.230 942.440 28.550 ;
        RECT 1628.500 28.230 1628.760 28.550 ;
        RECT 942.240 2.400 942.380 28.230 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 960.090 28.120 960.410 28.180 ;
        RECT 1642.270 28.120 1642.590 28.180 ;
        RECT 960.090 27.980 1642.590 28.120 ;
        RECT 960.090 27.920 960.410 27.980 ;
        RECT 1642.270 27.920 1642.590 27.980 ;
      LAYER via ;
        RECT 960.120 27.920 960.380 28.180 ;
        RECT 1642.300 27.920 1642.560 28.180 ;
      LAYER met2 ;
        RECT 1642.680 1700.410 1642.960 1702.400 ;
        RECT 1642.360 1700.270 1642.960 1700.410 ;
        RECT 1642.360 28.210 1642.500 1700.270 ;
        RECT 1642.680 1700.000 1642.960 1700.270 ;
        RECT 960.120 27.890 960.380 28.210 ;
        RECT 1642.300 27.890 1642.560 28.210 ;
        RECT 960.180 2.400 960.320 27.890 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 978.030 27.780 978.350 27.840 ;
        RECT 1649.170 27.780 1649.490 27.840 ;
        RECT 978.030 27.640 1649.490 27.780 ;
        RECT 978.030 27.580 978.350 27.640 ;
        RECT 1649.170 27.580 1649.490 27.640 ;
      LAYER via ;
        RECT 978.060 27.580 978.320 27.840 ;
        RECT 1649.200 27.580 1649.460 27.840 ;
      LAYER met2 ;
        RECT 1651.880 1700.410 1652.160 1702.400 ;
        RECT 1649.260 1700.270 1652.160 1700.410 ;
        RECT 1649.260 27.870 1649.400 1700.270 ;
        RECT 1651.880 1700.000 1652.160 1700.270 ;
        RECT 978.060 27.550 978.320 27.870 ;
        RECT 1649.200 27.550 1649.460 27.870 ;
        RECT 978.120 2.400 978.260 27.550 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 65.860 662.330 65.920 ;
        RECT 1484.490 65.860 1484.810 65.920 ;
        RECT 662.010 65.720 1484.810 65.860 ;
        RECT 662.010 65.660 662.330 65.720 ;
        RECT 1484.490 65.660 1484.810 65.720 ;
      LAYER via ;
        RECT 662.040 65.660 662.300 65.920 ;
        RECT 1484.520 65.660 1484.780 65.920 ;
      LAYER met2 ;
        RECT 1486.740 1700.410 1487.020 1702.400 ;
        RECT 1484.580 1700.270 1487.020 1700.410 ;
        RECT 1484.580 65.950 1484.720 1700.270 ;
        RECT 1486.740 1700.000 1487.020 1700.270 ;
        RECT 662.040 65.630 662.300 65.950 ;
        RECT 1484.520 65.630 1484.780 65.950 ;
        RECT 662.100 17.410 662.240 65.630 ;
        RECT 657.040 17.270 662.240 17.410 ;
        RECT 657.040 2.400 657.180 17.270 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1657.065 1442.025 1657.235 1490.475 ;
        RECT 1657.065 1007.505 1657.235 1014.815 ;
        RECT 1657.065 758.965 1657.235 807.075 ;
        RECT 1657.065 386.325 1657.235 434.435 ;
        RECT 1657.065 241.485 1657.235 278.375 ;
      LAYER mcon ;
        RECT 1657.065 1490.305 1657.235 1490.475 ;
        RECT 1657.065 1014.645 1657.235 1014.815 ;
        RECT 1657.065 806.905 1657.235 807.075 ;
        RECT 1657.065 434.265 1657.235 434.435 ;
        RECT 1657.065 278.205 1657.235 278.375 ;
      LAYER met1 ;
        RECT 1657.450 1642.440 1657.770 1642.500 ;
        RECT 1658.370 1642.440 1658.690 1642.500 ;
        RECT 1657.450 1642.300 1658.690 1642.440 ;
        RECT 1657.450 1642.240 1657.770 1642.300 ;
        RECT 1658.370 1642.240 1658.690 1642.300 ;
        RECT 1656.990 1497.260 1657.310 1497.320 ;
        RECT 1657.450 1497.260 1657.770 1497.320 ;
        RECT 1656.990 1497.120 1657.770 1497.260 ;
        RECT 1656.990 1497.060 1657.310 1497.120 ;
        RECT 1657.450 1497.060 1657.770 1497.120 ;
        RECT 1656.990 1490.460 1657.310 1490.520 ;
        RECT 1656.795 1490.320 1657.310 1490.460 ;
        RECT 1656.990 1490.260 1657.310 1490.320 ;
        RECT 1656.990 1442.180 1657.310 1442.240 ;
        RECT 1656.795 1442.040 1657.310 1442.180 ;
        RECT 1656.990 1441.980 1657.310 1442.040 ;
        RECT 1656.990 1414.440 1657.310 1414.700 ;
        RECT 1657.080 1413.960 1657.220 1414.440 ;
        RECT 1657.450 1413.960 1657.770 1414.020 ;
        RECT 1657.080 1413.820 1657.770 1413.960 ;
        RECT 1657.450 1413.760 1657.770 1413.820 ;
        RECT 1655.610 1400.700 1655.930 1400.760 ;
        RECT 1657.450 1400.700 1657.770 1400.760 ;
        RECT 1655.610 1400.560 1657.770 1400.700 ;
        RECT 1655.610 1400.500 1655.930 1400.560 ;
        RECT 1657.450 1400.500 1657.770 1400.560 ;
        RECT 1656.530 1317.740 1656.850 1317.800 ;
        RECT 1656.530 1317.600 1657.680 1317.740 ;
        RECT 1656.530 1317.540 1656.850 1317.600 ;
        RECT 1657.540 1317.460 1657.680 1317.600 ;
        RECT 1657.450 1317.200 1657.770 1317.460 ;
        RECT 1655.610 1304.140 1655.930 1304.200 ;
        RECT 1657.450 1304.140 1657.770 1304.200 ;
        RECT 1655.610 1304.000 1657.770 1304.140 ;
        RECT 1655.610 1303.940 1655.930 1304.000 ;
        RECT 1657.450 1303.940 1657.770 1304.000 ;
        RECT 1655.610 1207.580 1655.930 1207.640 ;
        RECT 1657.450 1207.580 1657.770 1207.640 ;
        RECT 1655.610 1207.440 1657.770 1207.580 ;
        RECT 1655.610 1207.380 1655.930 1207.440 ;
        RECT 1657.450 1207.380 1657.770 1207.440 ;
        RECT 1657.450 1159.100 1657.770 1159.360 ;
        RECT 1657.540 1158.680 1657.680 1159.100 ;
        RECT 1657.450 1158.420 1657.770 1158.680 ;
        RECT 1656.530 1104.220 1656.850 1104.280 ;
        RECT 1657.910 1104.220 1658.230 1104.280 ;
        RECT 1656.530 1104.080 1658.230 1104.220 ;
        RECT 1656.530 1104.020 1656.850 1104.080 ;
        RECT 1657.910 1104.020 1658.230 1104.080 ;
        RECT 1655.610 1097.080 1655.930 1097.140 ;
        RECT 1656.530 1097.080 1656.850 1097.140 ;
        RECT 1655.610 1096.940 1656.850 1097.080 ;
        RECT 1655.610 1096.880 1655.930 1096.940 ;
        RECT 1656.530 1096.880 1656.850 1096.940 ;
        RECT 1657.005 1014.800 1657.295 1014.845 ;
        RECT 1657.450 1014.800 1657.770 1014.860 ;
        RECT 1657.005 1014.660 1657.770 1014.800 ;
        RECT 1657.005 1014.615 1657.295 1014.660 ;
        RECT 1657.450 1014.600 1657.770 1014.660 ;
        RECT 1656.990 1007.660 1657.310 1007.720 ;
        RECT 1656.795 1007.520 1657.310 1007.660 ;
        RECT 1656.990 1007.460 1657.310 1007.520 ;
        RECT 1655.150 983.180 1655.470 983.240 ;
        RECT 1656.990 983.180 1657.310 983.240 ;
        RECT 1655.150 983.040 1657.310 983.180 ;
        RECT 1655.150 982.980 1655.470 983.040 ;
        RECT 1656.990 982.980 1657.310 983.040 ;
        RECT 1655.610 917.900 1655.930 917.960 ;
        RECT 1657.450 917.900 1657.770 917.960 ;
        RECT 1655.610 917.760 1657.770 917.900 ;
        RECT 1655.610 917.700 1655.930 917.760 ;
        RECT 1657.450 917.700 1657.770 917.760 ;
        RECT 1656.990 807.060 1657.310 807.120 ;
        RECT 1656.795 806.920 1657.310 807.060 ;
        RECT 1656.990 806.860 1657.310 806.920 ;
        RECT 1656.990 759.120 1657.310 759.180 ;
        RECT 1656.795 758.980 1657.310 759.120 ;
        RECT 1656.990 758.920 1657.310 758.980 ;
        RECT 1656.990 738.520 1657.310 738.780 ;
        RECT 1657.080 738.100 1657.220 738.520 ;
        RECT 1656.990 737.840 1657.310 738.100 ;
        RECT 1656.990 531.320 1657.310 531.380 ;
        RECT 1657.450 531.320 1657.770 531.380 ;
        RECT 1656.990 531.180 1657.770 531.320 ;
        RECT 1656.990 531.120 1657.310 531.180 ;
        RECT 1657.450 531.120 1657.770 531.180 ;
        RECT 1656.990 434.420 1657.310 434.480 ;
        RECT 1656.795 434.280 1657.310 434.420 ;
        RECT 1656.990 434.220 1657.310 434.280 ;
        RECT 1656.990 386.480 1657.310 386.540 ;
        RECT 1656.795 386.340 1657.310 386.480 ;
        RECT 1656.990 386.280 1657.310 386.340 ;
        RECT 1656.990 278.360 1657.310 278.420 ;
        RECT 1656.795 278.220 1657.310 278.360 ;
        RECT 1656.990 278.160 1657.310 278.220 ;
        RECT 1657.005 241.640 1657.295 241.685 ;
        RECT 1657.450 241.640 1657.770 241.700 ;
        RECT 1657.005 241.500 1657.770 241.640 ;
        RECT 1657.005 241.455 1657.295 241.500 ;
        RECT 1657.450 241.440 1657.770 241.500 ;
        RECT 1657.450 186.900 1657.770 186.960 ;
        RECT 1657.080 186.760 1657.770 186.900 ;
        RECT 1657.080 186.620 1657.220 186.760 ;
        RECT 1657.450 186.700 1657.770 186.760 ;
        RECT 1656.990 186.360 1657.310 186.620 ;
        RECT 1000.110 65.180 1000.430 65.240 ;
        RECT 1656.990 65.180 1657.310 65.240 ;
        RECT 1000.110 65.040 1657.310 65.180 ;
        RECT 1000.110 64.980 1000.430 65.040 ;
        RECT 1656.990 64.980 1657.310 65.040 ;
      LAYER via ;
        RECT 1657.480 1642.240 1657.740 1642.500 ;
        RECT 1658.400 1642.240 1658.660 1642.500 ;
        RECT 1657.020 1497.060 1657.280 1497.320 ;
        RECT 1657.480 1497.060 1657.740 1497.320 ;
        RECT 1657.020 1490.260 1657.280 1490.520 ;
        RECT 1657.020 1441.980 1657.280 1442.240 ;
        RECT 1657.020 1414.440 1657.280 1414.700 ;
        RECT 1657.480 1413.760 1657.740 1414.020 ;
        RECT 1655.640 1400.500 1655.900 1400.760 ;
        RECT 1657.480 1400.500 1657.740 1400.760 ;
        RECT 1656.560 1317.540 1656.820 1317.800 ;
        RECT 1657.480 1317.200 1657.740 1317.460 ;
        RECT 1655.640 1303.940 1655.900 1304.200 ;
        RECT 1657.480 1303.940 1657.740 1304.200 ;
        RECT 1655.640 1207.380 1655.900 1207.640 ;
        RECT 1657.480 1207.380 1657.740 1207.640 ;
        RECT 1657.480 1159.100 1657.740 1159.360 ;
        RECT 1657.480 1158.420 1657.740 1158.680 ;
        RECT 1656.560 1104.020 1656.820 1104.280 ;
        RECT 1657.940 1104.020 1658.200 1104.280 ;
        RECT 1655.640 1096.880 1655.900 1097.140 ;
        RECT 1656.560 1096.880 1656.820 1097.140 ;
        RECT 1657.480 1014.600 1657.740 1014.860 ;
        RECT 1657.020 1007.460 1657.280 1007.720 ;
        RECT 1655.180 982.980 1655.440 983.240 ;
        RECT 1657.020 982.980 1657.280 983.240 ;
        RECT 1655.640 917.700 1655.900 917.960 ;
        RECT 1657.480 917.700 1657.740 917.960 ;
        RECT 1657.020 806.860 1657.280 807.120 ;
        RECT 1657.020 758.920 1657.280 759.180 ;
        RECT 1657.020 738.520 1657.280 738.780 ;
        RECT 1657.020 737.840 1657.280 738.100 ;
        RECT 1657.020 531.120 1657.280 531.380 ;
        RECT 1657.480 531.120 1657.740 531.380 ;
        RECT 1657.020 434.220 1657.280 434.480 ;
        RECT 1657.020 386.280 1657.280 386.540 ;
        RECT 1657.020 278.160 1657.280 278.420 ;
        RECT 1657.480 241.440 1657.740 241.700 ;
        RECT 1657.480 186.700 1657.740 186.960 ;
        RECT 1657.020 186.360 1657.280 186.620 ;
        RECT 1000.140 64.980 1000.400 65.240 ;
        RECT 1657.020 64.980 1657.280 65.240 ;
      LAYER met2 ;
        RECT 1661.080 1701.090 1661.360 1702.400 ;
        RECT 1658.460 1700.950 1661.360 1701.090 ;
        RECT 1658.460 1642.530 1658.600 1700.950 ;
        RECT 1661.080 1700.000 1661.360 1700.950 ;
        RECT 1657.480 1642.210 1657.740 1642.530 ;
        RECT 1658.400 1642.210 1658.660 1642.530 ;
        RECT 1657.540 1546.050 1657.680 1642.210 ;
        RECT 1657.080 1545.910 1657.680 1546.050 ;
        RECT 1657.080 1510.010 1657.220 1545.910 ;
        RECT 1657.080 1509.870 1657.680 1510.010 ;
        RECT 1657.540 1497.350 1657.680 1509.870 ;
        RECT 1657.020 1497.030 1657.280 1497.350 ;
        RECT 1657.480 1497.030 1657.740 1497.350 ;
        RECT 1657.080 1490.550 1657.220 1497.030 ;
        RECT 1657.020 1490.230 1657.280 1490.550 ;
        RECT 1657.020 1441.950 1657.280 1442.270 ;
        RECT 1657.080 1414.730 1657.220 1441.950 ;
        RECT 1657.020 1414.410 1657.280 1414.730 ;
        RECT 1657.480 1413.730 1657.740 1414.050 ;
        RECT 1657.540 1400.790 1657.680 1413.730 ;
        RECT 1655.640 1400.470 1655.900 1400.790 ;
        RECT 1657.480 1400.470 1657.740 1400.790 ;
        RECT 1655.700 1353.045 1655.840 1400.470 ;
        RECT 1655.630 1352.675 1655.910 1353.045 ;
        RECT 1656.550 1351.995 1656.830 1352.365 ;
        RECT 1656.620 1317.830 1656.760 1351.995 ;
        RECT 1656.560 1317.510 1656.820 1317.830 ;
        RECT 1657.480 1317.170 1657.740 1317.490 ;
        RECT 1657.540 1304.230 1657.680 1317.170 ;
        RECT 1655.640 1303.910 1655.900 1304.230 ;
        RECT 1657.480 1303.910 1657.740 1304.230 ;
        RECT 1655.700 1256.485 1655.840 1303.910 ;
        RECT 1655.630 1256.115 1655.910 1256.485 ;
        RECT 1655.630 1255.435 1655.910 1255.805 ;
        RECT 1655.700 1207.670 1655.840 1255.435 ;
        RECT 1655.640 1207.350 1655.900 1207.670 ;
        RECT 1657.480 1207.350 1657.740 1207.670 ;
        RECT 1657.540 1159.390 1657.680 1207.350 ;
        RECT 1657.480 1159.070 1657.740 1159.390 ;
        RECT 1657.480 1158.390 1657.740 1158.710 ;
        RECT 1657.540 1111.530 1657.680 1158.390 ;
        RECT 1657.540 1111.390 1658.140 1111.530 ;
        RECT 1658.000 1104.310 1658.140 1111.390 ;
        RECT 1656.560 1103.990 1656.820 1104.310 ;
        RECT 1657.940 1103.990 1658.200 1104.310 ;
        RECT 1656.620 1097.170 1656.760 1103.990 ;
        RECT 1655.640 1096.850 1655.900 1097.170 ;
        RECT 1656.560 1096.850 1656.820 1097.170 ;
        RECT 1655.700 1049.085 1655.840 1096.850 ;
        RECT 1655.630 1048.715 1655.910 1049.085 ;
        RECT 1657.470 1048.715 1657.750 1049.085 ;
        RECT 1657.540 1014.890 1657.680 1048.715 ;
        RECT 1657.480 1014.570 1657.740 1014.890 ;
        RECT 1657.020 1007.430 1657.280 1007.750 ;
        RECT 1657.080 983.270 1657.220 1007.430 ;
        RECT 1655.180 982.950 1655.440 983.270 ;
        RECT 1657.020 982.950 1657.280 983.270 ;
        RECT 1655.240 966.010 1655.380 982.950 ;
        RECT 1655.240 965.870 1655.840 966.010 ;
        RECT 1655.700 917.990 1655.840 965.870 ;
        RECT 1655.640 917.670 1655.900 917.990 ;
        RECT 1657.480 917.670 1657.740 917.990 ;
        RECT 1657.540 863.445 1657.680 917.670 ;
        RECT 1657.470 863.075 1657.750 863.445 ;
        RECT 1657.010 862.395 1657.290 862.765 ;
        RECT 1657.080 807.150 1657.220 862.395 ;
        RECT 1657.020 806.830 1657.280 807.150 ;
        RECT 1657.020 758.890 1657.280 759.210 ;
        RECT 1657.080 738.810 1657.220 758.890 ;
        RECT 1657.020 738.490 1657.280 738.810 ;
        RECT 1657.020 737.810 1657.280 738.130 ;
        RECT 1657.080 724.610 1657.220 737.810 ;
        RECT 1657.080 724.470 1657.680 724.610 ;
        RECT 1657.540 676.330 1657.680 724.470 ;
        RECT 1657.080 676.190 1657.680 676.330 ;
        RECT 1657.080 628.050 1657.220 676.190 ;
        RECT 1657.080 627.910 1657.680 628.050 ;
        RECT 1657.540 594.730 1657.680 627.910 ;
        RECT 1657.540 594.590 1658.140 594.730 ;
        RECT 1658.000 593.370 1658.140 594.590 ;
        RECT 1657.540 593.230 1658.140 593.370 ;
        RECT 1657.540 531.410 1657.680 593.230 ;
        RECT 1657.020 531.090 1657.280 531.410 ;
        RECT 1657.480 531.090 1657.740 531.410 ;
        RECT 1657.080 434.510 1657.220 531.090 ;
        RECT 1657.020 434.190 1657.280 434.510 ;
        RECT 1657.020 386.250 1657.280 386.570 ;
        RECT 1657.080 278.450 1657.220 386.250 ;
        RECT 1657.020 278.130 1657.280 278.450 ;
        RECT 1657.480 241.410 1657.740 241.730 ;
        RECT 1657.540 186.990 1657.680 241.410 ;
        RECT 1657.480 186.670 1657.740 186.990 ;
        RECT 1657.020 186.330 1657.280 186.650 ;
        RECT 1657.080 65.270 1657.220 186.330 ;
        RECT 1000.140 64.950 1000.400 65.270 ;
        RECT 1657.020 64.950 1657.280 65.270 ;
        RECT 1000.200 17.410 1000.340 64.950 ;
        RECT 996.060 17.270 1000.340 17.410 ;
        RECT 996.060 2.400 996.200 17.270 ;
        RECT 995.850 -4.800 996.410 2.400 ;
      LAYER via2 ;
        RECT 1655.630 1352.720 1655.910 1353.000 ;
        RECT 1656.550 1352.040 1656.830 1352.320 ;
        RECT 1655.630 1256.160 1655.910 1256.440 ;
        RECT 1655.630 1255.480 1655.910 1255.760 ;
        RECT 1655.630 1048.760 1655.910 1049.040 ;
        RECT 1657.470 1048.760 1657.750 1049.040 ;
        RECT 1657.470 863.120 1657.750 863.400 ;
        RECT 1657.010 862.440 1657.290 862.720 ;
      LAYER met3 ;
        RECT 1655.605 1353.010 1655.935 1353.025 ;
        RECT 1655.605 1352.710 1656.610 1353.010 ;
        RECT 1655.605 1352.695 1655.935 1352.710 ;
        RECT 1656.310 1352.345 1656.610 1352.710 ;
        RECT 1656.310 1352.030 1656.855 1352.345 ;
        RECT 1656.525 1352.015 1656.855 1352.030 ;
        RECT 1655.605 1256.450 1655.935 1256.465 ;
        RECT 1655.605 1256.150 1656.610 1256.450 ;
        RECT 1655.605 1256.135 1655.935 1256.150 ;
        RECT 1655.605 1255.770 1655.935 1255.785 ;
        RECT 1656.310 1255.770 1656.610 1256.150 ;
        RECT 1655.605 1255.470 1656.610 1255.770 ;
        RECT 1655.605 1255.455 1655.935 1255.470 ;
        RECT 1655.605 1049.050 1655.935 1049.065 ;
        RECT 1657.445 1049.050 1657.775 1049.065 ;
        RECT 1655.605 1048.750 1657.775 1049.050 ;
        RECT 1655.605 1048.735 1655.935 1048.750 ;
        RECT 1657.445 1048.735 1657.775 1048.750 ;
        RECT 1657.445 863.410 1657.775 863.425 ;
        RECT 1656.310 863.110 1657.775 863.410 ;
        RECT 1656.310 862.730 1656.610 863.110 ;
        RECT 1657.445 863.095 1657.775 863.110 ;
        RECT 1656.985 862.730 1657.315 862.745 ;
        RECT 1656.310 862.430 1657.315 862.730 ;
        RECT 1656.985 862.415 1657.315 862.430 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1670.330 1677.120 1670.650 1677.180 ;
        RECT 1670.330 1676.980 1671.020 1677.120 ;
        RECT 1670.330 1676.920 1670.650 1676.980 ;
        RECT 1670.880 1676.160 1671.020 1676.980 ;
        RECT 1670.790 1675.900 1671.110 1676.160 ;
        RECT 1013.910 68.920 1014.230 68.980 ;
        RECT 1670.790 68.920 1671.110 68.980 ;
        RECT 1013.910 68.780 1671.110 68.920 ;
        RECT 1013.910 68.720 1014.230 68.780 ;
        RECT 1670.790 68.720 1671.110 68.780 ;
      LAYER via ;
        RECT 1670.360 1676.920 1670.620 1677.180 ;
        RECT 1670.820 1675.900 1671.080 1676.160 ;
        RECT 1013.940 68.720 1014.200 68.980 ;
        RECT 1670.820 68.720 1671.080 68.980 ;
      LAYER met2 ;
        RECT 1670.280 1700.000 1670.560 1702.400 ;
        RECT 1670.420 1677.210 1670.560 1700.000 ;
        RECT 1670.360 1676.890 1670.620 1677.210 ;
        RECT 1670.820 1675.870 1671.080 1676.190 ;
        RECT 1670.880 69.010 1671.020 1675.870 ;
        RECT 1013.940 68.690 1014.200 69.010 ;
        RECT 1670.820 68.690 1671.080 69.010 ;
        RECT 1014.000 17.410 1014.140 68.690 ;
        RECT 1013.540 17.270 1014.140 17.410 ;
        RECT 1013.540 2.400 1013.680 17.270 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1034.610 64.840 1034.930 64.900 ;
        RECT 1677.230 64.840 1677.550 64.900 ;
        RECT 1034.610 64.700 1677.550 64.840 ;
        RECT 1034.610 64.640 1034.930 64.700 ;
        RECT 1677.230 64.640 1677.550 64.700 ;
        RECT 1031.390 2.960 1031.710 3.020 ;
        RECT 1034.610 2.960 1034.930 3.020 ;
        RECT 1031.390 2.820 1034.930 2.960 ;
        RECT 1031.390 2.760 1031.710 2.820 ;
        RECT 1034.610 2.760 1034.930 2.820 ;
      LAYER via ;
        RECT 1034.640 64.640 1034.900 64.900 ;
        RECT 1677.260 64.640 1677.520 64.900 ;
        RECT 1031.420 2.760 1031.680 3.020 ;
        RECT 1034.640 2.760 1034.900 3.020 ;
      LAYER met2 ;
        RECT 1679.480 1700.410 1679.760 1702.400 ;
        RECT 1677.320 1700.270 1679.760 1700.410 ;
        RECT 1677.320 64.930 1677.460 1700.270 ;
        RECT 1679.480 1700.000 1679.760 1700.270 ;
        RECT 1034.640 64.610 1034.900 64.930 ;
        RECT 1677.260 64.610 1677.520 64.930 ;
        RECT 1034.700 3.050 1034.840 64.610 ;
        RECT 1031.420 2.730 1031.680 3.050 ;
        RECT 1034.640 2.730 1034.900 3.050 ;
        RECT 1031.480 2.400 1031.620 2.730 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1684.665 234.685 1684.835 282.795 ;
        RECT 1684.205 89.845 1684.375 137.955 ;
      LAYER mcon ;
        RECT 1684.665 282.625 1684.835 282.795 ;
        RECT 1684.205 137.785 1684.375 137.955 ;
      LAYER met1 ;
        RECT 1684.590 1642.440 1684.910 1642.500 ;
        RECT 1685.970 1642.440 1686.290 1642.500 ;
        RECT 1684.590 1642.300 1686.290 1642.440 ;
        RECT 1684.590 1642.240 1684.910 1642.300 ;
        RECT 1685.970 1642.240 1686.290 1642.300 ;
        RECT 1684.130 1545.880 1684.450 1545.940 ;
        RECT 1684.590 1545.880 1684.910 1545.940 ;
        RECT 1684.130 1545.740 1684.910 1545.880 ;
        RECT 1684.130 1545.680 1684.450 1545.740 ;
        RECT 1684.590 1545.680 1684.910 1545.740 ;
        RECT 1684.130 786.460 1684.450 786.720 ;
        RECT 1684.220 786.320 1684.360 786.460 ;
        RECT 1684.590 786.320 1684.910 786.380 ;
        RECT 1684.220 786.180 1684.910 786.320 ;
        RECT 1684.590 786.120 1684.910 786.180 ;
        RECT 1684.590 593.880 1684.910 593.940 ;
        RECT 1684.220 593.740 1684.910 593.880 ;
        RECT 1684.220 593.600 1684.360 593.740 ;
        RECT 1684.590 593.680 1684.910 593.740 ;
        RECT 1684.130 593.340 1684.450 593.600 ;
        RECT 1684.130 331.060 1684.450 331.120 ;
        RECT 1684.590 331.060 1684.910 331.120 ;
        RECT 1684.130 330.920 1684.910 331.060 ;
        RECT 1684.130 330.860 1684.450 330.920 ;
        RECT 1684.590 330.860 1684.910 330.920 ;
        RECT 1684.590 282.780 1684.910 282.840 ;
        RECT 1684.395 282.640 1684.910 282.780 ;
        RECT 1684.590 282.580 1684.910 282.640 ;
        RECT 1684.590 234.840 1684.910 234.900 ;
        RECT 1684.395 234.700 1684.910 234.840 ;
        RECT 1684.590 234.640 1684.910 234.700 ;
        RECT 1684.145 137.940 1684.435 137.985 ;
        RECT 1684.590 137.940 1684.910 138.000 ;
        RECT 1684.145 137.800 1684.910 137.940 ;
        RECT 1684.145 137.755 1684.435 137.800 ;
        RECT 1684.590 137.740 1684.910 137.800 ;
        RECT 1684.130 90.000 1684.450 90.060 ;
        RECT 1683.935 89.860 1684.450 90.000 ;
        RECT 1684.130 89.800 1684.450 89.860 ;
        RECT 1055.310 64.160 1055.630 64.220 ;
        RECT 1684.130 64.160 1684.450 64.220 ;
        RECT 1055.310 64.020 1684.450 64.160 ;
        RECT 1055.310 63.960 1055.630 64.020 ;
        RECT 1684.130 63.960 1684.450 64.020 ;
        RECT 1049.330 20.980 1049.650 21.040 ;
        RECT 1055.310 20.980 1055.630 21.040 ;
        RECT 1049.330 20.840 1055.630 20.980 ;
        RECT 1049.330 20.780 1049.650 20.840 ;
        RECT 1055.310 20.780 1055.630 20.840 ;
      LAYER via ;
        RECT 1684.620 1642.240 1684.880 1642.500 ;
        RECT 1686.000 1642.240 1686.260 1642.500 ;
        RECT 1684.160 1545.680 1684.420 1545.940 ;
        RECT 1684.620 1545.680 1684.880 1545.940 ;
        RECT 1684.160 786.460 1684.420 786.720 ;
        RECT 1684.620 786.120 1684.880 786.380 ;
        RECT 1684.620 593.680 1684.880 593.940 ;
        RECT 1684.160 593.340 1684.420 593.600 ;
        RECT 1684.160 330.860 1684.420 331.120 ;
        RECT 1684.620 330.860 1684.880 331.120 ;
        RECT 1684.620 282.580 1684.880 282.840 ;
        RECT 1684.620 234.640 1684.880 234.900 ;
        RECT 1684.620 137.740 1684.880 138.000 ;
        RECT 1684.160 89.800 1684.420 90.060 ;
        RECT 1055.340 63.960 1055.600 64.220 ;
        RECT 1684.160 63.960 1684.420 64.220 ;
        RECT 1049.360 20.780 1049.620 21.040 ;
        RECT 1055.340 20.780 1055.600 21.040 ;
      LAYER met2 ;
        RECT 1688.680 1701.090 1688.960 1702.400 ;
        RECT 1686.060 1700.950 1688.960 1701.090 ;
        RECT 1686.060 1642.530 1686.200 1700.950 ;
        RECT 1688.680 1700.000 1688.960 1700.950 ;
        RECT 1684.620 1642.210 1684.880 1642.530 ;
        RECT 1686.000 1642.210 1686.260 1642.530 ;
        RECT 1684.680 1545.970 1684.820 1642.210 ;
        RECT 1684.160 1545.650 1684.420 1545.970 ;
        RECT 1684.620 1545.650 1684.880 1545.970 ;
        RECT 1684.220 1511.370 1684.360 1545.650 ;
        RECT 1683.760 1511.230 1684.360 1511.370 ;
        RECT 1683.760 1510.690 1683.900 1511.230 ;
        RECT 1683.760 1510.550 1684.360 1510.690 ;
        RECT 1684.220 1414.810 1684.360 1510.550 ;
        RECT 1683.760 1414.670 1684.360 1414.810 ;
        RECT 1683.760 1414.130 1683.900 1414.670 ;
        RECT 1683.760 1413.990 1684.360 1414.130 ;
        RECT 1684.220 1318.250 1684.360 1413.990 ;
        RECT 1683.760 1318.110 1684.360 1318.250 ;
        RECT 1683.760 1317.570 1683.900 1318.110 ;
        RECT 1683.760 1317.430 1684.360 1317.570 ;
        RECT 1684.220 1221.690 1684.360 1317.430 ;
        RECT 1683.760 1221.550 1684.360 1221.690 ;
        RECT 1683.760 1221.010 1683.900 1221.550 ;
        RECT 1683.760 1220.870 1684.360 1221.010 ;
        RECT 1684.220 1125.130 1684.360 1220.870 ;
        RECT 1683.760 1124.990 1684.360 1125.130 ;
        RECT 1683.760 1124.450 1683.900 1124.990 ;
        RECT 1683.760 1124.310 1684.360 1124.450 ;
        RECT 1684.220 1028.570 1684.360 1124.310 ;
        RECT 1683.760 1028.430 1684.360 1028.570 ;
        RECT 1683.760 1027.890 1683.900 1028.430 ;
        RECT 1683.760 1027.750 1684.360 1027.890 ;
        RECT 1684.220 932.010 1684.360 1027.750 ;
        RECT 1683.760 931.870 1684.360 932.010 ;
        RECT 1683.760 931.330 1683.900 931.870 ;
        RECT 1683.760 931.190 1684.360 931.330 ;
        RECT 1684.220 835.450 1684.360 931.190 ;
        RECT 1683.760 835.310 1684.360 835.450 ;
        RECT 1683.760 834.770 1683.900 835.310 ;
        RECT 1683.760 834.630 1684.360 834.770 ;
        RECT 1684.220 786.750 1684.360 834.630 ;
        RECT 1684.160 786.430 1684.420 786.750 ;
        RECT 1684.620 786.090 1684.880 786.410 ;
        RECT 1684.680 690.610 1684.820 786.090 ;
        RECT 1684.680 690.470 1685.280 690.610 ;
        RECT 1685.140 688.570 1685.280 690.470 ;
        RECT 1684.680 688.430 1685.280 688.570 ;
        RECT 1684.680 593.970 1684.820 688.430 ;
        RECT 1684.620 593.650 1684.880 593.970 ;
        RECT 1684.160 593.310 1684.420 593.630 ;
        RECT 1684.220 545.770 1684.360 593.310 ;
        RECT 1683.760 545.630 1684.360 545.770 ;
        RECT 1683.760 545.090 1683.900 545.630 ;
        RECT 1683.760 544.950 1684.360 545.090 ;
        RECT 1684.220 449.210 1684.360 544.950 ;
        RECT 1683.760 449.070 1684.360 449.210 ;
        RECT 1683.760 448.530 1683.900 449.070 ;
        RECT 1683.760 448.390 1684.360 448.530 ;
        RECT 1684.220 331.150 1684.360 448.390 ;
        RECT 1684.160 330.830 1684.420 331.150 ;
        RECT 1684.620 330.830 1684.880 331.150 ;
        RECT 1684.680 282.870 1684.820 330.830 ;
        RECT 1684.620 282.550 1684.880 282.870 ;
        RECT 1684.620 234.610 1684.880 234.930 ;
        RECT 1684.680 138.030 1684.820 234.610 ;
        RECT 1684.620 137.710 1684.880 138.030 ;
        RECT 1684.160 89.770 1684.420 90.090 ;
        RECT 1684.220 64.250 1684.360 89.770 ;
        RECT 1055.340 63.930 1055.600 64.250 ;
        RECT 1684.160 63.930 1684.420 64.250 ;
        RECT 1055.400 21.070 1055.540 63.930 ;
        RECT 1049.360 20.750 1049.620 21.070 ;
        RECT 1055.340 20.750 1055.600 21.070 ;
        RECT 1049.420 2.400 1049.560 20.750 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 64.500 1069.430 64.560 ;
        RECT 1698.390 64.500 1698.710 64.560 ;
        RECT 1069.110 64.360 1698.710 64.500 ;
        RECT 1069.110 64.300 1069.430 64.360 ;
        RECT 1698.390 64.300 1698.710 64.360 ;
      LAYER via ;
        RECT 1069.140 64.300 1069.400 64.560 ;
        RECT 1698.420 64.300 1698.680 64.560 ;
      LAYER met2 ;
        RECT 1697.880 1700.410 1698.160 1702.400 ;
        RECT 1697.880 1700.270 1698.620 1700.410 ;
        RECT 1697.880 1700.000 1698.160 1700.270 ;
        RECT 1698.480 64.590 1698.620 1700.270 ;
        RECT 1069.140 64.270 1069.400 64.590 ;
        RECT 1698.420 64.270 1698.680 64.590 ;
        RECT 1069.200 17.410 1069.340 64.270 ;
        RECT 1067.360 17.270 1069.340 17.410 ;
        RECT 1067.360 2.400 1067.500 17.270 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 63.820 1090.130 63.880 ;
        RECT 1704.830 63.820 1705.150 63.880 ;
        RECT 1089.810 63.680 1705.150 63.820 ;
        RECT 1089.810 63.620 1090.130 63.680 ;
        RECT 1704.830 63.620 1705.150 63.680 ;
      LAYER via ;
        RECT 1089.840 63.620 1090.100 63.880 ;
        RECT 1704.860 63.620 1705.120 63.880 ;
      LAYER met2 ;
        RECT 1707.080 1700.410 1707.360 1702.400 ;
        RECT 1704.920 1700.270 1707.360 1700.410 ;
        RECT 1704.920 63.910 1705.060 1700.270 ;
        RECT 1707.080 1700.000 1707.360 1700.270 ;
        RECT 1089.840 63.590 1090.100 63.910 ;
        RECT 1704.860 63.590 1705.120 63.910 ;
        RECT 1089.900 17.410 1090.040 63.590 ;
        RECT 1085.300 17.270 1090.040 17.410 ;
        RECT 1085.300 2.400 1085.440 17.270 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1713.185 1642.285 1713.355 1656.395 ;
        RECT 1712.265 1497.785 1712.435 1545.215 ;
        RECT 1712.725 1401.225 1712.895 1414.655 ;
        RECT 1712.725 1304.325 1712.895 1318.095 ;
        RECT 1712.265 1256.045 1712.435 1303.815 ;
        RECT 1712.265 544.765 1712.435 579.615 ;
        RECT 1712.265 386.325 1712.435 434.775 ;
        RECT 1712.265 186.405 1712.435 234.515 ;
      LAYER mcon ;
        RECT 1713.185 1656.225 1713.355 1656.395 ;
        RECT 1712.265 1545.045 1712.435 1545.215 ;
        RECT 1712.725 1414.485 1712.895 1414.655 ;
        RECT 1712.725 1317.925 1712.895 1318.095 ;
        RECT 1712.265 1303.645 1712.435 1303.815 ;
        RECT 1712.265 579.445 1712.435 579.615 ;
        RECT 1712.265 434.605 1712.435 434.775 ;
        RECT 1712.265 234.345 1712.435 234.515 ;
      LAYER met1 ;
        RECT 1713.110 1656.380 1713.430 1656.440 ;
        RECT 1712.915 1656.240 1713.430 1656.380 ;
        RECT 1713.110 1656.180 1713.430 1656.240 ;
        RECT 1713.110 1642.440 1713.430 1642.500 ;
        RECT 1712.915 1642.300 1713.430 1642.440 ;
        RECT 1713.110 1642.240 1713.430 1642.300 ;
        RECT 1713.110 1546.220 1713.430 1546.280 ;
        RECT 1712.280 1546.080 1713.430 1546.220 ;
        RECT 1712.280 1545.940 1712.420 1546.080 ;
        RECT 1713.110 1546.020 1713.430 1546.080 ;
        RECT 1712.190 1545.680 1712.510 1545.940 ;
        RECT 1712.190 1545.200 1712.510 1545.260 ;
        RECT 1711.995 1545.060 1712.510 1545.200 ;
        RECT 1712.190 1545.000 1712.510 1545.060 ;
        RECT 1712.205 1497.940 1712.495 1497.985 ;
        RECT 1712.650 1497.940 1712.970 1498.000 ;
        RECT 1712.205 1497.800 1712.970 1497.940 ;
        RECT 1712.205 1497.755 1712.495 1497.800 ;
        RECT 1712.650 1497.740 1712.970 1497.800 ;
        RECT 1712.650 1414.640 1712.970 1414.700 ;
        RECT 1712.455 1414.500 1712.970 1414.640 ;
        RECT 1712.650 1414.440 1712.970 1414.500 ;
        RECT 1712.650 1401.380 1712.970 1401.440 ;
        RECT 1712.455 1401.240 1712.970 1401.380 ;
        RECT 1712.650 1401.180 1712.970 1401.240 ;
        RECT 1712.650 1318.080 1712.970 1318.140 ;
        RECT 1712.455 1317.940 1712.970 1318.080 ;
        RECT 1712.650 1317.880 1712.970 1317.940 ;
        RECT 1712.650 1304.480 1712.970 1304.540 ;
        RECT 1712.455 1304.340 1712.970 1304.480 ;
        RECT 1712.650 1304.280 1712.970 1304.340 ;
        RECT 1712.205 1303.800 1712.495 1303.845 ;
        RECT 1712.650 1303.800 1712.970 1303.860 ;
        RECT 1712.205 1303.660 1712.970 1303.800 ;
        RECT 1712.205 1303.615 1712.495 1303.660 ;
        RECT 1712.650 1303.600 1712.970 1303.660 ;
        RECT 1712.190 1256.200 1712.510 1256.260 ;
        RECT 1711.995 1256.060 1712.510 1256.200 ;
        RECT 1712.190 1256.000 1712.510 1256.060 ;
        RECT 1713.110 1014.460 1713.430 1014.520 ;
        RECT 1713.570 1014.460 1713.890 1014.520 ;
        RECT 1713.110 1014.320 1713.890 1014.460 ;
        RECT 1713.110 1014.260 1713.430 1014.320 ;
        RECT 1713.570 1014.260 1713.890 1014.320 ;
        RECT 1713.570 983.180 1713.890 983.240 ;
        RECT 1714.490 983.180 1714.810 983.240 ;
        RECT 1713.570 983.040 1714.810 983.180 ;
        RECT 1713.570 982.980 1713.890 983.040 ;
        RECT 1714.490 982.980 1714.810 983.040 ;
        RECT 1711.730 772.720 1712.050 772.780 ;
        RECT 1712.650 772.720 1712.970 772.780 ;
        RECT 1711.730 772.580 1712.970 772.720 ;
        RECT 1711.730 772.520 1712.050 772.580 ;
        RECT 1712.650 772.520 1712.970 772.580 ;
        RECT 1712.650 690.240 1712.970 690.500 ;
        RECT 1712.740 689.820 1712.880 690.240 ;
        RECT 1712.650 689.560 1712.970 689.820 ;
        RECT 1712.190 579.600 1712.510 579.660 ;
        RECT 1711.995 579.460 1712.510 579.600 ;
        RECT 1712.190 579.400 1712.510 579.460 ;
        RECT 1712.190 544.920 1712.510 544.980 ;
        RECT 1711.995 544.780 1712.510 544.920 ;
        RECT 1712.190 544.720 1712.510 544.780 ;
        RECT 1712.190 434.760 1712.510 434.820 ;
        RECT 1711.995 434.620 1712.510 434.760 ;
        RECT 1712.190 434.560 1712.510 434.620 ;
        RECT 1712.190 386.480 1712.510 386.540 ;
        RECT 1711.995 386.340 1712.510 386.480 ;
        RECT 1712.190 386.280 1712.510 386.340 ;
        RECT 1712.190 255.380 1712.510 255.640 ;
        RECT 1712.280 254.960 1712.420 255.380 ;
        RECT 1712.190 254.700 1712.510 254.960 ;
        RECT 1712.190 234.500 1712.510 234.560 ;
        RECT 1711.995 234.360 1712.510 234.500 ;
        RECT 1712.190 234.300 1712.510 234.360 ;
        RECT 1712.205 186.560 1712.495 186.605 ;
        RECT 1712.650 186.560 1712.970 186.620 ;
        RECT 1712.205 186.420 1712.970 186.560 ;
        RECT 1712.205 186.375 1712.495 186.420 ;
        RECT 1712.650 186.360 1712.970 186.420 ;
        RECT 1103.610 63.480 1103.930 63.540 ;
        RECT 1711.730 63.480 1712.050 63.540 ;
        RECT 1103.610 63.340 1712.050 63.480 ;
        RECT 1103.610 63.280 1103.930 63.340 ;
        RECT 1711.730 63.280 1712.050 63.340 ;
        RECT 1102.690 2.960 1103.010 3.020 ;
        RECT 1103.610 2.960 1103.930 3.020 ;
        RECT 1102.690 2.820 1103.930 2.960 ;
        RECT 1102.690 2.760 1103.010 2.820 ;
        RECT 1103.610 2.760 1103.930 2.820 ;
      LAYER via ;
        RECT 1713.140 1656.180 1713.400 1656.440 ;
        RECT 1713.140 1642.240 1713.400 1642.500 ;
        RECT 1713.140 1546.020 1713.400 1546.280 ;
        RECT 1712.220 1545.680 1712.480 1545.940 ;
        RECT 1712.220 1545.000 1712.480 1545.260 ;
        RECT 1712.680 1497.740 1712.940 1498.000 ;
        RECT 1712.680 1414.440 1712.940 1414.700 ;
        RECT 1712.680 1401.180 1712.940 1401.440 ;
        RECT 1712.680 1317.880 1712.940 1318.140 ;
        RECT 1712.680 1304.280 1712.940 1304.540 ;
        RECT 1712.680 1303.600 1712.940 1303.860 ;
        RECT 1712.220 1256.000 1712.480 1256.260 ;
        RECT 1713.140 1014.260 1713.400 1014.520 ;
        RECT 1713.600 1014.260 1713.860 1014.520 ;
        RECT 1713.600 982.980 1713.860 983.240 ;
        RECT 1714.520 982.980 1714.780 983.240 ;
        RECT 1711.760 772.520 1712.020 772.780 ;
        RECT 1712.680 772.520 1712.940 772.780 ;
        RECT 1712.680 690.240 1712.940 690.500 ;
        RECT 1712.680 689.560 1712.940 689.820 ;
        RECT 1712.220 579.400 1712.480 579.660 ;
        RECT 1712.220 544.720 1712.480 544.980 ;
        RECT 1712.220 434.560 1712.480 434.820 ;
        RECT 1712.220 386.280 1712.480 386.540 ;
        RECT 1712.220 255.380 1712.480 255.640 ;
        RECT 1712.220 254.700 1712.480 254.960 ;
        RECT 1712.220 234.300 1712.480 234.560 ;
        RECT 1712.680 186.360 1712.940 186.620 ;
        RECT 1103.640 63.280 1103.900 63.540 ;
        RECT 1711.760 63.280 1712.020 63.540 ;
        RECT 1102.720 2.760 1102.980 3.020 ;
        RECT 1103.640 2.760 1103.900 3.020 ;
      LAYER met2 ;
        RECT 1716.280 1701.090 1716.560 1702.400 ;
        RECT 1713.660 1700.950 1716.560 1701.090 ;
        RECT 1713.660 1690.210 1713.800 1700.950 ;
        RECT 1716.280 1700.000 1716.560 1700.950 ;
        RECT 1713.200 1690.070 1713.800 1690.210 ;
        RECT 1713.200 1656.470 1713.340 1690.070 ;
        RECT 1713.140 1656.150 1713.400 1656.470 ;
        RECT 1713.140 1642.210 1713.400 1642.530 ;
        RECT 1713.200 1546.310 1713.340 1642.210 ;
        RECT 1713.140 1545.990 1713.400 1546.310 ;
        RECT 1712.220 1545.650 1712.480 1545.970 ;
        RECT 1712.280 1545.290 1712.420 1545.650 ;
        RECT 1712.220 1544.970 1712.480 1545.290 ;
        RECT 1712.680 1497.710 1712.940 1498.030 ;
        RECT 1712.740 1497.260 1712.880 1497.710 ;
        RECT 1712.740 1497.120 1713.800 1497.260 ;
        RECT 1713.660 1449.490 1713.800 1497.120 ;
        RECT 1712.740 1449.350 1713.800 1449.490 ;
        RECT 1712.740 1414.730 1712.880 1449.350 ;
        RECT 1712.680 1414.410 1712.940 1414.730 ;
        RECT 1712.680 1401.150 1712.940 1401.470 ;
        RECT 1712.740 1400.700 1712.880 1401.150 ;
        RECT 1712.740 1400.560 1713.800 1400.700 ;
        RECT 1713.660 1352.930 1713.800 1400.560 ;
        RECT 1712.740 1352.790 1713.800 1352.930 ;
        RECT 1712.740 1318.170 1712.880 1352.790 ;
        RECT 1712.680 1317.850 1712.940 1318.170 ;
        RECT 1712.680 1304.250 1712.940 1304.570 ;
        RECT 1712.740 1303.890 1712.880 1304.250 ;
        RECT 1712.680 1303.570 1712.940 1303.890 ;
        RECT 1712.220 1255.970 1712.480 1256.290 ;
        RECT 1712.280 1255.805 1712.420 1255.970 ;
        RECT 1712.210 1255.435 1712.490 1255.805 ;
        RECT 1713.130 1255.435 1713.410 1255.805 ;
        RECT 1713.200 1207.580 1713.340 1255.435 ;
        RECT 1713.200 1207.440 1713.800 1207.580 ;
        RECT 1713.660 1172.730 1713.800 1207.440 ;
        RECT 1712.280 1172.590 1713.800 1172.730 ;
        RECT 1712.280 1159.245 1712.420 1172.590 ;
        RECT 1712.210 1158.875 1712.490 1159.245 ;
        RECT 1713.590 1158.875 1713.870 1159.245 ;
        RECT 1713.660 1064.045 1713.800 1158.875 ;
        RECT 1713.590 1063.675 1713.870 1064.045 ;
        RECT 1712.210 1062.570 1712.490 1062.855 ;
        RECT 1712.210 1062.485 1713.340 1062.570 ;
        RECT 1712.280 1062.430 1713.340 1062.485 ;
        RECT 1713.200 1014.550 1713.340 1062.430 ;
        RECT 1713.140 1014.230 1713.400 1014.550 ;
        RECT 1713.600 1014.230 1713.860 1014.550 ;
        RECT 1713.660 983.270 1713.800 1014.230 ;
        RECT 1713.600 982.950 1713.860 983.270 ;
        RECT 1714.520 982.950 1714.780 983.270 ;
        RECT 1714.580 959.325 1714.720 982.950 ;
        RECT 1713.590 958.955 1713.870 959.325 ;
        RECT 1714.510 958.955 1714.790 959.325 ;
        RECT 1713.660 862.765 1713.800 958.955 ;
        RECT 1712.210 862.395 1712.490 862.765 ;
        RECT 1713.590 862.395 1713.870 862.765 ;
        RECT 1712.280 833.410 1712.420 862.395 ;
        RECT 1712.280 833.270 1712.880 833.410 ;
        RECT 1712.740 821.000 1712.880 833.270 ;
        RECT 1712.280 820.860 1712.880 821.000 ;
        RECT 1712.280 787.170 1712.420 820.860 ;
        RECT 1711.820 787.030 1712.420 787.170 ;
        RECT 1711.820 773.685 1711.960 787.030 ;
        RECT 1711.750 773.315 1712.030 773.685 ;
        RECT 1712.210 772.890 1712.490 773.005 ;
        RECT 1712.210 772.810 1712.880 772.890 ;
        RECT 1711.760 772.490 1712.020 772.810 ;
        RECT 1712.210 772.750 1712.940 772.810 ;
        RECT 1712.210 772.635 1712.490 772.750 ;
        RECT 1712.680 772.490 1712.940 772.750 ;
        RECT 1711.820 724.725 1711.960 772.490 ;
        RECT 1712.740 772.335 1712.880 772.490 ;
        RECT 1711.750 724.355 1712.030 724.725 ;
        RECT 1712.670 724.355 1712.950 724.725 ;
        RECT 1712.740 690.530 1712.880 724.355 ;
        RECT 1712.680 690.210 1712.940 690.530 ;
        RECT 1712.680 689.530 1712.940 689.850 ;
        RECT 1712.740 580.565 1712.880 689.530 ;
        RECT 1712.670 580.195 1712.950 580.565 ;
        RECT 1712.210 579.515 1712.490 579.885 ;
        RECT 1712.220 579.370 1712.480 579.515 ;
        RECT 1712.220 544.690 1712.480 545.010 ;
        RECT 1712.280 507.010 1712.420 544.690 ;
        RECT 1711.820 506.870 1712.420 507.010 ;
        RECT 1711.820 496.810 1711.960 506.870 ;
        RECT 1711.820 496.670 1712.420 496.810 ;
        RECT 1712.280 434.850 1712.420 496.670 ;
        RECT 1712.220 434.530 1712.480 434.850 ;
        RECT 1712.220 386.250 1712.480 386.570 ;
        RECT 1712.280 255.670 1712.420 386.250 ;
        RECT 1712.220 255.350 1712.480 255.670 ;
        RECT 1712.220 254.670 1712.480 254.990 ;
        RECT 1712.280 234.590 1712.420 254.670 ;
        RECT 1712.220 234.270 1712.480 234.590 ;
        RECT 1712.680 186.330 1712.940 186.650 ;
        RECT 1712.740 144.740 1712.880 186.330 ;
        RECT 1711.820 144.600 1712.880 144.740 ;
        RECT 1711.820 63.570 1711.960 144.600 ;
        RECT 1103.640 63.250 1103.900 63.570 ;
        RECT 1711.760 63.250 1712.020 63.570 ;
        RECT 1103.700 3.050 1103.840 63.250 ;
        RECT 1102.720 2.730 1102.980 3.050 ;
        RECT 1103.640 2.730 1103.900 3.050 ;
        RECT 1102.780 2.400 1102.920 2.730 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
      LAYER via2 ;
        RECT 1712.210 1255.480 1712.490 1255.760 ;
        RECT 1713.130 1255.480 1713.410 1255.760 ;
        RECT 1712.210 1158.920 1712.490 1159.200 ;
        RECT 1713.590 1158.920 1713.870 1159.200 ;
        RECT 1713.590 1063.720 1713.870 1064.000 ;
        RECT 1712.210 1062.530 1712.490 1062.810 ;
        RECT 1713.590 959.000 1713.870 959.280 ;
        RECT 1714.510 959.000 1714.790 959.280 ;
        RECT 1712.210 862.440 1712.490 862.720 ;
        RECT 1713.590 862.440 1713.870 862.720 ;
        RECT 1711.750 773.360 1712.030 773.640 ;
        RECT 1712.210 772.680 1712.490 772.960 ;
        RECT 1711.750 724.400 1712.030 724.680 ;
        RECT 1712.670 724.400 1712.950 724.680 ;
        RECT 1712.670 580.240 1712.950 580.520 ;
        RECT 1712.210 579.560 1712.490 579.840 ;
      LAYER met3 ;
        RECT 1712.185 1255.770 1712.515 1255.785 ;
        RECT 1713.105 1255.770 1713.435 1255.785 ;
        RECT 1712.185 1255.470 1713.435 1255.770 ;
        RECT 1712.185 1255.455 1712.515 1255.470 ;
        RECT 1713.105 1255.455 1713.435 1255.470 ;
        RECT 1712.185 1159.210 1712.515 1159.225 ;
        RECT 1713.565 1159.210 1713.895 1159.225 ;
        RECT 1712.185 1158.910 1713.895 1159.210 ;
        RECT 1712.185 1158.895 1712.515 1158.910 ;
        RECT 1713.565 1158.895 1713.895 1158.910 ;
        RECT 1713.565 1064.010 1713.895 1064.025 ;
        RECT 1711.510 1063.710 1713.895 1064.010 ;
        RECT 1711.510 1062.820 1711.810 1063.710 ;
        RECT 1713.565 1063.695 1713.895 1063.710 ;
        RECT 1712.185 1062.820 1712.515 1062.835 ;
        RECT 1711.510 1062.520 1712.515 1062.820 ;
        RECT 1712.185 1062.505 1712.515 1062.520 ;
        RECT 1713.565 959.290 1713.895 959.305 ;
        RECT 1714.485 959.290 1714.815 959.305 ;
        RECT 1713.565 958.990 1714.815 959.290 ;
        RECT 1713.565 958.975 1713.895 958.990 ;
        RECT 1714.485 958.975 1714.815 958.990 ;
        RECT 1712.185 862.730 1712.515 862.745 ;
        RECT 1713.565 862.730 1713.895 862.745 ;
        RECT 1712.185 862.430 1713.895 862.730 ;
        RECT 1712.185 862.415 1712.515 862.430 ;
        RECT 1713.565 862.415 1713.895 862.430 ;
        RECT 1711.725 773.650 1712.055 773.665 ;
        RECT 1711.510 773.335 1712.055 773.650 ;
        RECT 1711.510 772.970 1711.810 773.335 ;
        RECT 1712.185 772.970 1712.515 772.985 ;
        RECT 1711.510 772.670 1712.515 772.970 ;
        RECT 1712.185 772.655 1712.515 772.670 ;
        RECT 1711.725 724.690 1712.055 724.705 ;
        RECT 1712.645 724.690 1712.975 724.705 ;
        RECT 1711.725 724.390 1712.975 724.690 ;
        RECT 1711.725 724.375 1712.055 724.390 ;
        RECT 1712.645 724.375 1712.975 724.390 ;
        RECT 1712.645 580.530 1712.975 580.545 ;
        RECT 1712.430 580.215 1712.975 580.530 ;
        RECT 1712.430 579.865 1712.730 580.215 ;
        RECT 1712.185 579.550 1712.730 579.865 ;
        RECT 1712.185 579.535 1712.515 579.550 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1120.630 35.940 1120.950 36.000 ;
        RECT 1725.530 35.940 1725.850 36.000 ;
        RECT 1120.630 35.800 1725.850 35.940 ;
        RECT 1120.630 35.740 1120.950 35.800 ;
        RECT 1725.530 35.740 1725.850 35.800 ;
      LAYER via ;
        RECT 1120.660 35.740 1120.920 36.000 ;
        RECT 1725.560 35.740 1725.820 36.000 ;
      LAYER met2 ;
        RECT 1725.480 1700.000 1725.760 1702.400 ;
        RECT 1725.620 36.030 1725.760 1700.000 ;
        RECT 1120.660 35.710 1120.920 36.030 ;
        RECT 1725.560 35.710 1725.820 36.030 ;
        RECT 1120.720 2.400 1120.860 35.710 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1138.570 35.600 1138.890 35.660 ;
        RECT 1731.970 35.600 1732.290 35.660 ;
        RECT 1138.570 35.460 1732.290 35.600 ;
        RECT 1138.570 35.400 1138.890 35.460 ;
        RECT 1731.970 35.400 1732.290 35.460 ;
      LAYER via ;
        RECT 1138.600 35.400 1138.860 35.660 ;
        RECT 1732.000 35.400 1732.260 35.660 ;
      LAYER met2 ;
        RECT 1734.680 1700.410 1734.960 1702.400 ;
        RECT 1732.060 1700.270 1734.960 1700.410 ;
        RECT 1732.060 35.690 1732.200 1700.270 ;
        RECT 1734.680 1700.000 1734.960 1700.270 ;
        RECT 1138.600 35.370 1138.860 35.690 ;
        RECT 1732.000 35.370 1732.260 35.690 ;
        RECT 1138.660 2.400 1138.800 35.370 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1740.325 1207.425 1740.495 1273.215 ;
        RECT 1740.325 1151.665 1740.495 1193.655 ;
        RECT 1739.865 778.685 1740.035 821.015 ;
        RECT 1739.865 723.945 1740.035 765.935 ;
        RECT 1739.405 61.965 1739.575 113.815 ;
      LAYER mcon ;
        RECT 1740.325 1273.045 1740.495 1273.215 ;
        RECT 1740.325 1193.485 1740.495 1193.655 ;
        RECT 1739.865 820.845 1740.035 821.015 ;
        RECT 1739.865 765.765 1740.035 765.935 ;
        RECT 1739.405 113.645 1739.575 113.815 ;
      LAYER met1 ;
        RECT 1739.790 1593.820 1740.110 1593.880 ;
        RECT 1740.250 1593.820 1740.570 1593.880 ;
        RECT 1739.790 1593.680 1740.570 1593.820 ;
        RECT 1739.790 1593.620 1740.110 1593.680 ;
        RECT 1740.250 1593.620 1740.570 1593.680 ;
        RECT 1739.790 1511.340 1740.110 1511.600 ;
        RECT 1739.880 1510.920 1740.020 1511.340 ;
        RECT 1739.790 1510.660 1740.110 1510.920 ;
        RECT 1739.790 1448.780 1740.110 1449.040 ;
        RECT 1739.880 1448.640 1740.020 1448.780 ;
        RECT 1740.250 1448.640 1740.570 1448.700 ;
        RECT 1739.880 1448.500 1740.570 1448.640 ;
        RECT 1740.250 1448.440 1740.570 1448.500 ;
        RECT 1740.250 1394.240 1740.570 1394.300 ;
        RECT 1739.880 1394.100 1740.570 1394.240 ;
        RECT 1739.880 1393.960 1740.020 1394.100 ;
        RECT 1740.250 1394.040 1740.570 1394.100 ;
        RECT 1739.790 1393.700 1740.110 1393.960 ;
        RECT 1740.250 1304.280 1740.570 1304.540 ;
        RECT 1740.340 1304.140 1740.480 1304.280 ;
        RECT 1740.710 1304.140 1741.030 1304.200 ;
        RECT 1740.340 1304.000 1741.030 1304.140 ;
        RECT 1740.710 1303.940 1741.030 1304.000 ;
        RECT 1740.265 1273.200 1740.555 1273.245 ;
        RECT 1740.710 1273.200 1741.030 1273.260 ;
        RECT 1740.265 1273.060 1741.030 1273.200 ;
        RECT 1740.265 1273.015 1740.555 1273.060 ;
        RECT 1740.710 1273.000 1741.030 1273.060 ;
        RECT 1740.250 1207.580 1740.570 1207.640 ;
        RECT 1740.055 1207.440 1740.570 1207.580 ;
        RECT 1740.250 1207.380 1740.570 1207.440 ;
        RECT 1740.250 1193.640 1740.570 1193.700 ;
        RECT 1740.055 1193.500 1740.570 1193.640 ;
        RECT 1740.250 1193.440 1740.570 1193.500 ;
        RECT 1740.250 1151.820 1740.570 1151.880 ;
        RECT 1740.055 1151.680 1740.570 1151.820 ;
        RECT 1740.250 1151.620 1740.570 1151.680 ;
        RECT 1739.790 1062.740 1740.110 1062.800 ;
        RECT 1740.710 1062.740 1741.030 1062.800 ;
        RECT 1739.790 1062.600 1741.030 1062.740 ;
        RECT 1739.790 1062.540 1740.110 1062.600 ;
        RECT 1740.710 1062.540 1741.030 1062.600 ;
        RECT 1739.790 1028.200 1740.110 1028.460 ;
        RECT 1739.880 1027.720 1740.020 1028.200 ;
        RECT 1740.250 1027.720 1740.570 1027.780 ;
        RECT 1739.880 1027.580 1740.570 1027.720 ;
        RECT 1740.250 1027.520 1740.570 1027.580 ;
        RECT 1739.790 966.180 1740.110 966.240 ;
        RECT 1740.710 966.180 1741.030 966.240 ;
        RECT 1739.790 966.040 1741.030 966.180 ;
        RECT 1739.790 965.980 1740.110 966.040 ;
        RECT 1740.710 965.980 1741.030 966.040 ;
        RECT 1739.790 869.620 1740.110 869.680 ;
        RECT 1740.710 869.620 1741.030 869.680 ;
        RECT 1739.790 869.480 1741.030 869.620 ;
        RECT 1739.790 869.420 1740.110 869.480 ;
        RECT 1740.710 869.420 1741.030 869.480 ;
        RECT 1739.790 821.000 1740.110 821.060 ;
        RECT 1739.595 820.860 1740.110 821.000 ;
        RECT 1739.790 820.800 1740.110 820.860 ;
        RECT 1739.790 778.840 1740.110 778.900 ;
        RECT 1739.595 778.700 1740.110 778.840 ;
        RECT 1739.790 778.640 1740.110 778.700 ;
        RECT 1739.790 765.920 1740.110 765.980 ;
        RECT 1739.595 765.780 1740.110 765.920 ;
        RECT 1739.790 765.720 1740.110 765.780 ;
        RECT 1739.790 724.100 1740.110 724.160 ;
        RECT 1739.595 723.960 1740.110 724.100 ;
        RECT 1739.790 723.900 1740.110 723.960 ;
        RECT 1739.790 579.600 1740.110 579.660 ;
        RECT 1740.250 579.600 1740.570 579.660 ;
        RECT 1739.790 579.460 1740.570 579.600 ;
        RECT 1739.790 579.400 1740.110 579.460 ;
        RECT 1740.250 579.400 1740.570 579.460 ;
        RECT 1739.330 386.620 1739.650 386.880 ;
        RECT 1739.420 386.200 1739.560 386.620 ;
        RECT 1739.330 385.940 1739.650 386.200 ;
        RECT 1739.330 338.200 1739.650 338.260 ;
        RECT 1740.250 338.200 1740.570 338.260 ;
        RECT 1739.330 338.060 1740.570 338.200 ;
        RECT 1739.330 338.000 1739.650 338.060 ;
        RECT 1740.250 338.000 1740.570 338.060 ;
        RECT 1739.790 289.920 1740.110 289.980 ;
        RECT 1740.250 289.920 1740.570 289.980 ;
        RECT 1739.790 289.780 1740.570 289.920 ;
        RECT 1739.790 289.720 1740.110 289.780 ;
        RECT 1740.250 289.720 1740.570 289.780 ;
        RECT 1740.250 144.740 1740.570 144.800 ;
        RECT 1740.710 144.740 1741.030 144.800 ;
        RECT 1740.250 144.600 1741.030 144.740 ;
        RECT 1740.250 144.540 1740.570 144.600 ;
        RECT 1740.710 144.540 1741.030 144.600 ;
        RECT 1739.345 113.800 1739.635 113.845 ;
        RECT 1740.710 113.800 1741.030 113.860 ;
        RECT 1739.345 113.660 1741.030 113.800 ;
        RECT 1739.345 113.615 1739.635 113.660 ;
        RECT 1740.710 113.600 1741.030 113.660 ;
        RECT 1739.330 62.120 1739.650 62.180 ;
        RECT 1739.135 61.980 1739.650 62.120 ;
        RECT 1739.330 61.920 1739.650 61.980 ;
        RECT 1156.510 37.980 1156.830 38.040 ;
        RECT 1739.330 37.980 1739.650 38.040 ;
        RECT 1156.510 37.840 1739.650 37.980 ;
        RECT 1156.510 37.780 1156.830 37.840 ;
        RECT 1739.330 37.780 1739.650 37.840 ;
      LAYER via ;
        RECT 1739.820 1593.620 1740.080 1593.880 ;
        RECT 1740.280 1593.620 1740.540 1593.880 ;
        RECT 1739.820 1511.340 1740.080 1511.600 ;
        RECT 1739.820 1510.660 1740.080 1510.920 ;
        RECT 1739.820 1448.780 1740.080 1449.040 ;
        RECT 1740.280 1448.440 1740.540 1448.700 ;
        RECT 1740.280 1394.040 1740.540 1394.300 ;
        RECT 1739.820 1393.700 1740.080 1393.960 ;
        RECT 1740.280 1304.280 1740.540 1304.540 ;
        RECT 1740.740 1303.940 1741.000 1304.200 ;
        RECT 1740.740 1273.000 1741.000 1273.260 ;
        RECT 1740.280 1207.380 1740.540 1207.640 ;
        RECT 1740.280 1193.440 1740.540 1193.700 ;
        RECT 1740.280 1151.620 1740.540 1151.880 ;
        RECT 1739.820 1062.540 1740.080 1062.800 ;
        RECT 1740.740 1062.540 1741.000 1062.800 ;
        RECT 1739.820 1028.200 1740.080 1028.460 ;
        RECT 1740.280 1027.520 1740.540 1027.780 ;
        RECT 1739.820 965.980 1740.080 966.240 ;
        RECT 1740.740 965.980 1741.000 966.240 ;
        RECT 1739.820 869.420 1740.080 869.680 ;
        RECT 1740.740 869.420 1741.000 869.680 ;
        RECT 1739.820 820.800 1740.080 821.060 ;
        RECT 1739.820 778.640 1740.080 778.900 ;
        RECT 1739.820 765.720 1740.080 765.980 ;
        RECT 1739.820 723.900 1740.080 724.160 ;
        RECT 1739.820 579.400 1740.080 579.660 ;
        RECT 1740.280 579.400 1740.540 579.660 ;
        RECT 1739.360 386.620 1739.620 386.880 ;
        RECT 1739.360 385.940 1739.620 386.200 ;
        RECT 1739.360 338.000 1739.620 338.260 ;
        RECT 1740.280 338.000 1740.540 338.260 ;
        RECT 1739.820 289.720 1740.080 289.980 ;
        RECT 1740.280 289.720 1740.540 289.980 ;
        RECT 1740.280 144.540 1740.540 144.800 ;
        RECT 1740.740 144.540 1741.000 144.800 ;
        RECT 1740.740 113.600 1741.000 113.860 ;
        RECT 1739.360 61.920 1739.620 62.180 ;
        RECT 1156.540 37.780 1156.800 38.040 ;
        RECT 1739.360 37.780 1739.620 38.040 ;
      LAYER met2 ;
        RECT 1743.880 1701.090 1744.160 1702.400 ;
        RECT 1741.260 1700.950 1744.160 1701.090 ;
        RECT 1741.260 1677.970 1741.400 1700.950 ;
        RECT 1743.880 1700.000 1744.160 1700.950 ;
        RECT 1739.880 1677.830 1741.400 1677.970 ;
        RECT 1739.880 1618.130 1740.020 1677.830 ;
        RECT 1739.880 1617.990 1740.480 1618.130 ;
        RECT 1740.340 1593.910 1740.480 1617.990 ;
        RECT 1739.820 1593.590 1740.080 1593.910 ;
        RECT 1740.280 1593.590 1740.540 1593.910 ;
        RECT 1739.880 1511.630 1740.020 1593.590 ;
        RECT 1739.820 1511.310 1740.080 1511.630 ;
        RECT 1739.820 1510.630 1740.080 1510.950 ;
        RECT 1739.880 1449.070 1740.020 1510.630 ;
        RECT 1739.820 1448.750 1740.080 1449.070 ;
        RECT 1740.280 1448.410 1740.540 1448.730 ;
        RECT 1740.340 1394.330 1740.480 1448.410 ;
        RECT 1739.880 1393.990 1740.020 1394.145 ;
        RECT 1740.280 1394.010 1740.540 1394.330 ;
        RECT 1739.820 1393.730 1740.080 1393.990 ;
        RECT 1739.820 1393.670 1740.480 1393.730 ;
        RECT 1739.880 1393.590 1740.480 1393.670 ;
        RECT 1740.340 1387.045 1740.480 1393.590 ;
        RECT 1739.350 1386.675 1739.630 1387.045 ;
        RECT 1740.270 1386.675 1740.550 1387.045 ;
        RECT 1739.420 1344.090 1739.560 1386.675 ;
        RECT 1739.420 1343.950 1740.480 1344.090 ;
        RECT 1740.340 1304.570 1740.480 1343.950 ;
        RECT 1740.280 1304.250 1740.540 1304.570 ;
        RECT 1740.740 1303.910 1741.000 1304.230 ;
        RECT 1740.800 1273.290 1740.940 1303.910 ;
        RECT 1740.740 1272.970 1741.000 1273.290 ;
        RECT 1740.280 1207.350 1740.540 1207.670 ;
        RECT 1740.340 1193.730 1740.480 1207.350 ;
        RECT 1740.280 1193.410 1740.540 1193.730 ;
        RECT 1740.280 1151.590 1740.540 1151.910 ;
        RECT 1740.340 1087.050 1740.480 1151.590 ;
        RECT 1740.340 1086.910 1740.940 1087.050 ;
        RECT 1740.800 1062.830 1740.940 1086.910 ;
        RECT 1739.820 1062.510 1740.080 1062.830 ;
        RECT 1740.740 1062.510 1741.000 1062.830 ;
        RECT 1739.880 1028.490 1740.020 1062.510 ;
        RECT 1739.820 1028.170 1740.080 1028.490 ;
        RECT 1740.280 1027.490 1740.540 1027.810 ;
        RECT 1740.340 990.490 1740.480 1027.490 ;
        RECT 1740.340 990.350 1740.940 990.490 ;
        RECT 1740.800 966.270 1740.940 990.350 ;
        RECT 1739.820 966.125 1740.080 966.270 ;
        RECT 1740.740 966.125 1741.000 966.270 ;
        RECT 1739.810 965.755 1740.090 966.125 ;
        RECT 1740.730 965.755 1741.010 966.125 ;
        RECT 1740.800 931.330 1740.940 965.755 ;
        RECT 1740.340 931.190 1740.940 931.330 ;
        RECT 1740.340 893.930 1740.480 931.190 ;
        RECT 1740.340 893.790 1740.940 893.930 ;
        RECT 1740.800 869.710 1740.940 893.790 ;
        RECT 1739.820 869.390 1740.080 869.710 ;
        RECT 1740.740 869.390 1741.000 869.710 ;
        RECT 1739.880 821.090 1740.020 869.390 ;
        RECT 1739.820 820.770 1740.080 821.090 ;
        RECT 1739.820 778.610 1740.080 778.930 ;
        RECT 1739.880 766.010 1740.020 778.610 ;
        RECT 1739.820 765.690 1740.080 766.010 ;
        RECT 1739.820 723.870 1740.080 724.190 ;
        RECT 1739.880 640.970 1740.020 723.870 ;
        RECT 1739.880 640.830 1740.480 640.970 ;
        RECT 1740.340 580.565 1740.480 640.830 ;
        RECT 1740.270 580.195 1740.550 580.565 ;
        RECT 1739.810 579.515 1740.090 579.885 ;
        RECT 1739.820 579.370 1740.080 579.515 ;
        RECT 1740.280 579.370 1740.540 579.690 ;
        RECT 1740.340 507.010 1740.480 579.370 ;
        RECT 1739.880 506.870 1740.480 507.010 ;
        RECT 1739.880 435.725 1740.020 506.870 ;
        RECT 1739.810 435.355 1740.090 435.725 ;
        RECT 1739.350 434.675 1739.630 435.045 ;
        RECT 1739.420 386.910 1739.560 434.675 ;
        RECT 1739.360 386.590 1739.620 386.910 ;
        RECT 1739.360 385.910 1739.620 386.230 ;
        RECT 1739.420 338.290 1739.560 385.910 ;
        RECT 1739.360 337.970 1739.620 338.290 ;
        RECT 1740.280 337.970 1740.540 338.290 ;
        RECT 1740.340 290.010 1740.480 337.970 ;
        RECT 1739.820 289.690 1740.080 290.010 ;
        RECT 1740.280 289.690 1740.540 290.010 ;
        RECT 1739.880 289.410 1740.020 289.690 ;
        RECT 1739.880 289.270 1740.480 289.410 ;
        RECT 1740.340 144.830 1740.480 289.270 ;
        RECT 1740.280 144.510 1740.540 144.830 ;
        RECT 1740.740 144.510 1741.000 144.830 ;
        RECT 1740.800 113.890 1740.940 144.510 ;
        RECT 1740.740 113.570 1741.000 113.890 ;
        RECT 1739.360 61.890 1739.620 62.210 ;
        RECT 1739.420 38.070 1739.560 61.890 ;
        RECT 1156.540 37.750 1156.800 38.070 ;
        RECT 1739.360 37.750 1739.620 38.070 ;
        RECT 1156.600 2.400 1156.740 37.750 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
      LAYER via2 ;
        RECT 1739.350 1386.720 1739.630 1387.000 ;
        RECT 1740.270 1386.720 1740.550 1387.000 ;
        RECT 1739.810 965.800 1740.090 966.080 ;
        RECT 1740.730 965.800 1741.010 966.080 ;
        RECT 1740.270 580.240 1740.550 580.520 ;
        RECT 1739.810 579.560 1740.090 579.840 ;
        RECT 1739.810 435.400 1740.090 435.680 ;
        RECT 1739.350 434.720 1739.630 435.000 ;
      LAYER met3 ;
        RECT 1739.325 1387.010 1739.655 1387.025 ;
        RECT 1740.245 1387.010 1740.575 1387.025 ;
        RECT 1739.325 1386.710 1740.575 1387.010 ;
        RECT 1739.325 1386.695 1739.655 1386.710 ;
        RECT 1740.245 1386.695 1740.575 1386.710 ;
        RECT 1739.785 966.090 1740.115 966.105 ;
        RECT 1740.705 966.090 1741.035 966.105 ;
        RECT 1739.785 965.790 1741.035 966.090 ;
        RECT 1739.785 965.775 1740.115 965.790 ;
        RECT 1740.705 965.775 1741.035 965.790 ;
        RECT 1740.245 580.530 1740.575 580.545 ;
        RECT 1740.030 580.215 1740.575 580.530 ;
        RECT 1740.030 579.865 1740.330 580.215 ;
        RECT 1739.785 579.550 1740.330 579.865 ;
        RECT 1739.785 579.535 1740.115 579.550 ;
        RECT 1739.785 435.690 1740.115 435.705 ;
        RECT 1739.110 435.390 1740.115 435.690 ;
        RECT 1739.110 435.025 1739.410 435.390 ;
        RECT 1739.785 435.375 1740.115 435.390 ;
        RECT 1739.110 434.710 1739.655 435.025 ;
        RECT 1739.325 434.695 1739.655 434.710 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1491.925 1435.225 1492.095 1483.335 ;
        RECT 1491.005 1213.205 1491.175 1255.875 ;
        RECT 1491.465 1056.125 1491.635 1077.375 ;
        RECT 1491.465 1027.905 1491.635 1055.615 ;
        RECT 1491.465 959.225 1491.635 966.195 ;
        RECT 1491.925 917.745 1492.095 932.535 ;
        RECT 1491.465 834.785 1491.635 862.495 ;
        RECT 1491.925 620.925 1492.095 669.035 ;
        RECT 1491.925 572.645 1492.095 596.955 ;
        RECT 1491.005 524.365 1491.175 572.135 ;
        RECT 1491.925 476.085 1492.095 497.335 ;
        RECT 1491.925 427.805 1492.095 448.715 ;
        RECT 1491.465 338.045 1491.635 403.835 ;
        RECT 1491.465 234.685 1491.635 282.795 ;
        RECT 1491.925 161.925 1492.095 210.375 ;
      LAYER mcon ;
        RECT 1491.925 1483.165 1492.095 1483.335 ;
        RECT 1491.005 1255.705 1491.175 1255.875 ;
        RECT 1491.465 1077.205 1491.635 1077.375 ;
        RECT 1491.465 1055.445 1491.635 1055.615 ;
        RECT 1491.465 966.025 1491.635 966.195 ;
        RECT 1491.925 932.365 1492.095 932.535 ;
        RECT 1491.465 862.325 1491.635 862.495 ;
        RECT 1491.925 668.865 1492.095 669.035 ;
        RECT 1491.925 596.785 1492.095 596.955 ;
        RECT 1491.005 571.965 1491.175 572.135 ;
        RECT 1491.925 497.165 1492.095 497.335 ;
        RECT 1491.925 448.545 1492.095 448.715 ;
        RECT 1491.465 403.665 1491.635 403.835 ;
        RECT 1491.465 282.625 1491.635 282.795 ;
        RECT 1491.925 210.205 1492.095 210.375 ;
      LAYER met1 ;
        RECT 1491.390 1511.340 1491.710 1511.600 ;
        RECT 1491.480 1510.520 1491.620 1511.340 ;
        RECT 1491.850 1510.520 1492.170 1510.580 ;
        RECT 1491.480 1510.380 1492.170 1510.520 ;
        RECT 1491.850 1510.320 1492.170 1510.380 ;
        RECT 1491.850 1483.320 1492.170 1483.380 ;
        RECT 1491.655 1483.180 1492.170 1483.320 ;
        RECT 1491.850 1483.120 1492.170 1483.180 ;
        RECT 1491.865 1435.380 1492.155 1435.425 ;
        RECT 1492.310 1435.380 1492.630 1435.440 ;
        RECT 1491.865 1435.240 1492.630 1435.380 ;
        RECT 1491.865 1435.195 1492.155 1435.240 ;
        RECT 1492.310 1435.180 1492.630 1435.240 ;
        RECT 1492.310 1400.700 1492.630 1400.760 ;
        RECT 1491.480 1400.560 1492.630 1400.700 ;
        RECT 1491.480 1400.420 1491.620 1400.560 ;
        RECT 1492.310 1400.500 1492.630 1400.560 ;
        RECT 1491.390 1400.160 1491.710 1400.420 ;
        RECT 1490.945 1255.860 1491.235 1255.905 ;
        RECT 1491.390 1255.860 1491.710 1255.920 ;
        RECT 1490.945 1255.720 1491.710 1255.860 ;
        RECT 1490.945 1255.675 1491.235 1255.720 ;
        RECT 1491.390 1255.660 1491.710 1255.720 ;
        RECT 1490.930 1213.360 1491.250 1213.420 ;
        RECT 1490.735 1213.220 1491.250 1213.360 ;
        RECT 1490.930 1213.160 1491.250 1213.220 ;
        RECT 1490.930 1200.440 1491.250 1200.500 ;
        RECT 1491.390 1200.440 1491.710 1200.500 ;
        RECT 1490.930 1200.300 1491.710 1200.440 ;
        RECT 1490.930 1200.240 1491.250 1200.300 ;
        RECT 1491.390 1200.240 1491.710 1200.300 ;
        RECT 1491.390 1193.640 1491.710 1193.700 ;
        RECT 1492.770 1193.640 1493.090 1193.700 ;
        RECT 1491.390 1193.500 1493.090 1193.640 ;
        RECT 1491.390 1193.440 1491.710 1193.500 ;
        RECT 1492.770 1193.440 1493.090 1193.500 ;
        RECT 1491.850 1104.220 1492.170 1104.280 ;
        RECT 1492.770 1104.220 1493.090 1104.280 ;
        RECT 1491.850 1104.080 1493.090 1104.220 ;
        RECT 1491.850 1104.020 1492.170 1104.080 ;
        RECT 1492.770 1104.020 1493.090 1104.080 ;
        RECT 1491.405 1077.360 1491.695 1077.405 ;
        RECT 1491.850 1077.360 1492.170 1077.420 ;
        RECT 1491.405 1077.220 1492.170 1077.360 ;
        RECT 1491.405 1077.175 1491.695 1077.220 ;
        RECT 1491.850 1077.160 1492.170 1077.220 ;
        RECT 1491.390 1056.280 1491.710 1056.340 ;
        RECT 1491.195 1056.140 1491.710 1056.280 ;
        RECT 1491.390 1056.080 1491.710 1056.140 ;
        RECT 1491.390 1055.600 1491.710 1055.660 ;
        RECT 1491.195 1055.460 1491.710 1055.600 ;
        RECT 1491.390 1055.400 1491.710 1055.460 ;
        RECT 1491.390 1028.060 1491.710 1028.120 ;
        RECT 1491.195 1027.920 1491.710 1028.060 ;
        RECT 1491.390 1027.860 1491.710 1027.920 ;
        RECT 1491.405 966.180 1491.695 966.225 ;
        RECT 1491.850 966.180 1492.170 966.240 ;
        RECT 1491.405 966.040 1492.170 966.180 ;
        RECT 1491.405 965.995 1491.695 966.040 ;
        RECT 1491.850 965.980 1492.170 966.040 ;
        RECT 1491.390 959.380 1491.710 959.440 ;
        RECT 1491.195 959.240 1491.710 959.380 ;
        RECT 1491.390 959.180 1491.710 959.240 ;
        RECT 1491.390 932.520 1491.710 932.580 ;
        RECT 1491.865 932.520 1492.155 932.565 ;
        RECT 1491.390 932.380 1492.155 932.520 ;
        RECT 1491.390 932.320 1491.710 932.380 ;
        RECT 1491.865 932.335 1492.155 932.380 ;
        RECT 1491.850 917.900 1492.170 917.960 ;
        RECT 1491.655 917.760 1492.170 917.900 ;
        RECT 1491.850 917.700 1492.170 917.760 ;
        RECT 1491.850 883.900 1492.170 883.960 ;
        RECT 1491.480 883.760 1492.170 883.900 ;
        RECT 1491.480 883.280 1491.620 883.760 ;
        RECT 1491.850 883.700 1492.170 883.760 ;
        RECT 1491.390 883.020 1491.710 883.280 ;
        RECT 1491.390 862.480 1491.710 862.540 ;
        RECT 1491.195 862.340 1491.710 862.480 ;
        RECT 1491.390 862.280 1491.710 862.340 ;
        RECT 1491.390 834.940 1491.710 835.000 ;
        RECT 1491.195 834.800 1491.710 834.940 ;
        RECT 1491.390 834.740 1491.710 834.800 ;
        RECT 1491.850 669.020 1492.170 669.080 ;
        RECT 1491.655 668.880 1492.170 669.020 ;
        RECT 1491.850 668.820 1492.170 668.880 ;
        RECT 1491.850 621.080 1492.170 621.140 ;
        RECT 1491.655 620.940 1492.170 621.080 ;
        RECT 1491.850 620.880 1492.170 620.940 ;
        RECT 1491.850 596.940 1492.170 597.000 ;
        RECT 1491.655 596.800 1492.170 596.940 ;
        RECT 1491.850 596.740 1492.170 596.800 ;
        RECT 1490.930 572.800 1491.250 572.860 ;
        RECT 1491.865 572.800 1492.155 572.845 ;
        RECT 1490.930 572.660 1492.155 572.800 ;
        RECT 1490.930 572.600 1491.250 572.660 ;
        RECT 1491.865 572.615 1492.155 572.660 ;
        RECT 1490.930 572.120 1491.250 572.180 ;
        RECT 1490.735 571.980 1491.250 572.120 ;
        RECT 1490.930 571.920 1491.250 571.980 ;
        RECT 1490.945 524.520 1491.235 524.565 ;
        RECT 1491.850 524.520 1492.170 524.580 ;
        RECT 1490.945 524.380 1492.170 524.520 ;
        RECT 1490.945 524.335 1491.235 524.380 ;
        RECT 1491.850 524.320 1492.170 524.380 ;
        RECT 1491.850 497.320 1492.170 497.380 ;
        RECT 1491.655 497.180 1492.170 497.320 ;
        RECT 1491.850 497.120 1492.170 497.180 ;
        RECT 1491.850 476.240 1492.170 476.300 ;
        RECT 1491.655 476.100 1492.170 476.240 ;
        RECT 1491.850 476.040 1492.170 476.100 ;
        RECT 1491.850 448.700 1492.170 448.760 ;
        RECT 1491.655 448.560 1492.170 448.700 ;
        RECT 1491.850 448.500 1492.170 448.560 ;
        RECT 1491.850 427.960 1492.170 428.020 ;
        RECT 1491.655 427.820 1492.170 427.960 ;
        RECT 1491.850 427.760 1492.170 427.820 ;
        RECT 1491.405 403.820 1491.695 403.865 ;
        RECT 1491.850 403.820 1492.170 403.880 ;
        RECT 1491.405 403.680 1492.170 403.820 ;
        RECT 1491.405 403.635 1491.695 403.680 ;
        RECT 1491.850 403.620 1492.170 403.680 ;
        RECT 1491.405 338.200 1491.695 338.245 ;
        RECT 1491.850 338.200 1492.170 338.260 ;
        RECT 1491.405 338.060 1492.170 338.200 ;
        RECT 1491.405 338.015 1491.695 338.060 ;
        RECT 1491.850 338.000 1492.170 338.060 ;
        RECT 1491.390 282.780 1491.710 282.840 ;
        RECT 1491.195 282.640 1491.710 282.780 ;
        RECT 1491.390 282.580 1491.710 282.640 ;
        RECT 1491.405 234.840 1491.695 234.885 ;
        RECT 1491.850 234.840 1492.170 234.900 ;
        RECT 1491.405 234.700 1492.170 234.840 ;
        RECT 1491.405 234.655 1491.695 234.700 ;
        RECT 1491.850 234.640 1492.170 234.700 ;
        RECT 1491.850 210.360 1492.170 210.420 ;
        RECT 1491.655 210.220 1492.170 210.360 ;
        RECT 1491.850 210.160 1492.170 210.220 ;
        RECT 1490.930 162.080 1491.250 162.140 ;
        RECT 1491.865 162.080 1492.155 162.125 ;
        RECT 1490.930 161.940 1492.155 162.080 ;
        RECT 1490.930 161.880 1491.250 161.940 ;
        RECT 1491.865 161.895 1492.155 161.940 ;
      LAYER via ;
        RECT 1491.420 1511.340 1491.680 1511.600 ;
        RECT 1491.880 1510.320 1492.140 1510.580 ;
        RECT 1491.880 1483.120 1492.140 1483.380 ;
        RECT 1492.340 1435.180 1492.600 1435.440 ;
        RECT 1492.340 1400.500 1492.600 1400.760 ;
        RECT 1491.420 1400.160 1491.680 1400.420 ;
        RECT 1491.420 1255.660 1491.680 1255.920 ;
        RECT 1490.960 1213.160 1491.220 1213.420 ;
        RECT 1490.960 1200.240 1491.220 1200.500 ;
        RECT 1491.420 1200.240 1491.680 1200.500 ;
        RECT 1491.420 1193.440 1491.680 1193.700 ;
        RECT 1492.800 1193.440 1493.060 1193.700 ;
        RECT 1491.880 1104.020 1492.140 1104.280 ;
        RECT 1492.800 1104.020 1493.060 1104.280 ;
        RECT 1491.880 1077.160 1492.140 1077.420 ;
        RECT 1491.420 1056.080 1491.680 1056.340 ;
        RECT 1491.420 1055.400 1491.680 1055.660 ;
        RECT 1491.420 1027.860 1491.680 1028.120 ;
        RECT 1491.880 965.980 1492.140 966.240 ;
        RECT 1491.420 959.180 1491.680 959.440 ;
        RECT 1491.420 932.320 1491.680 932.580 ;
        RECT 1491.880 917.700 1492.140 917.960 ;
        RECT 1491.880 883.700 1492.140 883.960 ;
        RECT 1491.420 883.020 1491.680 883.280 ;
        RECT 1491.420 862.280 1491.680 862.540 ;
        RECT 1491.420 834.740 1491.680 835.000 ;
        RECT 1491.880 668.820 1492.140 669.080 ;
        RECT 1491.880 620.880 1492.140 621.140 ;
        RECT 1491.880 596.740 1492.140 597.000 ;
        RECT 1490.960 572.600 1491.220 572.860 ;
        RECT 1490.960 571.920 1491.220 572.180 ;
        RECT 1491.880 524.320 1492.140 524.580 ;
        RECT 1491.880 497.120 1492.140 497.380 ;
        RECT 1491.880 476.040 1492.140 476.300 ;
        RECT 1491.880 448.500 1492.140 448.760 ;
        RECT 1491.880 427.760 1492.140 428.020 ;
        RECT 1491.880 403.620 1492.140 403.880 ;
        RECT 1491.880 338.000 1492.140 338.260 ;
        RECT 1491.420 282.580 1491.680 282.840 ;
        RECT 1491.880 234.640 1492.140 234.900 ;
        RECT 1491.880 210.160 1492.140 210.420 ;
        RECT 1490.960 161.880 1491.220 162.140 ;
      LAYER met2 ;
        RECT 1495.940 1700.410 1496.220 1702.400 ;
        RECT 1493.320 1700.270 1496.220 1700.410 ;
        RECT 1493.320 1678.140 1493.460 1700.270 ;
        RECT 1495.940 1700.000 1496.220 1700.270 ;
        RECT 1491.940 1678.000 1493.460 1678.140 ;
        RECT 1491.940 1559.650 1492.080 1678.000 ;
        RECT 1491.480 1559.510 1492.080 1559.650 ;
        RECT 1491.480 1511.630 1491.620 1559.510 ;
        RECT 1491.420 1511.310 1491.680 1511.630 ;
        RECT 1491.880 1510.290 1492.140 1510.610 ;
        RECT 1491.940 1483.410 1492.080 1510.290 ;
        RECT 1491.880 1483.090 1492.140 1483.410 ;
        RECT 1492.340 1435.150 1492.600 1435.470 ;
        RECT 1492.400 1400.790 1492.540 1435.150 ;
        RECT 1492.340 1400.470 1492.600 1400.790 ;
        RECT 1491.420 1400.130 1491.680 1400.450 ;
        RECT 1491.480 1393.845 1491.620 1400.130 ;
        RECT 1491.410 1393.475 1491.690 1393.845 ;
        RECT 1492.790 1393.475 1493.070 1393.845 ;
        RECT 1492.860 1268.610 1493.000 1393.475 ;
        RECT 1491.480 1268.470 1493.000 1268.610 ;
        RECT 1491.480 1255.950 1491.620 1268.470 ;
        RECT 1491.420 1255.630 1491.680 1255.950 ;
        RECT 1490.960 1213.130 1491.220 1213.450 ;
        RECT 1491.020 1200.530 1491.160 1213.130 ;
        RECT 1490.960 1200.210 1491.220 1200.530 ;
        RECT 1491.420 1200.210 1491.680 1200.530 ;
        RECT 1491.480 1193.730 1491.620 1200.210 ;
        RECT 1491.420 1193.410 1491.680 1193.730 ;
        RECT 1492.800 1193.410 1493.060 1193.730 ;
        RECT 1492.860 1104.310 1493.000 1193.410 ;
        RECT 1491.880 1103.990 1492.140 1104.310 ;
        RECT 1492.800 1103.990 1493.060 1104.310 ;
        RECT 1491.940 1077.450 1492.080 1103.990 ;
        RECT 1491.880 1077.130 1492.140 1077.450 ;
        RECT 1491.420 1056.050 1491.680 1056.370 ;
        RECT 1491.480 1055.690 1491.620 1056.050 ;
        RECT 1491.420 1055.370 1491.680 1055.690 ;
        RECT 1491.420 1027.830 1491.680 1028.150 ;
        RECT 1491.480 1007.490 1491.620 1027.830 ;
        RECT 1491.480 1007.350 1492.080 1007.490 ;
        RECT 1491.940 966.270 1492.080 1007.350 ;
        RECT 1491.880 965.950 1492.140 966.270 ;
        RECT 1491.420 959.150 1491.680 959.470 ;
        RECT 1491.480 932.610 1491.620 959.150 ;
        RECT 1491.420 932.290 1491.680 932.610 ;
        RECT 1491.880 917.670 1492.140 917.990 ;
        RECT 1491.940 883.990 1492.080 917.670 ;
        RECT 1491.880 883.670 1492.140 883.990 ;
        RECT 1491.420 882.990 1491.680 883.310 ;
        RECT 1491.480 862.570 1491.620 882.990 ;
        RECT 1491.420 862.250 1491.680 862.570 ;
        RECT 1491.420 834.710 1491.680 835.030 ;
        RECT 1491.480 814.370 1491.620 834.710 ;
        RECT 1491.480 814.230 1492.080 814.370 ;
        RECT 1491.940 669.110 1492.080 814.230 ;
        RECT 1491.880 668.790 1492.140 669.110 ;
        RECT 1491.880 620.850 1492.140 621.170 ;
        RECT 1491.940 597.030 1492.080 620.850 ;
        RECT 1491.880 596.710 1492.140 597.030 ;
        RECT 1490.960 572.570 1491.220 572.890 ;
        RECT 1491.020 572.210 1491.160 572.570 ;
        RECT 1490.960 571.890 1491.220 572.210 ;
        RECT 1491.880 524.290 1492.140 524.610 ;
        RECT 1491.940 497.410 1492.080 524.290 ;
        RECT 1491.880 497.090 1492.140 497.410 ;
        RECT 1491.880 476.010 1492.140 476.330 ;
        RECT 1491.940 448.790 1492.080 476.010 ;
        RECT 1491.880 448.470 1492.140 448.790 ;
        RECT 1491.880 427.730 1492.140 428.050 ;
        RECT 1491.940 403.910 1492.080 427.730 ;
        RECT 1491.880 403.590 1492.140 403.910 ;
        RECT 1491.880 337.970 1492.140 338.290 ;
        RECT 1491.940 289.580 1492.080 337.970 ;
        RECT 1491.480 289.440 1492.080 289.580 ;
        RECT 1491.480 282.870 1491.620 289.440 ;
        RECT 1491.420 282.550 1491.680 282.870 ;
        RECT 1491.880 234.610 1492.140 234.930 ;
        RECT 1491.940 210.450 1492.080 234.610 ;
        RECT 1491.880 210.130 1492.140 210.450 ;
        RECT 1490.960 161.850 1491.220 162.170 ;
        RECT 1491.020 96.970 1491.160 161.850 ;
        RECT 1491.020 96.830 1491.620 96.970 ;
        RECT 1491.480 72.490 1491.620 96.830 ;
        RECT 1491.020 72.350 1491.620 72.490 ;
        RECT 1491.020 48.010 1491.160 72.350 ;
        RECT 1491.020 47.870 1491.620 48.010 ;
        RECT 1491.480 37.925 1491.620 47.870 ;
        RECT 674.450 37.555 674.730 37.925 ;
        RECT 1491.410 37.555 1491.690 37.925 ;
        RECT 674.520 2.400 674.660 37.555 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 1491.410 1393.520 1491.690 1393.800 ;
        RECT 1492.790 1393.520 1493.070 1393.800 ;
        RECT 674.450 37.600 674.730 37.880 ;
        RECT 1491.410 37.600 1491.690 37.880 ;
      LAYER met3 ;
        RECT 1491.385 1393.810 1491.715 1393.825 ;
        RECT 1492.765 1393.810 1493.095 1393.825 ;
        RECT 1491.385 1393.510 1493.095 1393.810 ;
        RECT 1491.385 1393.495 1491.715 1393.510 ;
        RECT 1492.765 1393.495 1493.095 1393.510 ;
        RECT 674.425 37.890 674.755 37.905 ;
        RECT 1491.385 37.890 1491.715 37.905 ;
        RECT 674.425 37.590 1491.715 37.890 ;
        RECT 674.425 37.575 674.755 37.590 ;
        RECT 1491.385 37.575 1491.715 37.590 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1173.990 38.320 1174.310 38.380 ;
        RECT 1753.130 38.320 1753.450 38.380 ;
        RECT 1173.990 38.180 1753.450 38.320 ;
        RECT 1173.990 38.120 1174.310 38.180 ;
        RECT 1753.130 38.120 1753.450 38.180 ;
      LAYER via ;
        RECT 1174.020 38.120 1174.280 38.380 ;
        RECT 1753.160 38.120 1753.420 38.380 ;
      LAYER met2 ;
        RECT 1753.080 1700.000 1753.360 1702.400 ;
        RECT 1753.220 38.410 1753.360 1700.000 ;
        RECT 1174.020 38.090 1174.280 38.410 ;
        RECT 1753.160 38.090 1753.420 38.410 ;
        RECT 1174.080 2.400 1174.220 38.090 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1191.930 35.260 1192.250 35.320 ;
        RECT 1759.570 35.260 1759.890 35.320 ;
        RECT 1191.930 35.120 1759.890 35.260 ;
        RECT 1191.930 35.060 1192.250 35.120 ;
        RECT 1759.570 35.060 1759.890 35.120 ;
      LAYER via ;
        RECT 1191.960 35.060 1192.220 35.320 ;
        RECT 1759.600 35.060 1759.860 35.320 ;
      LAYER met2 ;
        RECT 1762.280 1700.410 1762.560 1702.400 ;
        RECT 1759.660 1700.270 1762.560 1700.410 ;
        RECT 1759.660 35.350 1759.800 1700.270 ;
        RECT 1762.280 1700.000 1762.560 1700.270 ;
        RECT 1191.960 35.030 1192.220 35.350 ;
        RECT 1759.600 35.030 1759.860 35.350 ;
        RECT 1192.020 2.400 1192.160 35.030 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1767.465 1442.025 1767.635 1490.475 ;
        RECT 1767.925 1207.425 1768.095 1273.215 ;
        RECT 1767.465 766.105 1767.635 814.215 ;
        RECT 1767.465 723.945 1767.635 765.595 ;
        RECT 1767.925 572.645 1768.095 579.955 ;
        RECT 1767.465 476.085 1767.635 524.195 ;
        RECT 1767.925 331.245 1768.095 379.355 ;
        RECT 1768.385 96.305 1768.555 137.955 ;
      LAYER mcon ;
        RECT 1767.465 1490.305 1767.635 1490.475 ;
        RECT 1767.925 1273.045 1768.095 1273.215 ;
        RECT 1767.465 814.045 1767.635 814.215 ;
        RECT 1767.465 765.425 1767.635 765.595 ;
        RECT 1767.925 579.785 1768.095 579.955 ;
        RECT 1767.465 524.025 1767.635 524.195 ;
        RECT 1767.925 379.185 1768.095 379.355 ;
        RECT 1768.385 137.785 1768.555 137.955 ;
      LAYER met1 ;
        RECT 1767.390 1593.820 1767.710 1593.880 ;
        RECT 1767.850 1593.820 1768.170 1593.880 ;
        RECT 1767.390 1593.680 1768.170 1593.820 ;
        RECT 1767.390 1593.620 1767.710 1593.680 ;
        RECT 1767.850 1593.620 1768.170 1593.680 ;
        RECT 1767.390 1490.460 1767.710 1490.520 ;
        RECT 1767.195 1490.320 1767.710 1490.460 ;
        RECT 1767.390 1490.260 1767.710 1490.320 ;
        RECT 1767.405 1442.180 1767.695 1442.225 ;
        RECT 1767.850 1442.180 1768.170 1442.240 ;
        RECT 1767.405 1442.040 1768.170 1442.180 ;
        RECT 1767.405 1441.995 1767.695 1442.040 ;
        RECT 1767.850 1441.980 1768.170 1442.040 ;
        RECT 1767.850 1400.700 1768.170 1400.760 ;
        RECT 1768.310 1400.700 1768.630 1400.760 ;
        RECT 1767.850 1400.560 1768.630 1400.700 ;
        RECT 1767.850 1400.500 1768.170 1400.560 ;
        RECT 1768.310 1400.500 1768.630 1400.560 ;
        RECT 1767.865 1273.200 1768.155 1273.245 ;
        RECT 1768.310 1273.200 1768.630 1273.260 ;
        RECT 1767.865 1273.060 1768.630 1273.200 ;
        RECT 1767.865 1273.015 1768.155 1273.060 ;
        RECT 1768.310 1273.000 1768.630 1273.060 ;
        RECT 1767.850 1207.580 1768.170 1207.640 ;
        RECT 1767.655 1207.440 1768.170 1207.580 ;
        RECT 1767.850 1207.380 1768.170 1207.440 ;
        RECT 1767.850 1173.380 1768.170 1173.640 ;
        RECT 1767.940 1172.960 1768.080 1173.380 ;
        RECT 1767.850 1172.700 1768.170 1172.960 ;
        RECT 1767.390 1062.740 1767.710 1062.800 ;
        RECT 1768.310 1062.740 1768.630 1062.800 ;
        RECT 1767.390 1062.600 1768.630 1062.740 ;
        RECT 1767.390 1062.540 1767.710 1062.600 ;
        RECT 1768.310 1062.540 1768.630 1062.600 ;
        RECT 1767.390 1028.200 1767.710 1028.460 ;
        RECT 1767.480 1028.060 1767.620 1028.200 ;
        RECT 1767.850 1028.060 1768.170 1028.120 ;
        RECT 1767.480 1027.920 1768.170 1028.060 ;
        RECT 1767.850 1027.860 1768.170 1027.920 ;
        RECT 1767.390 966.180 1767.710 966.240 ;
        RECT 1768.310 966.180 1768.630 966.240 ;
        RECT 1767.390 966.040 1768.630 966.180 ;
        RECT 1767.390 965.980 1767.710 966.040 ;
        RECT 1768.310 965.980 1768.630 966.040 ;
        RECT 1767.390 869.620 1767.710 869.680 ;
        RECT 1768.310 869.620 1768.630 869.680 ;
        RECT 1767.390 869.480 1768.630 869.620 ;
        RECT 1767.390 869.420 1767.710 869.480 ;
        RECT 1768.310 869.420 1768.630 869.480 ;
        RECT 1767.390 821.000 1767.710 821.060 ;
        RECT 1767.850 821.000 1768.170 821.060 ;
        RECT 1767.390 820.860 1768.170 821.000 ;
        RECT 1767.390 820.800 1767.710 820.860 ;
        RECT 1767.850 820.800 1768.170 820.860 ;
        RECT 1767.390 814.200 1767.710 814.260 ;
        RECT 1767.195 814.060 1767.710 814.200 ;
        RECT 1767.390 814.000 1767.710 814.060 ;
        RECT 1767.390 766.260 1767.710 766.320 ;
        RECT 1767.195 766.120 1767.710 766.260 ;
        RECT 1767.390 766.060 1767.710 766.120 ;
        RECT 1767.390 765.580 1767.710 765.640 ;
        RECT 1767.195 765.440 1767.710 765.580 ;
        RECT 1767.390 765.380 1767.710 765.440 ;
        RECT 1767.390 724.100 1767.710 724.160 ;
        RECT 1767.195 723.960 1767.710 724.100 ;
        RECT 1767.390 723.900 1767.710 723.960 ;
        RECT 1767.850 579.940 1768.170 580.000 ;
        RECT 1767.655 579.800 1768.170 579.940 ;
        RECT 1767.850 579.740 1768.170 579.800 ;
        RECT 1767.850 572.800 1768.170 572.860 ;
        RECT 1767.655 572.660 1768.170 572.800 ;
        RECT 1767.850 572.600 1768.170 572.660 ;
        RECT 1767.390 531.320 1767.710 531.380 ;
        RECT 1767.850 531.320 1768.170 531.380 ;
        RECT 1767.390 531.180 1768.170 531.320 ;
        RECT 1767.390 531.120 1767.710 531.180 ;
        RECT 1767.850 531.120 1768.170 531.180 ;
        RECT 1767.390 524.180 1767.710 524.240 ;
        RECT 1767.195 524.040 1767.710 524.180 ;
        RECT 1767.390 523.980 1767.710 524.040 ;
        RECT 1767.390 476.240 1767.710 476.300 ;
        RECT 1767.195 476.100 1767.710 476.240 ;
        RECT 1767.390 476.040 1767.710 476.100 ;
        RECT 1767.390 434.760 1767.710 434.820 ;
        RECT 1767.850 434.760 1768.170 434.820 ;
        RECT 1767.390 434.620 1768.170 434.760 ;
        RECT 1767.390 434.560 1767.710 434.620 ;
        RECT 1767.850 434.560 1768.170 434.620 ;
        RECT 1767.390 427.420 1767.710 427.680 ;
        RECT 1767.480 427.280 1767.620 427.420 ;
        RECT 1767.850 427.280 1768.170 427.340 ;
        RECT 1767.480 427.140 1768.170 427.280 ;
        RECT 1767.850 427.080 1768.170 427.140 ;
        RECT 1767.850 379.340 1768.170 379.400 ;
        RECT 1767.655 379.200 1768.170 379.340 ;
        RECT 1767.850 379.140 1768.170 379.200 ;
        RECT 1767.865 331.400 1768.155 331.445 ;
        RECT 1768.310 331.400 1768.630 331.460 ;
        RECT 1767.865 331.260 1768.630 331.400 ;
        RECT 1767.865 331.215 1768.155 331.260 ;
        RECT 1768.310 331.200 1768.630 331.260 ;
        RECT 1767.850 144.740 1768.170 144.800 ;
        RECT 1768.310 144.740 1768.630 144.800 ;
        RECT 1767.850 144.600 1768.630 144.740 ;
        RECT 1767.850 144.540 1768.170 144.600 ;
        RECT 1768.310 144.540 1768.630 144.600 ;
        RECT 1768.310 137.940 1768.630 138.000 ;
        RECT 1768.115 137.800 1768.630 137.940 ;
        RECT 1768.310 137.740 1768.630 137.800 ;
        RECT 1768.310 96.460 1768.630 96.520 ;
        RECT 1768.115 96.320 1768.630 96.460 ;
        RECT 1768.310 96.260 1768.630 96.320 ;
        RECT 1209.870 34.920 1210.190 34.980 ;
        RECT 1766.930 34.920 1767.250 34.980 ;
        RECT 1209.870 34.780 1767.250 34.920 ;
        RECT 1209.870 34.720 1210.190 34.780 ;
        RECT 1766.930 34.720 1767.250 34.780 ;
      LAYER via ;
        RECT 1767.420 1593.620 1767.680 1593.880 ;
        RECT 1767.880 1593.620 1768.140 1593.880 ;
        RECT 1767.420 1490.260 1767.680 1490.520 ;
        RECT 1767.880 1441.980 1768.140 1442.240 ;
        RECT 1767.880 1400.500 1768.140 1400.760 ;
        RECT 1768.340 1400.500 1768.600 1400.760 ;
        RECT 1768.340 1273.000 1768.600 1273.260 ;
        RECT 1767.880 1207.380 1768.140 1207.640 ;
        RECT 1767.880 1173.380 1768.140 1173.640 ;
        RECT 1767.880 1172.700 1768.140 1172.960 ;
        RECT 1767.420 1062.540 1767.680 1062.800 ;
        RECT 1768.340 1062.540 1768.600 1062.800 ;
        RECT 1767.420 1028.200 1767.680 1028.460 ;
        RECT 1767.880 1027.860 1768.140 1028.120 ;
        RECT 1767.420 965.980 1767.680 966.240 ;
        RECT 1768.340 965.980 1768.600 966.240 ;
        RECT 1767.420 869.420 1767.680 869.680 ;
        RECT 1768.340 869.420 1768.600 869.680 ;
        RECT 1767.420 820.800 1767.680 821.060 ;
        RECT 1767.880 820.800 1768.140 821.060 ;
        RECT 1767.420 814.000 1767.680 814.260 ;
        RECT 1767.420 766.060 1767.680 766.320 ;
        RECT 1767.420 765.380 1767.680 765.640 ;
        RECT 1767.420 723.900 1767.680 724.160 ;
        RECT 1767.880 579.740 1768.140 580.000 ;
        RECT 1767.880 572.600 1768.140 572.860 ;
        RECT 1767.420 531.120 1767.680 531.380 ;
        RECT 1767.880 531.120 1768.140 531.380 ;
        RECT 1767.420 523.980 1767.680 524.240 ;
        RECT 1767.420 476.040 1767.680 476.300 ;
        RECT 1767.420 434.560 1767.680 434.820 ;
        RECT 1767.880 434.560 1768.140 434.820 ;
        RECT 1767.420 427.420 1767.680 427.680 ;
        RECT 1767.880 427.080 1768.140 427.340 ;
        RECT 1767.880 379.140 1768.140 379.400 ;
        RECT 1768.340 331.200 1768.600 331.460 ;
        RECT 1767.880 144.540 1768.140 144.800 ;
        RECT 1768.340 144.540 1768.600 144.800 ;
        RECT 1768.340 137.740 1768.600 138.000 ;
        RECT 1768.340 96.260 1768.600 96.520 ;
        RECT 1209.900 34.720 1210.160 34.980 ;
        RECT 1766.960 34.720 1767.220 34.980 ;
      LAYER met2 ;
        RECT 1771.020 1700.410 1771.300 1702.400 ;
        RECT 1768.860 1700.270 1771.300 1700.410 ;
        RECT 1768.860 1678.140 1769.000 1700.270 ;
        RECT 1771.020 1700.000 1771.300 1700.270 ;
        RECT 1767.480 1678.000 1769.000 1678.140 ;
        RECT 1767.480 1618.130 1767.620 1678.000 ;
        RECT 1767.480 1617.990 1768.080 1618.130 ;
        RECT 1767.940 1593.910 1768.080 1617.990 ;
        RECT 1767.420 1593.590 1767.680 1593.910 ;
        RECT 1767.880 1593.590 1768.140 1593.910 ;
        RECT 1767.480 1490.550 1767.620 1593.590 ;
        RECT 1767.420 1490.230 1767.680 1490.550 ;
        RECT 1767.880 1441.950 1768.140 1442.270 ;
        RECT 1767.940 1400.790 1768.080 1441.950 ;
        RECT 1767.880 1400.470 1768.140 1400.790 ;
        RECT 1768.340 1400.470 1768.600 1400.790 ;
        RECT 1768.400 1351.570 1768.540 1400.470 ;
        RECT 1768.400 1351.430 1769.000 1351.570 ;
        RECT 1768.860 1350.210 1769.000 1351.430 ;
        RECT 1768.400 1350.070 1769.000 1350.210 ;
        RECT 1768.400 1273.290 1768.540 1350.070 ;
        RECT 1768.340 1272.970 1768.600 1273.290 ;
        RECT 1767.880 1207.350 1768.140 1207.670 ;
        RECT 1767.940 1173.670 1768.080 1207.350 ;
        RECT 1767.880 1173.350 1768.140 1173.670 ;
        RECT 1767.880 1172.670 1768.140 1172.990 ;
        RECT 1767.940 1087.050 1768.080 1172.670 ;
        RECT 1767.940 1086.910 1768.540 1087.050 ;
        RECT 1768.400 1062.830 1768.540 1086.910 ;
        RECT 1767.420 1062.510 1767.680 1062.830 ;
        RECT 1768.340 1062.510 1768.600 1062.830 ;
        RECT 1767.480 1028.490 1767.620 1062.510 ;
        RECT 1767.420 1028.170 1767.680 1028.490 ;
        RECT 1767.880 1027.830 1768.140 1028.150 ;
        RECT 1767.940 990.490 1768.080 1027.830 ;
        RECT 1767.940 990.350 1768.540 990.490 ;
        RECT 1768.400 966.270 1768.540 990.350 ;
        RECT 1767.420 966.125 1767.680 966.270 ;
        RECT 1768.340 966.125 1768.600 966.270 ;
        RECT 1767.410 965.755 1767.690 966.125 ;
        RECT 1768.330 965.755 1768.610 966.125 ;
        RECT 1768.400 931.330 1768.540 965.755 ;
        RECT 1767.940 931.190 1768.540 931.330 ;
        RECT 1767.940 893.930 1768.080 931.190 ;
        RECT 1767.940 893.790 1768.540 893.930 ;
        RECT 1768.400 869.710 1768.540 893.790 ;
        RECT 1767.420 869.565 1767.680 869.710 ;
        RECT 1767.410 869.195 1767.690 869.565 ;
        RECT 1768.340 869.390 1768.600 869.710 ;
        RECT 1767.870 868.515 1768.150 868.885 ;
        RECT 1767.940 821.090 1768.080 868.515 ;
        RECT 1767.420 820.770 1767.680 821.090 ;
        RECT 1767.880 820.770 1768.140 821.090 ;
        RECT 1767.480 814.290 1767.620 820.770 ;
        RECT 1767.420 813.970 1767.680 814.290 ;
        RECT 1767.420 766.030 1767.680 766.350 ;
        RECT 1767.480 765.670 1767.620 766.030 ;
        RECT 1767.420 765.350 1767.680 765.670 ;
        RECT 1767.420 723.870 1767.680 724.190 ;
        RECT 1767.480 651.850 1767.620 723.870 ;
        RECT 1767.480 651.710 1768.540 651.850 ;
        RECT 1768.400 641.650 1768.540 651.710 ;
        RECT 1767.940 641.510 1768.540 641.650 ;
        RECT 1767.940 580.030 1768.080 641.510 ;
        RECT 1767.880 579.710 1768.140 580.030 ;
        RECT 1767.880 572.570 1768.140 572.890 ;
        RECT 1767.940 531.410 1768.080 572.570 ;
        RECT 1767.420 531.090 1767.680 531.410 ;
        RECT 1767.880 531.090 1768.140 531.410 ;
        RECT 1767.480 524.270 1767.620 531.090 ;
        RECT 1767.420 523.950 1767.680 524.270 ;
        RECT 1767.420 476.010 1767.680 476.330 ;
        RECT 1767.480 458.730 1767.620 476.010 ;
        RECT 1767.480 458.590 1768.080 458.730 ;
        RECT 1767.940 434.850 1768.080 458.590 ;
        RECT 1767.420 434.530 1767.680 434.850 ;
        RECT 1767.880 434.530 1768.140 434.850 ;
        RECT 1767.480 427.710 1767.620 434.530 ;
        RECT 1767.420 427.390 1767.680 427.710 ;
        RECT 1767.880 427.050 1768.140 427.370 ;
        RECT 1767.940 379.430 1768.080 427.050 ;
        RECT 1767.880 379.110 1768.140 379.430 ;
        RECT 1768.340 331.170 1768.600 331.490 ;
        RECT 1768.400 241.810 1768.540 331.170 ;
        RECT 1767.940 241.670 1768.540 241.810 ;
        RECT 1767.940 144.830 1768.080 241.670 ;
        RECT 1767.880 144.510 1768.140 144.830 ;
        RECT 1768.340 144.510 1768.600 144.830 ;
        RECT 1768.400 138.030 1768.540 144.510 ;
        RECT 1768.340 137.710 1768.600 138.030 ;
        RECT 1768.340 96.230 1768.600 96.550 ;
        RECT 1768.400 60.930 1768.540 96.230 ;
        RECT 1767.020 60.790 1768.540 60.930 ;
        RECT 1767.020 35.010 1767.160 60.790 ;
        RECT 1209.900 34.690 1210.160 35.010 ;
        RECT 1766.960 34.690 1767.220 35.010 ;
        RECT 1209.960 2.400 1210.100 34.690 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
      LAYER via2 ;
        RECT 1767.410 965.800 1767.690 966.080 ;
        RECT 1768.330 965.800 1768.610 966.080 ;
        RECT 1767.410 869.240 1767.690 869.520 ;
        RECT 1767.870 868.560 1768.150 868.840 ;
      LAYER met3 ;
        RECT 1767.385 966.090 1767.715 966.105 ;
        RECT 1768.305 966.090 1768.635 966.105 ;
        RECT 1767.385 965.790 1768.635 966.090 ;
        RECT 1767.385 965.775 1767.715 965.790 ;
        RECT 1768.305 965.775 1768.635 965.790 ;
        RECT 1767.385 869.530 1767.715 869.545 ;
        RECT 1767.385 869.215 1767.930 869.530 ;
        RECT 1767.630 868.865 1767.930 869.215 ;
        RECT 1767.630 868.550 1768.175 868.865 ;
        RECT 1767.845 868.535 1768.175 868.550 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 38.660 1228.130 38.720 ;
        RECT 1780.730 38.660 1781.050 38.720 ;
        RECT 1227.810 38.520 1781.050 38.660 ;
        RECT 1227.810 38.460 1228.130 38.520 ;
        RECT 1780.730 38.460 1781.050 38.520 ;
      LAYER via ;
        RECT 1227.840 38.460 1228.100 38.720 ;
        RECT 1780.760 38.460 1781.020 38.720 ;
      LAYER met2 ;
        RECT 1780.220 1700.410 1780.500 1702.400 ;
        RECT 1780.220 1700.270 1780.960 1700.410 ;
        RECT 1780.220 1700.000 1780.500 1700.270 ;
        RECT 1780.820 38.750 1780.960 1700.270 ;
        RECT 1227.840 38.430 1228.100 38.750 ;
        RECT 1780.760 38.430 1781.020 38.750 ;
        RECT 1227.900 2.400 1228.040 38.430 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1245.750 39.000 1246.070 39.060 ;
        RECT 1787.170 39.000 1787.490 39.060 ;
        RECT 1245.750 38.860 1787.490 39.000 ;
        RECT 1245.750 38.800 1246.070 38.860 ;
        RECT 1787.170 38.800 1787.490 38.860 ;
      LAYER via ;
        RECT 1245.780 38.800 1246.040 39.060 ;
        RECT 1787.200 38.800 1787.460 39.060 ;
      LAYER met2 ;
        RECT 1789.420 1700.410 1789.700 1702.400 ;
        RECT 1787.260 1700.270 1789.700 1700.410 ;
        RECT 1787.260 39.090 1787.400 1700.270 ;
        RECT 1789.420 1700.000 1789.700 1700.270 ;
        RECT 1245.780 38.770 1246.040 39.090 ;
        RECT 1787.200 38.770 1787.460 39.090 ;
        RECT 1245.840 2.400 1245.980 38.770 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1795.065 1594.005 1795.235 1608.115 ;
        RECT 1795.065 1256.385 1795.235 1304.155 ;
        RECT 1795.065 1220.685 1795.235 1255.875 ;
        RECT 1794.605 1041.845 1794.775 1063.095 ;
        RECT 1795.065 772.905 1795.235 786.675 ;
        RECT 1795.065 365.925 1795.235 414.035 ;
        RECT 1795.525 269.025 1795.695 317.475 ;
        RECT 1795.065 179.605 1795.235 227.715 ;
        RECT 1795.065 89.845 1795.235 137.955 ;
      LAYER mcon ;
        RECT 1795.065 1607.945 1795.235 1608.115 ;
        RECT 1795.065 1303.985 1795.235 1304.155 ;
        RECT 1795.065 1255.705 1795.235 1255.875 ;
        RECT 1794.605 1062.925 1794.775 1063.095 ;
        RECT 1795.065 786.505 1795.235 786.675 ;
        RECT 1795.065 413.865 1795.235 414.035 ;
        RECT 1795.525 317.305 1795.695 317.475 ;
        RECT 1795.065 227.545 1795.235 227.715 ;
        RECT 1795.065 137.785 1795.235 137.955 ;
      LAYER met1 ;
        RECT 1795.450 1659.440 1795.770 1659.500 ;
        RECT 1796.370 1659.440 1796.690 1659.500 ;
        RECT 1795.450 1659.300 1796.690 1659.440 ;
        RECT 1795.450 1659.240 1795.770 1659.300 ;
        RECT 1796.370 1659.240 1796.690 1659.300 ;
        RECT 1795.005 1608.100 1795.295 1608.145 ;
        RECT 1795.450 1608.100 1795.770 1608.160 ;
        RECT 1795.005 1607.960 1795.770 1608.100 ;
        RECT 1795.005 1607.915 1795.295 1607.960 ;
        RECT 1795.450 1607.900 1795.770 1607.960 ;
        RECT 1794.990 1594.160 1795.310 1594.220 ;
        RECT 1794.795 1594.020 1795.310 1594.160 ;
        RECT 1794.990 1593.960 1795.310 1594.020 ;
        RECT 1794.990 1400.700 1795.310 1400.760 ;
        RECT 1795.450 1400.700 1795.770 1400.760 ;
        RECT 1794.990 1400.560 1795.770 1400.700 ;
        RECT 1794.990 1400.500 1795.310 1400.560 ;
        RECT 1795.450 1400.500 1795.770 1400.560 ;
        RECT 1794.530 1317.740 1794.850 1317.800 ;
        RECT 1794.530 1317.600 1795.680 1317.740 ;
        RECT 1794.530 1317.540 1794.850 1317.600 ;
        RECT 1795.540 1317.460 1795.680 1317.600 ;
        RECT 1795.450 1317.200 1795.770 1317.460 ;
        RECT 1795.005 1304.140 1795.295 1304.185 ;
        RECT 1795.450 1304.140 1795.770 1304.200 ;
        RECT 1795.005 1304.000 1795.770 1304.140 ;
        RECT 1795.005 1303.955 1795.295 1304.000 ;
        RECT 1795.450 1303.940 1795.770 1304.000 ;
        RECT 1794.990 1256.540 1795.310 1256.600 ;
        RECT 1794.795 1256.400 1795.310 1256.540 ;
        RECT 1794.990 1256.340 1795.310 1256.400 ;
        RECT 1794.990 1255.860 1795.310 1255.920 ;
        RECT 1794.795 1255.720 1795.310 1255.860 ;
        RECT 1794.990 1255.660 1795.310 1255.720 ;
        RECT 1794.990 1220.840 1795.310 1220.900 ;
        RECT 1794.795 1220.700 1795.310 1220.840 ;
        RECT 1794.990 1220.640 1795.310 1220.700 ;
        RECT 1794.990 1159.980 1795.310 1160.040 ;
        RECT 1794.990 1159.840 1795.680 1159.980 ;
        RECT 1794.990 1159.780 1795.310 1159.840 ;
        RECT 1795.540 1159.360 1795.680 1159.840 ;
        RECT 1795.450 1159.100 1795.770 1159.360 ;
        RECT 1794.545 1063.080 1794.835 1063.125 ;
        RECT 1794.990 1063.080 1795.310 1063.140 ;
        RECT 1794.545 1062.940 1795.310 1063.080 ;
        RECT 1794.545 1062.895 1794.835 1062.940 ;
        RECT 1794.990 1062.880 1795.310 1062.940 ;
        RECT 1794.530 1042.000 1794.850 1042.060 ;
        RECT 1794.335 1041.860 1794.850 1042.000 ;
        RECT 1794.530 1041.800 1794.850 1041.860 ;
        RECT 1794.530 980.120 1794.850 980.180 ;
        RECT 1795.450 980.120 1795.770 980.180 ;
        RECT 1794.530 979.980 1795.770 980.120 ;
        RECT 1794.530 979.920 1794.850 979.980 ;
        RECT 1795.450 979.920 1795.770 979.980 ;
        RECT 1795.450 894.100 1795.770 894.160 ;
        RECT 1795.080 893.960 1795.770 894.100 ;
        RECT 1795.080 893.820 1795.220 893.960 ;
        RECT 1795.450 893.900 1795.770 893.960 ;
        RECT 1794.990 893.560 1795.310 893.820 ;
        RECT 1794.990 835.080 1795.310 835.340 ;
        RECT 1795.080 834.600 1795.220 835.080 ;
        RECT 1795.450 834.600 1795.770 834.660 ;
        RECT 1795.080 834.460 1795.770 834.600 ;
        RECT 1795.450 834.400 1795.770 834.460 ;
        RECT 1795.005 786.660 1795.295 786.705 ;
        RECT 1795.450 786.660 1795.770 786.720 ;
        RECT 1795.005 786.520 1795.770 786.660 ;
        RECT 1795.005 786.475 1795.295 786.520 ;
        RECT 1795.450 786.460 1795.770 786.520 ;
        RECT 1794.990 773.060 1795.310 773.120 ;
        RECT 1794.795 772.920 1795.310 773.060 ;
        RECT 1794.990 772.860 1795.310 772.920 ;
        RECT 1794.990 738.520 1795.310 738.780 ;
        RECT 1795.080 738.100 1795.220 738.520 ;
        RECT 1794.990 737.840 1795.310 738.100 ;
        RECT 1794.990 676.640 1795.310 676.900 ;
        RECT 1795.080 676.220 1795.220 676.640 ;
        RECT 1794.990 675.960 1795.310 676.220 ;
        RECT 1794.990 414.020 1795.310 414.080 ;
        RECT 1794.795 413.880 1795.310 414.020 ;
        RECT 1794.990 413.820 1795.310 413.880 ;
        RECT 1794.990 366.080 1795.310 366.140 ;
        RECT 1794.795 365.940 1795.310 366.080 ;
        RECT 1794.990 365.880 1795.310 365.940 ;
        RECT 1795.450 317.460 1795.770 317.520 ;
        RECT 1795.255 317.320 1795.770 317.460 ;
        RECT 1795.450 317.260 1795.770 317.320 ;
        RECT 1795.465 269.180 1795.755 269.225 ;
        RECT 1795.910 269.180 1796.230 269.240 ;
        RECT 1795.465 269.040 1796.230 269.180 ;
        RECT 1795.465 268.995 1795.755 269.040 ;
        RECT 1795.910 268.980 1796.230 269.040 ;
        RECT 1794.990 234.500 1795.310 234.560 ;
        RECT 1795.910 234.500 1796.230 234.560 ;
        RECT 1794.990 234.360 1796.230 234.500 ;
        RECT 1794.990 234.300 1795.310 234.360 ;
        RECT 1795.910 234.300 1796.230 234.360 ;
        RECT 1794.990 227.700 1795.310 227.760 ;
        RECT 1794.795 227.560 1795.310 227.700 ;
        RECT 1794.990 227.500 1795.310 227.560 ;
        RECT 1794.990 179.760 1795.310 179.820 ;
        RECT 1794.795 179.620 1795.310 179.760 ;
        RECT 1794.990 179.560 1795.310 179.620 ;
        RECT 1794.990 137.940 1795.310 138.000 ;
        RECT 1794.795 137.800 1795.310 137.940 ;
        RECT 1794.990 137.740 1795.310 137.800 ;
        RECT 1794.990 90.000 1795.310 90.060 ;
        RECT 1794.795 89.860 1795.310 90.000 ;
        RECT 1794.990 89.800 1795.310 89.860 ;
        RECT 1263.230 39.340 1263.550 39.400 ;
        RECT 1794.990 39.340 1795.310 39.400 ;
        RECT 1263.230 39.200 1795.310 39.340 ;
        RECT 1263.230 39.140 1263.550 39.200 ;
        RECT 1794.990 39.140 1795.310 39.200 ;
      LAYER via ;
        RECT 1795.480 1659.240 1795.740 1659.500 ;
        RECT 1796.400 1659.240 1796.660 1659.500 ;
        RECT 1795.480 1607.900 1795.740 1608.160 ;
        RECT 1795.020 1593.960 1795.280 1594.220 ;
        RECT 1795.020 1400.500 1795.280 1400.760 ;
        RECT 1795.480 1400.500 1795.740 1400.760 ;
        RECT 1794.560 1317.540 1794.820 1317.800 ;
        RECT 1795.480 1317.200 1795.740 1317.460 ;
        RECT 1795.480 1303.940 1795.740 1304.200 ;
        RECT 1795.020 1256.340 1795.280 1256.600 ;
        RECT 1795.020 1255.660 1795.280 1255.920 ;
        RECT 1795.020 1220.640 1795.280 1220.900 ;
        RECT 1795.020 1159.780 1795.280 1160.040 ;
        RECT 1795.480 1159.100 1795.740 1159.360 ;
        RECT 1795.020 1062.880 1795.280 1063.140 ;
        RECT 1794.560 1041.800 1794.820 1042.060 ;
        RECT 1794.560 979.920 1794.820 980.180 ;
        RECT 1795.480 979.920 1795.740 980.180 ;
        RECT 1795.480 893.900 1795.740 894.160 ;
        RECT 1795.020 893.560 1795.280 893.820 ;
        RECT 1795.020 835.080 1795.280 835.340 ;
        RECT 1795.480 834.400 1795.740 834.660 ;
        RECT 1795.480 786.460 1795.740 786.720 ;
        RECT 1795.020 772.860 1795.280 773.120 ;
        RECT 1795.020 738.520 1795.280 738.780 ;
        RECT 1795.020 737.840 1795.280 738.100 ;
        RECT 1795.020 676.640 1795.280 676.900 ;
        RECT 1795.020 675.960 1795.280 676.220 ;
        RECT 1795.020 413.820 1795.280 414.080 ;
        RECT 1795.020 365.880 1795.280 366.140 ;
        RECT 1795.480 317.260 1795.740 317.520 ;
        RECT 1795.940 268.980 1796.200 269.240 ;
        RECT 1795.020 234.300 1795.280 234.560 ;
        RECT 1795.940 234.300 1796.200 234.560 ;
        RECT 1795.020 227.500 1795.280 227.760 ;
        RECT 1795.020 179.560 1795.280 179.820 ;
        RECT 1795.020 137.740 1795.280 138.000 ;
        RECT 1795.020 89.800 1795.280 90.060 ;
        RECT 1263.260 39.140 1263.520 39.400 ;
        RECT 1795.020 39.140 1795.280 39.400 ;
      LAYER met2 ;
        RECT 1798.620 1700.410 1798.900 1702.400 ;
        RECT 1796.460 1700.270 1798.900 1700.410 ;
        RECT 1796.460 1659.530 1796.600 1700.270 ;
        RECT 1798.620 1700.000 1798.900 1700.270 ;
        RECT 1795.480 1659.210 1795.740 1659.530 ;
        RECT 1796.400 1659.210 1796.660 1659.530 ;
        RECT 1795.540 1608.190 1795.680 1659.210 ;
        RECT 1795.480 1607.870 1795.740 1608.190 ;
        RECT 1795.020 1593.930 1795.280 1594.250 ;
        RECT 1795.080 1593.650 1795.220 1593.930 ;
        RECT 1795.080 1593.510 1795.680 1593.650 ;
        RECT 1795.540 1463.090 1795.680 1593.510 ;
        RECT 1795.080 1462.950 1795.680 1463.090 ;
        RECT 1795.080 1425.010 1795.220 1462.950 ;
        RECT 1794.620 1424.870 1795.220 1425.010 ;
        RECT 1794.620 1414.130 1794.760 1424.870 ;
        RECT 1794.620 1413.990 1795.680 1414.130 ;
        RECT 1795.540 1400.790 1795.680 1413.990 ;
        RECT 1795.020 1400.470 1795.280 1400.790 ;
        RECT 1795.480 1400.470 1795.740 1400.790 ;
        RECT 1795.080 1353.725 1795.220 1400.470 ;
        RECT 1795.010 1353.355 1795.290 1353.725 ;
        RECT 1794.550 1351.995 1794.830 1352.365 ;
        RECT 1794.620 1317.830 1794.760 1351.995 ;
        RECT 1794.560 1317.510 1794.820 1317.830 ;
        RECT 1795.480 1317.170 1795.740 1317.490 ;
        RECT 1795.540 1304.230 1795.680 1317.170 ;
        RECT 1795.480 1303.910 1795.740 1304.230 ;
        RECT 1795.020 1256.310 1795.280 1256.630 ;
        RECT 1795.080 1255.950 1795.220 1256.310 ;
        RECT 1795.020 1255.630 1795.280 1255.950 ;
        RECT 1795.020 1220.610 1795.280 1220.930 ;
        RECT 1795.080 1160.070 1795.220 1220.610 ;
        RECT 1795.020 1159.750 1795.280 1160.070 ;
        RECT 1795.480 1159.070 1795.740 1159.390 ;
        RECT 1795.540 1134.650 1795.680 1159.070 ;
        RECT 1795.080 1134.510 1795.680 1134.650 ;
        RECT 1795.080 1063.170 1795.220 1134.510 ;
        RECT 1795.020 1062.850 1795.280 1063.170 ;
        RECT 1794.560 1041.770 1794.820 1042.090 ;
        RECT 1794.620 1000.805 1794.760 1041.770 ;
        RECT 1794.550 1000.435 1794.830 1000.805 ;
        RECT 1795.470 1000.435 1795.750 1000.805 ;
        RECT 1795.540 980.210 1795.680 1000.435 ;
        RECT 1794.560 979.890 1794.820 980.210 ;
        RECT 1795.480 979.890 1795.740 980.210 ;
        RECT 1794.620 952.525 1794.760 979.890 ;
        RECT 1794.550 952.155 1794.830 952.525 ;
        RECT 1795.930 952.155 1796.210 952.525 ;
        RECT 1796.000 949.010 1796.140 952.155 ;
        RECT 1795.540 948.870 1796.140 949.010 ;
        RECT 1795.540 894.190 1795.680 948.870 ;
        RECT 1795.480 893.870 1795.740 894.190 ;
        RECT 1795.020 893.530 1795.280 893.850 ;
        RECT 1795.080 835.370 1795.220 893.530 ;
        RECT 1795.020 835.050 1795.280 835.370 ;
        RECT 1795.480 834.370 1795.740 834.690 ;
        RECT 1795.540 786.750 1795.680 834.370 ;
        RECT 1795.480 786.430 1795.740 786.750 ;
        RECT 1795.020 772.830 1795.280 773.150 ;
        RECT 1795.080 738.810 1795.220 772.830 ;
        RECT 1795.020 738.490 1795.280 738.810 ;
        RECT 1795.020 737.810 1795.280 738.130 ;
        RECT 1795.080 676.930 1795.220 737.810 ;
        RECT 1795.020 676.610 1795.280 676.930 ;
        RECT 1795.020 675.930 1795.280 676.250 ;
        RECT 1795.080 669.530 1795.220 675.930 ;
        RECT 1795.080 669.390 1795.680 669.530 ;
        RECT 1795.540 579.770 1795.680 669.390 ;
        RECT 1795.080 579.630 1795.680 579.770 ;
        RECT 1795.080 531.490 1795.220 579.630 ;
        RECT 1795.080 531.350 1795.680 531.490 ;
        RECT 1795.540 483.210 1795.680 531.350 ;
        RECT 1795.080 483.070 1795.680 483.210 ;
        RECT 1795.080 422.010 1795.220 483.070 ;
        RECT 1795.080 421.870 1795.680 422.010 ;
        RECT 1795.540 421.330 1795.680 421.870 ;
        RECT 1795.080 421.190 1795.680 421.330 ;
        RECT 1795.080 414.110 1795.220 421.190 ;
        RECT 1795.020 413.790 1795.280 414.110 ;
        RECT 1795.020 365.850 1795.280 366.170 ;
        RECT 1795.080 351.970 1795.220 365.850 ;
        RECT 1794.620 351.830 1795.220 351.970 ;
        RECT 1794.620 324.770 1794.760 351.830 ;
        RECT 1794.620 324.630 1795.680 324.770 ;
        RECT 1795.540 317.550 1795.680 324.630 ;
        RECT 1795.480 317.230 1795.740 317.550 ;
        RECT 1795.940 268.950 1796.200 269.270 ;
        RECT 1796.000 234.590 1796.140 268.950 ;
        RECT 1795.020 234.270 1795.280 234.590 ;
        RECT 1795.940 234.270 1796.200 234.590 ;
        RECT 1795.080 227.790 1795.220 234.270 ;
        RECT 1795.020 227.470 1795.280 227.790 ;
        RECT 1795.020 179.530 1795.280 179.850 ;
        RECT 1795.080 138.030 1795.220 179.530 ;
        RECT 1795.020 137.710 1795.280 138.030 ;
        RECT 1795.020 89.770 1795.280 90.090 ;
        RECT 1795.080 62.290 1795.220 89.770 ;
        RECT 1795.080 62.150 1795.680 62.290 ;
        RECT 1795.540 61.610 1795.680 62.150 ;
        RECT 1794.620 61.470 1795.680 61.610 ;
        RECT 1794.620 48.010 1794.760 61.470 ;
        RECT 1794.620 47.870 1795.220 48.010 ;
        RECT 1795.080 39.430 1795.220 47.870 ;
        RECT 1263.260 39.110 1263.520 39.430 ;
        RECT 1795.020 39.110 1795.280 39.430 ;
        RECT 1263.320 2.400 1263.460 39.110 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
      LAYER via2 ;
        RECT 1795.010 1353.400 1795.290 1353.680 ;
        RECT 1794.550 1352.040 1794.830 1352.320 ;
        RECT 1794.550 1000.480 1794.830 1000.760 ;
        RECT 1795.470 1000.480 1795.750 1000.760 ;
        RECT 1794.550 952.200 1794.830 952.480 ;
        RECT 1795.930 952.200 1796.210 952.480 ;
      LAYER met3 ;
        RECT 1794.985 1353.690 1795.315 1353.705 ;
        RECT 1794.310 1353.390 1795.315 1353.690 ;
        RECT 1794.310 1352.345 1794.610 1353.390 ;
        RECT 1794.985 1353.375 1795.315 1353.390 ;
        RECT 1794.310 1352.030 1794.855 1352.345 ;
        RECT 1794.525 1352.015 1794.855 1352.030 ;
        RECT 1794.525 1000.770 1794.855 1000.785 ;
        RECT 1795.445 1000.770 1795.775 1000.785 ;
        RECT 1794.525 1000.470 1795.775 1000.770 ;
        RECT 1794.525 1000.455 1794.855 1000.470 ;
        RECT 1795.445 1000.455 1795.775 1000.470 ;
        RECT 1794.525 952.490 1794.855 952.505 ;
        RECT 1795.905 952.490 1796.235 952.505 ;
        RECT 1794.525 952.190 1796.235 952.490 ;
        RECT 1794.525 952.175 1794.855 952.190 ;
        RECT 1795.905 952.175 1796.235 952.190 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1281.170 39.680 1281.490 39.740 ;
        RECT 1807.870 39.680 1808.190 39.740 ;
        RECT 1281.170 39.540 1808.190 39.680 ;
        RECT 1281.170 39.480 1281.490 39.540 ;
        RECT 1807.870 39.480 1808.190 39.540 ;
      LAYER via ;
        RECT 1281.200 39.480 1281.460 39.740 ;
        RECT 1807.900 39.480 1808.160 39.740 ;
      LAYER met2 ;
        RECT 1807.820 1700.000 1808.100 1702.400 ;
        RECT 1807.960 39.770 1808.100 1700.000 ;
        RECT 1281.200 39.450 1281.460 39.770 ;
        RECT 1807.900 39.450 1808.160 39.770 ;
        RECT 1281.260 2.400 1281.400 39.450 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1299.110 40.020 1299.430 40.080 ;
        RECT 1815.230 40.020 1815.550 40.080 ;
        RECT 1299.110 39.880 1815.550 40.020 ;
        RECT 1299.110 39.820 1299.430 39.880 ;
        RECT 1815.230 39.820 1815.550 39.880 ;
      LAYER via ;
        RECT 1299.140 39.820 1299.400 40.080 ;
        RECT 1815.260 39.820 1815.520 40.080 ;
      LAYER met2 ;
        RECT 1817.020 1700.410 1817.300 1702.400 ;
        RECT 1815.320 1700.270 1817.300 1700.410 ;
        RECT 1815.320 40.110 1815.460 1700.270 ;
        RECT 1817.020 1700.000 1817.300 1700.270 ;
        RECT 1299.140 39.790 1299.400 40.110 ;
        RECT 1815.260 39.790 1815.520 40.110 ;
        RECT 1299.200 2.400 1299.340 39.790 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1822.665 1365.865 1822.835 1400.715 ;
        RECT 1822.205 1090.125 1822.375 1179.715 ;
        RECT 1822.665 772.905 1822.835 838.355 ;
        RECT 1822.665 579.785 1822.835 627.895 ;
        RECT 1822.665 386.325 1822.835 434.435 ;
      LAYER mcon ;
        RECT 1822.665 1400.545 1822.835 1400.715 ;
        RECT 1822.205 1179.545 1822.375 1179.715 ;
        RECT 1822.665 838.185 1822.835 838.355 ;
        RECT 1822.665 627.725 1822.835 627.895 ;
        RECT 1822.665 434.265 1822.835 434.435 ;
      LAYER met1 ;
        RECT 1822.590 1657.060 1822.910 1657.120 ;
        RECT 1824.890 1657.060 1825.210 1657.120 ;
        RECT 1822.590 1656.920 1825.210 1657.060 ;
        RECT 1822.590 1656.860 1822.910 1656.920 ;
        RECT 1824.890 1656.860 1825.210 1656.920 ;
        RECT 1822.590 1414.440 1822.910 1414.700 ;
        RECT 1822.680 1413.960 1822.820 1414.440 ;
        RECT 1823.050 1413.960 1823.370 1414.020 ;
        RECT 1822.680 1413.820 1823.370 1413.960 ;
        RECT 1823.050 1413.760 1823.370 1413.820 ;
        RECT 1822.605 1400.700 1822.895 1400.745 ;
        RECT 1823.050 1400.700 1823.370 1400.760 ;
        RECT 1822.605 1400.560 1823.370 1400.700 ;
        RECT 1822.605 1400.515 1822.895 1400.560 ;
        RECT 1823.050 1400.500 1823.370 1400.560 ;
        RECT 1822.590 1366.020 1822.910 1366.080 ;
        RECT 1822.395 1365.880 1822.910 1366.020 ;
        RECT 1822.590 1365.820 1822.910 1365.880 ;
        RECT 1822.590 1317.880 1822.910 1318.140 ;
        RECT 1822.680 1317.400 1822.820 1317.880 ;
        RECT 1823.050 1317.400 1823.370 1317.460 ;
        RECT 1822.680 1317.260 1823.370 1317.400 ;
        RECT 1823.050 1317.200 1823.370 1317.260 ;
        RECT 1821.210 1304.140 1821.530 1304.200 ;
        RECT 1823.050 1304.140 1823.370 1304.200 ;
        RECT 1821.210 1304.000 1823.370 1304.140 ;
        RECT 1821.210 1303.940 1821.530 1304.000 ;
        RECT 1823.050 1303.940 1823.370 1304.000 ;
        RECT 1821.210 1210.980 1821.530 1211.040 ;
        RECT 1823.050 1210.980 1823.370 1211.040 ;
        RECT 1821.210 1210.840 1823.370 1210.980 ;
        RECT 1821.210 1210.780 1821.530 1210.840 ;
        RECT 1823.050 1210.780 1823.370 1210.840 ;
        RECT 1822.145 1179.700 1822.435 1179.745 ;
        RECT 1823.050 1179.700 1823.370 1179.760 ;
        RECT 1822.145 1179.560 1823.370 1179.700 ;
        RECT 1822.145 1179.515 1822.435 1179.560 ;
        RECT 1823.050 1179.500 1823.370 1179.560 ;
        RECT 1822.130 1090.280 1822.450 1090.340 ;
        RECT 1821.935 1090.140 1822.450 1090.280 ;
        RECT 1822.130 1090.080 1822.450 1090.140 ;
        RECT 1823.050 980.260 1823.370 980.520 ;
        RECT 1823.140 979.840 1823.280 980.260 ;
        RECT 1823.050 979.580 1823.370 979.840 ;
        RECT 1822.590 838.340 1822.910 838.400 ;
        RECT 1822.395 838.200 1822.910 838.340 ;
        RECT 1822.590 838.140 1822.910 838.200 ;
        RECT 1822.605 773.060 1822.895 773.105 ;
        RECT 1823.050 773.060 1823.370 773.120 ;
        RECT 1822.605 772.920 1823.370 773.060 ;
        RECT 1822.605 772.875 1822.895 772.920 ;
        RECT 1823.050 772.860 1823.370 772.920 ;
        RECT 1823.050 724.440 1823.370 724.500 ;
        RECT 1823.510 724.440 1823.830 724.500 ;
        RECT 1823.050 724.300 1823.830 724.440 ;
        RECT 1823.050 724.240 1823.370 724.300 ;
        RECT 1823.510 724.240 1823.830 724.300 ;
        RECT 1822.605 627.880 1822.895 627.925 ;
        RECT 1823.050 627.880 1823.370 627.940 ;
        RECT 1822.605 627.740 1823.370 627.880 ;
        RECT 1822.605 627.695 1822.895 627.740 ;
        RECT 1823.050 627.680 1823.370 627.740 ;
        RECT 1822.590 579.940 1822.910 580.000 ;
        RECT 1822.395 579.800 1822.910 579.940 ;
        RECT 1822.590 579.740 1822.910 579.800 ;
        RECT 1822.590 531.320 1822.910 531.380 ;
        RECT 1823.050 531.320 1823.370 531.380 ;
        RECT 1822.590 531.180 1823.370 531.320 ;
        RECT 1822.590 531.120 1822.910 531.180 ;
        RECT 1823.050 531.120 1823.370 531.180 ;
        RECT 1822.590 434.420 1822.910 434.480 ;
        RECT 1822.395 434.280 1822.910 434.420 ;
        RECT 1822.590 434.220 1822.910 434.280 ;
        RECT 1822.590 386.480 1822.910 386.540 ;
        RECT 1822.395 386.340 1822.910 386.480 ;
        RECT 1822.590 386.280 1822.910 386.340 ;
        RECT 1822.590 110.540 1822.910 110.800 ;
        RECT 1822.680 110.120 1822.820 110.540 ;
        RECT 1822.590 109.860 1822.910 110.120 ;
        RECT 1317.050 40.360 1317.370 40.420 ;
        RECT 1822.590 40.360 1822.910 40.420 ;
        RECT 1317.050 40.220 1822.910 40.360 ;
        RECT 1317.050 40.160 1317.370 40.220 ;
        RECT 1822.590 40.160 1822.910 40.220 ;
      LAYER via ;
        RECT 1822.620 1656.860 1822.880 1657.120 ;
        RECT 1824.920 1656.860 1825.180 1657.120 ;
        RECT 1822.620 1414.440 1822.880 1414.700 ;
        RECT 1823.080 1413.760 1823.340 1414.020 ;
        RECT 1823.080 1400.500 1823.340 1400.760 ;
        RECT 1822.620 1365.820 1822.880 1366.080 ;
        RECT 1822.620 1317.880 1822.880 1318.140 ;
        RECT 1823.080 1317.200 1823.340 1317.460 ;
        RECT 1821.240 1303.940 1821.500 1304.200 ;
        RECT 1823.080 1303.940 1823.340 1304.200 ;
        RECT 1821.240 1210.780 1821.500 1211.040 ;
        RECT 1823.080 1210.780 1823.340 1211.040 ;
        RECT 1823.080 1179.500 1823.340 1179.760 ;
        RECT 1822.160 1090.080 1822.420 1090.340 ;
        RECT 1823.080 980.260 1823.340 980.520 ;
        RECT 1823.080 979.580 1823.340 979.840 ;
        RECT 1822.620 838.140 1822.880 838.400 ;
        RECT 1823.080 772.860 1823.340 773.120 ;
        RECT 1823.080 724.240 1823.340 724.500 ;
        RECT 1823.540 724.240 1823.800 724.500 ;
        RECT 1823.080 627.680 1823.340 627.940 ;
        RECT 1822.620 579.740 1822.880 580.000 ;
        RECT 1822.620 531.120 1822.880 531.380 ;
        RECT 1823.080 531.120 1823.340 531.380 ;
        RECT 1822.620 434.220 1822.880 434.480 ;
        RECT 1822.620 386.280 1822.880 386.540 ;
        RECT 1822.620 110.540 1822.880 110.800 ;
        RECT 1822.620 109.860 1822.880 110.120 ;
        RECT 1317.080 40.160 1317.340 40.420 ;
        RECT 1822.620 40.160 1822.880 40.420 ;
      LAYER met2 ;
        RECT 1826.220 1700.410 1826.500 1702.400 ;
        RECT 1824.980 1700.270 1826.500 1700.410 ;
        RECT 1824.980 1657.150 1825.120 1700.270 ;
        RECT 1826.220 1700.000 1826.500 1700.270 ;
        RECT 1822.620 1656.830 1822.880 1657.150 ;
        RECT 1824.920 1656.830 1825.180 1657.150 ;
        RECT 1822.680 1655.530 1822.820 1656.830 ;
        RECT 1822.680 1655.390 1823.280 1655.530 ;
        RECT 1823.140 1606.570 1823.280 1655.390 ;
        RECT 1822.680 1606.430 1823.280 1606.570 ;
        RECT 1822.680 1593.650 1822.820 1606.430 ;
        RECT 1822.680 1593.510 1823.280 1593.650 ;
        RECT 1823.140 1463.090 1823.280 1593.510 ;
        RECT 1822.680 1462.950 1823.280 1463.090 ;
        RECT 1822.680 1414.730 1822.820 1462.950 ;
        RECT 1822.620 1414.410 1822.880 1414.730 ;
        RECT 1823.080 1413.730 1823.340 1414.050 ;
        RECT 1823.140 1400.790 1823.280 1413.730 ;
        RECT 1823.080 1400.470 1823.340 1400.790 ;
        RECT 1822.620 1365.790 1822.880 1366.110 ;
        RECT 1822.680 1318.170 1822.820 1365.790 ;
        RECT 1822.620 1317.850 1822.880 1318.170 ;
        RECT 1823.080 1317.170 1823.340 1317.490 ;
        RECT 1823.140 1304.230 1823.280 1317.170 ;
        RECT 1821.240 1303.910 1821.500 1304.230 ;
        RECT 1823.080 1303.910 1823.340 1304.230 ;
        RECT 1821.300 1256.485 1821.440 1303.910 ;
        RECT 1821.230 1256.115 1821.510 1256.485 ;
        RECT 1821.230 1255.435 1821.510 1255.805 ;
        RECT 1821.300 1211.070 1821.440 1255.435 ;
        RECT 1821.240 1210.750 1821.500 1211.070 ;
        RECT 1823.080 1210.750 1823.340 1211.070 ;
        RECT 1823.140 1179.790 1823.280 1210.750 ;
        RECT 1823.080 1179.470 1823.340 1179.790 ;
        RECT 1822.160 1090.050 1822.420 1090.370 ;
        RECT 1822.220 1089.885 1822.360 1090.050 ;
        RECT 1822.150 1089.515 1822.430 1089.885 ;
        RECT 1823.070 1089.515 1823.350 1089.885 ;
        RECT 1823.140 1061.890 1823.280 1089.515 ;
        RECT 1822.220 1061.750 1823.280 1061.890 ;
        RECT 1822.220 1000.805 1822.360 1061.750 ;
        RECT 1822.150 1000.435 1822.430 1000.805 ;
        RECT 1823.070 1000.435 1823.350 1000.805 ;
        RECT 1823.140 980.550 1823.280 1000.435 ;
        RECT 1823.080 980.230 1823.340 980.550 ;
        RECT 1823.080 979.550 1823.340 979.870 ;
        RECT 1823.140 952.525 1823.280 979.550 ;
        RECT 1823.070 952.155 1823.350 952.525 ;
        RECT 1823.990 952.155 1824.270 952.525 ;
        RECT 1824.060 917.050 1824.200 952.155 ;
        RECT 1823.600 916.910 1824.200 917.050 ;
        RECT 1823.600 862.765 1823.740 916.910 ;
        RECT 1822.610 862.395 1822.890 862.765 ;
        RECT 1823.530 862.395 1823.810 862.765 ;
        RECT 1822.680 838.430 1822.820 862.395 ;
        RECT 1822.620 838.110 1822.880 838.430 ;
        RECT 1823.080 772.890 1823.340 773.150 ;
        RECT 1822.680 772.830 1823.340 772.890 ;
        RECT 1822.680 772.750 1823.280 772.830 ;
        RECT 1822.680 759.970 1822.820 772.750 ;
        RECT 1822.680 759.830 1823.740 759.970 ;
        RECT 1823.600 737.530 1823.740 759.830 ;
        RECT 1823.140 737.390 1823.740 737.530 ;
        RECT 1823.140 724.530 1823.280 737.390 ;
        RECT 1823.080 724.210 1823.340 724.530 ;
        RECT 1823.540 724.210 1823.800 724.530 ;
        RECT 1823.600 676.445 1823.740 724.210 ;
        RECT 1822.610 676.075 1822.890 676.445 ;
        RECT 1823.530 676.075 1823.810 676.445 ;
        RECT 1822.680 651.850 1822.820 676.075 ;
        RECT 1822.680 651.710 1823.280 651.850 ;
        RECT 1823.140 627.970 1823.280 651.710 ;
        RECT 1823.080 627.650 1823.340 627.970 ;
        RECT 1822.620 579.710 1822.880 580.030 ;
        RECT 1822.680 555.290 1822.820 579.710 ;
        RECT 1822.220 555.150 1822.820 555.290 ;
        RECT 1822.220 544.410 1822.360 555.150 ;
        RECT 1822.220 544.270 1823.280 544.410 ;
        RECT 1823.140 531.410 1823.280 544.270 ;
        RECT 1822.620 531.090 1822.880 531.410 ;
        RECT 1823.080 531.090 1823.340 531.410 ;
        RECT 1822.680 434.510 1822.820 531.090 ;
        RECT 1822.620 434.190 1822.880 434.510 ;
        RECT 1822.620 386.250 1822.880 386.570 ;
        RECT 1822.680 110.830 1822.820 386.250 ;
        RECT 1822.620 110.510 1822.880 110.830 ;
        RECT 1822.620 109.830 1822.880 110.150 ;
        RECT 1822.680 40.450 1822.820 109.830 ;
        RECT 1317.080 40.130 1317.340 40.450 ;
        RECT 1822.620 40.130 1822.880 40.450 ;
        RECT 1317.140 2.400 1317.280 40.130 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
      LAYER via2 ;
        RECT 1821.230 1256.160 1821.510 1256.440 ;
        RECT 1821.230 1255.480 1821.510 1255.760 ;
        RECT 1822.150 1089.560 1822.430 1089.840 ;
        RECT 1823.070 1089.560 1823.350 1089.840 ;
        RECT 1822.150 1000.480 1822.430 1000.760 ;
        RECT 1823.070 1000.480 1823.350 1000.760 ;
        RECT 1823.070 952.200 1823.350 952.480 ;
        RECT 1823.990 952.200 1824.270 952.480 ;
        RECT 1822.610 862.440 1822.890 862.720 ;
        RECT 1823.530 862.440 1823.810 862.720 ;
        RECT 1822.610 676.120 1822.890 676.400 ;
        RECT 1823.530 676.120 1823.810 676.400 ;
      LAYER met3 ;
        RECT 1821.205 1256.450 1821.535 1256.465 ;
        RECT 1821.205 1256.150 1822.210 1256.450 ;
        RECT 1821.205 1256.135 1821.535 1256.150 ;
        RECT 1821.205 1255.770 1821.535 1255.785 ;
        RECT 1821.910 1255.770 1822.210 1256.150 ;
        RECT 1821.205 1255.470 1822.210 1255.770 ;
        RECT 1821.205 1255.455 1821.535 1255.470 ;
        RECT 1822.125 1089.850 1822.455 1089.865 ;
        RECT 1823.045 1089.850 1823.375 1089.865 ;
        RECT 1822.125 1089.550 1823.375 1089.850 ;
        RECT 1822.125 1089.535 1822.455 1089.550 ;
        RECT 1823.045 1089.535 1823.375 1089.550 ;
        RECT 1822.125 1000.770 1822.455 1000.785 ;
        RECT 1823.045 1000.770 1823.375 1000.785 ;
        RECT 1822.125 1000.470 1823.375 1000.770 ;
        RECT 1822.125 1000.455 1822.455 1000.470 ;
        RECT 1823.045 1000.455 1823.375 1000.470 ;
        RECT 1823.045 952.490 1823.375 952.505 ;
        RECT 1823.965 952.490 1824.295 952.505 ;
        RECT 1823.045 952.190 1824.295 952.490 ;
        RECT 1823.045 952.175 1823.375 952.190 ;
        RECT 1823.965 952.175 1824.295 952.190 ;
        RECT 1822.585 862.730 1822.915 862.745 ;
        RECT 1823.505 862.730 1823.835 862.745 ;
        RECT 1822.585 862.430 1823.835 862.730 ;
        RECT 1822.585 862.415 1822.915 862.430 ;
        RECT 1823.505 862.415 1823.835 862.430 ;
        RECT 1822.585 676.410 1822.915 676.425 ;
        RECT 1823.505 676.410 1823.835 676.425 ;
        RECT 1822.585 676.110 1823.835 676.410 ;
        RECT 1822.585 676.095 1822.915 676.110 ;
        RECT 1823.505 676.095 1823.835 676.110 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.990 40.700 1335.310 40.760 ;
        RECT 1835.470 40.700 1835.790 40.760 ;
        RECT 1334.990 40.560 1835.790 40.700 ;
        RECT 1334.990 40.500 1335.310 40.560 ;
        RECT 1835.470 40.500 1835.790 40.560 ;
      LAYER via ;
        RECT 1335.020 40.500 1335.280 40.760 ;
        RECT 1835.500 40.500 1835.760 40.760 ;
      LAYER met2 ;
        RECT 1835.420 1700.000 1835.700 1702.400 ;
        RECT 1835.560 40.790 1835.700 1700.000 ;
        RECT 1335.020 40.470 1335.280 40.790 ;
        RECT 1835.500 40.470 1835.760 40.790 ;
        RECT 1335.080 2.400 1335.220 40.470 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 692.370 36.620 692.690 36.680 ;
        RECT 1504.270 36.620 1504.590 36.680 ;
        RECT 692.370 36.480 1504.590 36.620 ;
        RECT 692.370 36.420 692.690 36.480 ;
        RECT 1504.270 36.420 1504.590 36.480 ;
      LAYER via ;
        RECT 692.400 36.420 692.660 36.680 ;
        RECT 1504.300 36.420 1504.560 36.680 ;
      LAYER met2 ;
        RECT 1504.680 1700.410 1504.960 1702.400 ;
        RECT 1504.360 1700.270 1504.960 1700.410 ;
        RECT 1504.360 36.710 1504.500 1700.270 ;
        RECT 1504.680 1700.000 1504.960 1700.270 ;
        RECT 692.400 36.390 692.660 36.710 ;
        RECT 1504.300 36.390 1504.560 36.710 ;
        RECT 692.460 2.400 692.600 36.390 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.470 41.040 1352.790 41.100 ;
        RECT 1842.830 41.040 1843.150 41.100 ;
        RECT 1352.470 40.900 1843.150 41.040 ;
        RECT 1352.470 40.840 1352.790 40.900 ;
        RECT 1842.830 40.840 1843.150 40.900 ;
      LAYER via ;
        RECT 1352.500 40.840 1352.760 41.100 ;
        RECT 1842.860 40.840 1843.120 41.100 ;
      LAYER met2 ;
        RECT 1844.620 1700.410 1844.900 1702.400 ;
        RECT 1842.920 1700.270 1844.900 1700.410 ;
        RECT 1842.920 41.130 1843.060 1700.270 ;
        RECT 1844.620 1700.000 1844.900 1700.270 ;
        RECT 1352.500 40.810 1352.760 41.130 ;
        RECT 1842.860 40.810 1843.120 41.130 ;
        RECT 1352.560 2.400 1352.700 40.810 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1850.265 1635.485 1850.435 1683.595 ;
        RECT 1850.725 1448.485 1850.895 1490.475 ;
        RECT 1849.805 1207.425 1849.975 1255.875 ;
        RECT 1850.265 737.885 1850.435 772.735 ;
        RECT 1850.265 641.325 1850.435 676.175 ;
        RECT 1850.725 531.505 1850.895 545.275 ;
        RECT 1850.265 386.325 1850.435 434.435 ;
        RECT 1850.265 241.485 1850.435 305.575 ;
        RECT 1849.805 192.865 1849.975 207.315 ;
      LAYER mcon ;
        RECT 1850.265 1683.425 1850.435 1683.595 ;
        RECT 1850.725 1490.305 1850.895 1490.475 ;
        RECT 1849.805 1255.705 1849.975 1255.875 ;
        RECT 1850.265 772.565 1850.435 772.735 ;
        RECT 1850.265 676.005 1850.435 676.175 ;
        RECT 1850.725 545.105 1850.895 545.275 ;
        RECT 1850.265 434.265 1850.435 434.435 ;
        RECT 1850.265 305.405 1850.435 305.575 ;
        RECT 1849.805 207.145 1849.975 207.315 ;
      LAYER met1 ;
        RECT 1850.205 1683.580 1850.495 1683.625 ;
        RECT 1852.490 1683.580 1852.810 1683.640 ;
        RECT 1850.205 1683.440 1852.810 1683.580 ;
        RECT 1850.205 1683.395 1850.495 1683.440 ;
        RECT 1852.490 1683.380 1852.810 1683.440 ;
        RECT 1850.190 1635.640 1850.510 1635.700 ;
        RECT 1849.995 1635.500 1850.510 1635.640 ;
        RECT 1850.190 1635.440 1850.510 1635.500 ;
        RECT 1850.650 1497.600 1850.970 1497.660 ;
        RECT 1851.110 1497.600 1851.430 1497.660 ;
        RECT 1850.650 1497.460 1851.430 1497.600 ;
        RECT 1850.650 1497.400 1850.970 1497.460 ;
        RECT 1851.110 1497.400 1851.430 1497.460 ;
        RECT 1850.650 1490.460 1850.970 1490.520 ;
        RECT 1850.455 1490.320 1850.970 1490.460 ;
        RECT 1850.650 1490.260 1850.970 1490.320 ;
        RECT 1850.665 1448.640 1850.955 1448.685 ;
        RECT 1851.110 1448.640 1851.430 1448.700 ;
        RECT 1850.665 1448.500 1851.430 1448.640 ;
        RECT 1850.665 1448.455 1850.955 1448.500 ;
        RECT 1851.110 1448.440 1851.430 1448.500 ;
        RECT 1849.730 1400.700 1850.050 1400.760 ;
        RECT 1851.110 1400.700 1851.430 1400.760 ;
        RECT 1849.730 1400.560 1851.430 1400.700 ;
        RECT 1849.730 1400.500 1850.050 1400.560 ;
        RECT 1851.110 1400.500 1851.430 1400.560 ;
        RECT 1849.745 1255.860 1850.035 1255.905 ;
        RECT 1850.190 1255.860 1850.510 1255.920 ;
        RECT 1849.745 1255.720 1850.510 1255.860 ;
        RECT 1849.745 1255.675 1850.035 1255.720 ;
        RECT 1850.190 1255.660 1850.510 1255.720 ;
        RECT 1849.730 1207.580 1850.050 1207.640 ;
        RECT 1849.535 1207.440 1850.050 1207.580 ;
        RECT 1849.730 1207.380 1850.050 1207.440 ;
        RECT 1849.730 1159.300 1850.050 1159.360 ;
        RECT 1850.190 1159.300 1850.510 1159.360 ;
        RECT 1849.730 1159.160 1850.510 1159.300 ;
        RECT 1849.730 1159.100 1850.050 1159.160 ;
        RECT 1850.190 1159.100 1850.510 1159.160 ;
        RECT 1850.190 1076.820 1850.510 1077.080 ;
        RECT 1850.280 1076.400 1850.420 1076.820 ;
        RECT 1850.190 1076.140 1850.510 1076.400 ;
        RECT 1850.190 1055.600 1850.510 1055.660 ;
        RECT 1851.110 1055.600 1851.430 1055.660 ;
        RECT 1850.190 1055.460 1851.430 1055.600 ;
        RECT 1850.190 1055.400 1850.510 1055.460 ;
        RECT 1851.110 1055.400 1851.430 1055.460 ;
        RECT 1850.190 980.260 1850.510 980.520 ;
        RECT 1850.280 979.840 1850.420 980.260 ;
        RECT 1850.190 979.580 1850.510 979.840 ;
        RECT 1848.810 959.040 1849.130 959.100 ;
        RECT 1850.190 959.040 1850.510 959.100 ;
        RECT 1848.810 958.900 1850.510 959.040 ;
        RECT 1848.810 958.840 1849.130 958.900 ;
        RECT 1850.190 958.840 1850.510 958.900 ;
        RECT 1849.730 910.760 1850.050 910.820 ;
        RECT 1852.030 910.760 1852.350 910.820 ;
        RECT 1849.730 910.620 1852.350 910.760 ;
        RECT 1849.730 910.560 1850.050 910.620 ;
        RECT 1852.030 910.560 1852.350 910.620 ;
        RECT 1850.190 772.720 1850.510 772.780 ;
        RECT 1849.995 772.580 1850.510 772.720 ;
        RECT 1850.190 772.520 1850.510 772.580 ;
        RECT 1850.190 738.040 1850.510 738.100 ;
        RECT 1849.995 737.900 1850.510 738.040 ;
        RECT 1850.190 737.840 1850.510 737.900 ;
        RECT 1850.190 676.160 1850.510 676.220 ;
        RECT 1849.995 676.020 1850.510 676.160 ;
        RECT 1850.190 675.960 1850.510 676.020 ;
        RECT 1850.190 641.480 1850.510 641.540 ;
        RECT 1849.995 641.340 1850.510 641.480 ;
        RECT 1850.190 641.280 1850.510 641.340 ;
        RECT 1850.650 603.540 1850.970 603.800 ;
        RECT 1850.740 603.120 1850.880 603.540 ;
        RECT 1850.650 602.860 1850.970 603.120 ;
        RECT 1850.650 545.260 1850.970 545.320 ;
        RECT 1850.455 545.120 1850.970 545.260 ;
        RECT 1850.650 545.060 1850.970 545.120 ;
        RECT 1850.650 531.660 1850.970 531.720 ;
        RECT 1850.455 531.520 1850.970 531.660 ;
        RECT 1850.650 531.460 1850.970 531.520 ;
        RECT 1850.190 434.420 1850.510 434.480 ;
        RECT 1849.995 434.280 1850.510 434.420 ;
        RECT 1850.190 434.220 1850.510 434.280 ;
        RECT 1850.190 386.480 1850.510 386.540 ;
        RECT 1849.995 386.340 1850.510 386.480 ;
        RECT 1850.190 386.280 1850.510 386.340 ;
        RECT 1850.190 305.560 1850.510 305.620 ;
        RECT 1849.995 305.420 1850.510 305.560 ;
        RECT 1850.190 305.360 1850.510 305.420 ;
        RECT 1850.205 241.640 1850.495 241.685 ;
        RECT 1850.650 241.640 1850.970 241.700 ;
        RECT 1850.205 241.500 1850.970 241.640 ;
        RECT 1850.205 241.455 1850.495 241.500 ;
        RECT 1850.650 241.440 1850.970 241.500 ;
        RECT 1849.745 207.300 1850.035 207.345 ;
        RECT 1850.650 207.300 1850.970 207.360 ;
        RECT 1849.745 207.160 1850.970 207.300 ;
        RECT 1849.745 207.115 1850.035 207.160 ;
        RECT 1850.650 207.100 1850.970 207.160 ;
        RECT 1849.730 193.020 1850.050 193.080 ;
        RECT 1849.535 192.880 1850.050 193.020 ;
        RECT 1849.730 192.820 1850.050 192.880 ;
        RECT 1849.730 169.220 1850.050 169.280 ;
        RECT 1851.110 169.220 1851.430 169.280 ;
        RECT 1849.730 169.080 1851.430 169.220 ;
        RECT 1849.730 169.020 1850.050 169.080 ;
        RECT 1851.110 169.020 1851.430 169.080 ;
        RECT 1850.190 96.800 1850.510 96.860 ;
        RECT 1851.110 96.800 1851.430 96.860 ;
        RECT 1850.190 96.660 1851.430 96.800 ;
        RECT 1850.190 96.600 1850.510 96.660 ;
        RECT 1851.110 96.600 1851.430 96.660 ;
        RECT 1370.410 41.380 1370.730 41.440 ;
        RECT 1850.650 41.380 1850.970 41.440 ;
        RECT 1370.410 41.240 1850.970 41.380 ;
        RECT 1370.410 41.180 1370.730 41.240 ;
        RECT 1850.650 41.180 1850.970 41.240 ;
      LAYER via ;
        RECT 1852.520 1683.380 1852.780 1683.640 ;
        RECT 1850.220 1635.440 1850.480 1635.700 ;
        RECT 1850.680 1497.400 1850.940 1497.660 ;
        RECT 1851.140 1497.400 1851.400 1497.660 ;
        RECT 1850.680 1490.260 1850.940 1490.520 ;
        RECT 1851.140 1448.440 1851.400 1448.700 ;
        RECT 1849.760 1400.500 1850.020 1400.760 ;
        RECT 1851.140 1400.500 1851.400 1400.760 ;
        RECT 1850.220 1255.660 1850.480 1255.920 ;
        RECT 1849.760 1207.380 1850.020 1207.640 ;
        RECT 1849.760 1159.100 1850.020 1159.360 ;
        RECT 1850.220 1159.100 1850.480 1159.360 ;
        RECT 1850.220 1076.820 1850.480 1077.080 ;
        RECT 1850.220 1076.140 1850.480 1076.400 ;
        RECT 1850.220 1055.400 1850.480 1055.660 ;
        RECT 1851.140 1055.400 1851.400 1055.660 ;
        RECT 1850.220 980.260 1850.480 980.520 ;
        RECT 1850.220 979.580 1850.480 979.840 ;
        RECT 1848.840 958.840 1849.100 959.100 ;
        RECT 1850.220 958.840 1850.480 959.100 ;
        RECT 1849.760 910.560 1850.020 910.820 ;
        RECT 1852.060 910.560 1852.320 910.820 ;
        RECT 1850.220 772.520 1850.480 772.780 ;
        RECT 1850.220 737.840 1850.480 738.100 ;
        RECT 1850.220 675.960 1850.480 676.220 ;
        RECT 1850.220 641.280 1850.480 641.540 ;
        RECT 1850.680 603.540 1850.940 603.800 ;
        RECT 1850.680 602.860 1850.940 603.120 ;
        RECT 1850.680 545.060 1850.940 545.320 ;
        RECT 1850.680 531.460 1850.940 531.720 ;
        RECT 1850.220 434.220 1850.480 434.480 ;
        RECT 1850.220 386.280 1850.480 386.540 ;
        RECT 1850.220 305.360 1850.480 305.620 ;
        RECT 1850.680 241.440 1850.940 241.700 ;
        RECT 1850.680 207.100 1850.940 207.360 ;
        RECT 1849.760 192.820 1850.020 193.080 ;
        RECT 1849.760 169.020 1850.020 169.280 ;
        RECT 1851.140 169.020 1851.400 169.280 ;
        RECT 1850.220 96.600 1850.480 96.860 ;
        RECT 1851.140 96.600 1851.400 96.860 ;
        RECT 1370.440 41.180 1370.700 41.440 ;
        RECT 1850.680 41.180 1850.940 41.440 ;
      LAYER met2 ;
        RECT 1853.820 1700.410 1854.100 1702.400 ;
        RECT 1852.580 1700.270 1854.100 1700.410 ;
        RECT 1852.580 1683.670 1852.720 1700.270 ;
        RECT 1853.820 1700.000 1854.100 1700.270 ;
        RECT 1852.520 1683.350 1852.780 1683.670 ;
        RECT 1850.220 1635.410 1850.480 1635.730 ;
        RECT 1850.280 1587.530 1850.420 1635.410 ;
        RECT 1850.280 1587.390 1851.340 1587.530 ;
        RECT 1851.200 1497.690 1851.340 1587.390 ;
        RECT 1850.680 1497.370 1850.940 1497.690 ;
        RECT 1851.140 1497.370 1851.400 1497.690 ;
        RECT 1850.740 1490.550 1850.880 1497.370 ;
        RECT 1850.680 1490.230 1850.940 1490.550 ;
        RECT 1851.140 1448.410 1851.400 1448.730 ;
        RECT 1851.200 1400.790 1851.340 1448.410 ;
        RECT 1849.760 1400.470 1850.020 1400.790 ;
        RECT 1851.140 1400.470 1851.400 1400.790 ;
        RECT 1849.820 1393.845 1849.960 1400.470 ;
        RECT 1849.750 1393.475 1850.030 1393.845 ;
        RECT 1851.590 1393.475 1851.870 1393.845 ;
        RECT 1851.660 1269.290 1851.800 1393.475 ;
        RECT 1850.280 1269.150 1851.800 1269.290 ;
        RECT 1850.280 1255.950 1850.420 1269.150 ;
        RECT 1850.220 1255.630 1850.480 1255.950 ;
        RECT 1849.760 1207.350 1850.020 1207.670 ;
        RECT 1849.820 1159.390 1849.960 1207.350 ;
        RECT 1849.760 1159.070 1850.020 1159.390 ;
        RECT 1850.220 1159.070 1850.480 1159.390 ;
        RECT 1850.280 1077.110 1850.420 1159.070 ;
        RECT 1850.220 1076.790 1850.480 1077.110 ;
        RECT 1850.220 1076.110 1850.480 1076.430 ;
        RECT 1850.280 1055.690 1850.420 1076.110 ;
        RECT 1850.220 1055.370 1850.480 1055.690 ;
        RECT 1851.140 1055.370 1851.400 1055.690 ;
        RECT 1851.200 1007.605 1851.340 1055.370 ;
        RECT 1850.210 1007.235 1850.490 1007.605 ;
        RECT 1851.130 1007.235 1851.410 1007.605 ;
        RECT 1850.280 980.550 1850.420 1007.235 ;
        RECT 1850.220 980.230 1850.480 980.550 ;
        RECT 1850.220 979.550 1850.480 979.870 ;
        RECT 1850.280 959.130 1850.420 979.550 ;
        RECT 1848.840 958.810 1849.100 959.130 ;
        RECT 1850.220 958.810 1850.480 959.130 ;
        RECT 1848.900 911.045 1849.040 958.810 ;
        RECT 1848.830 910.675 1849.110 911.045 ;
        RECT 1849.750 910.675 1850.030 911.045 ;
        RECT 1849.760 910.530 1850.020 910.675 ;
        RECT 1852.060 910.530 1852.320 910.850 ;
        RECT 1852.120 862.765 1852.260 910.530 ;
        RECT 1851.130 862.395 1851.410 862.765 ;
        RECT 1852.050 862.395 1852.330 862.765 ;
        RECT 1851.200 821.285 1851.340 862.395 ;
        RECT 1850.210 820.915 1850.490 821.285 ;
        RECT 1851.130 820.915 1851.410 821.285 ;
        RECT 1850.280 787.965 1850.420 820.915 ;
        RECT 1850.210 787.595 1850.490 787.965 ;
        RECT 1850.210 772.635 1850.490 773.005 ;
        RECT 1850.220 772.490 1850.480 772.635 ;
        RECT 1850.220 737.810 1850.480 738.130 ;
        RECT 1850.280 724.610 1850.420 737.810 ;
        RECT 1850.280 724.470 1850.880 724.610 ;
        RECT 1850.740 691.405 1850.880 724.470 ;
        RECT 1850.670 691.035 1850.950 691.405 ;
        RECT 1850.210 676.075 1850.490 676.445 ;
        RECT 1850.220 675.930 1850.480 676.075 ;
        RECT 1850.220 641.250 1850.480 641.570 ;
        RECT 1850.280 628.050 1850.420 641.250 ;
        RECT 1850.280 627.910 1850.880 628.050 ;
        RECT 1850.740 603.830 1850.880 627.910 ;
        RECT 1850.680 603.510 1850.940 603.830 ;
        RECT 1850.680 602.830 1850.940 603.150 ;
        RECT 1850.740 545.350 1850.880 602.830 ;
        RECT 1850.680 545.030 1850.940 545.350 ;
        RECT 1850.680 531.430 1850.940 531.750 ;
        RECT 1850.740 507.010 1850.880 531.430 ;
        RECT 1850.740 506.870 1851.340 507.010 ;
        RECT 1851.200 483.325 1851.340 506.870 ;
        RECT 1850.210 482.955 1850.490 483.325 ;
        RECT 1851.130 482.955 1851.410 483.325 ;
        RECT 1850.280 434.510 1850.420 482.955 ;
        RECT 1850.220 434.190 1850.480 434.510 ;
        RECT 1850.220 386.250 1850.480 386.570 ;
        RECT 1850.280 305.650 1850.420 386.250 ;
        RECT 1850.220 305.330 1850.480 305.650 ;
        RECT 1850.680 241.410 1850.940 241.730 ;
        RECT 1850.740 207.390 1850.880 241.410 ;
        RECT 1850.680 207.070 1850.940 207.390 ;
        RECT 1849.760 192.790 1850.020 193.110 ;
        RECT 1849.820 169.310 1849.960 192.790 ;
        RECT 1849.760 168.990 1850.020 169.310 ;
        RECT 1851.140 168.990 1851.400 169.310 ;
        RECT 1851.200 96.890 1851.340 168.990 ;
        RECT 1850.220 96.570 1850.480 96.890 ;
        RECT 1851.140 96.570 1851.400 96.890 ;
        RECT 1850.280 48.010 1850.420 96.570 ;
        RECT 1850.280 47.870 1850.880 48.010 ;
        RECT 1850.740 41.470 1850.880 47.870 ;
        RECT 1370.440 41.150 1370.700 41.470 ;
        RECT 1850.680 41.150 1850.940 41.470 ;
        RECT 1370.500 2.400 1370.640 41.150 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
      LAYER via2 ;
        RECT 1849.750 1393.520 1850.030 1393.800 ;
        RECT 1851.590 1393.520 1851.870 1393.800 ;
        RECT 1850.210 1007.280 1850.490 1007.560 ;
        RECT 1851.130 1007.280 1851.410 1007.560 ;
        RECT 1848.830 910.720 1849.110 911.000 ;
        RECT 1849.750 910.720 1850.030 911.000 ;
        RECT 1851.130 862.440 1851.410 862.720 ;
        RECT 1852.050 862.440 1852.330 862.720 ;
        RECT 1850.210 820.960 1850.490 821.240 ;
        RECT 1851.130 820.960 1851.410 821.240 ;
        RECT 1850.210 787.640 1850.490 787.920 ;
        RECT 1850.210 772.680 1850.490 772.960 ;
        RECT 1850.670 691.080 1850.950 691.360 ;
        RECT 1850.210 676.120 1850.490 676.400 ;
        RECT 1850.210 483.000 1850.490 483.280 ;
        RECT 1851.130 483.000 1851.410 483.280 ;
      LAYER met3 ;
        RECT 1849.725 1393.810 1850.055 1393.825 ;
        RECT 1851.565 1393.810 1851.895 1393.825 ;
        RECT 1849.725 1393.510 1851.895 1393.810 ;
        RECT 1849.725 1393.495 1850.055 1393.510 ;
        RECT 1851.565 1393.495 1851.895 1393.510 ;
        RECT 1850.185 1007.570 1850.515 1007.585 ;
        RECT 1851.105 1007.570 1851.435 1007.585 ;
        RECT 1850.185 1007.270 1851.435 1007.570 ;
        RECT 1850.185 1007.255 1850.515 1007.270 ;
        RECT 1851.105 1007.255 1851.435 1007.270 ;
        RECT 1848.805 911.010 1849.135 911.025 ;
        RECT 1849.725 911.010 1850.055 911.025 ;
        RECT 1848.805 910.710 1850.055 911.010 ;
        RECT 1848.805 910.695 1849.135 910.710 ;
        RECT 1849.725 910.695 1850.055 910.710 ;
        RECT 1851.105 862.730 1851.435 862.745 ;
        RECT 1852.025 862.730 1852.355 862.745 ;
        RECT 1851.105 862.430 1852.355 862.730 ;
        RECT 1851.105 862.415 1851.435 862.430 ;
        RECT 1852.025 862.415 1852.355 862.430 ;
        RECT 1850.185 821.250 1850.515 821.265 ;
        RECT 1851.105 821.250 1851.435 821.265 ;
        RECT 1850.185 820.950 1851.435 821.250 ;
        RECT 1850.185 820.935 1850.515 820.950 ;
        RECT 1851.105 820.935 1851.435 820.950 ;
        RECT 1850.185 787.940 1850.515 787.945 ;
        RECT 1850.185 787.930 1850.770 787.940 ;
        RECT 1850.185 787.630 1850.970 787.930 ;
        RECT 1850.185 787.620 1850.770 787.630 ;
        RECT 1850.185 787.615 1850.515 787.620 ;
        RECT 1850.185 772.980 1850.515 772.985 ;
        RECT 1850.185 772.970 1850.770 772.980 ;
        RECT 1849.960 772.670 1850.770 772.970 ;
        RECT 1850.185 772.660 1850.770 772.670 ;
        RECT 1850.185 772.655 1850.515 772.660 ;
        RECT 1850.645 691.380 1850.975 691.385 ;
        RECT 1850.390 691.370 1850.975 691.380 ;
        RECT 1850.190 691.070 1850.975 691.370 ;
        RECT 1850.390 691.060 1850.975 691.070 ;
        RECT 1850.645 691.055 1850.975 691.060 ;
        RECT 1850.185 676.420 1850.515 676.425 ;
        RECT 1850.185 676.410 1850.770 676.420 ;
        RECT 1849.960 676.110 1850.770 676.410 ;
        RECT 1850.185 676.100 1850.770 676.110 ;
        RECT 1850.185 676.095 1850.515 676.100 ;
        RECT 1850.185 483.290 1850.515 483.305 ;
        RECT 1851.105 483.290 1851.435 483.305 ;
        RECT 1850.185 482.990 1851.435 483.290 ;
        RECT 1850.185 482.975 1850.515 482.990 ;
        RECT 1851.105 482.975 1851.435 482.990 ;
      LAYER via3 ;
        RECT 1850.420 787.620 1850.740 787.940 ;
        RECT 1850.420 772.660 1850.740 772.980 ;
        RECT 1850.420 691.060 1850.740 691.380 ;
        RECT 1850.420 676.100 1850.740 676.420 ;
      LAYER met4 ;
        RECT 1850.415 787.615 1850.745 787.945 ;
        RECT 1850.430 772.985 1850.730 787.615 ;
        RECT 1850.415 772.655 1850.745 772.985 ;
        RECT 1850.415 691.055 1850.745 691.385 ;
        RECT 1850.430 676.425 1850.730 691.055 ;
        RECT 1850.415 676.095 1850.745 676.425 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1388.350 37.640 1388.670 37.700 ;
        RECT 1863.530 37.640 1863.850 37.700 ;
        RECT 1388.350 37.500 1863.850 37.640 ;
        RECT 1388.350 37.440 1388.670 37.500 ;
        RECT 1863.530 37.440 1863.850 37.500 ;
      LAYER via ;
        RECT 1388.380 37.440 1388.640 37.700 ;
        RECT 1863.560 37.440 1863.820 37.700 ;
      LAYER met2 ;
        RECT 1863.020 1700.410 1863.300 1702.400 ;
        RECT 1863.020 1700.270 1863.760 1700.410 ;
        RECT 1863.020 1700.000 1863.300 1700.270 ;
        RECT 1863.620 37.730 1863.760 1700.270 ;
        RECT 1388.380 37.410 1388.640 37.730 ;
        RECT 1863.560 37.410 1863.820 37.730 ;
        RECT 1388.440 2.400 1388.580 37.410 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1406.290 37.300 1406.610 37.360 ;
        RECT 1870.430 37.300 1870.750 37.360 ;
        RECT 1406.290 37.160 1870.750 37.300 ;
        RECT 1406.290 37.100 1406.610 37.160 ;
        RECT 1870.430 37.100 1870.750 37.160 ;
      LAYER via ;
        RECT 1406.320 37.100 1406.580 37.360 ;
        RECT 1870.460 37.100 1870.720 37.360 ;
      LAYER met2 ;
        RECT 1872.220 1700.410 1872.500 1702.400 ;
        RECT 1870.520 1700.270 1872.500 1700.410 ;
        RECT 1870.520 37.390 1870.660 1700.270 ;
        RECT 1872.220 1700.000 1872.500 1700.270 ;
        RECT 1406.320 37.070 1406.580 37.390 ;
        RECT 1870.460 37.070 1870.720 37.390 ;
        RECT 1406.380 2.400 1406.520 37.070 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1877.865 1635.485 1878.035 1683.595 ;
        RECT 1878.785 1545.385 1878.955 1587.035 ;
        RECT 1877.405 1317.245 1877.575 1393.575 ;
        RECT 1877.865 1256.045 1878.035 1304.155 ;
        RECT 1877.865 241.485 1878.035 305.575 ;
        RECT 1877.405 186.405 1877.575 207.995 ;
      LAYER mcon ;
        RECT 1877.865 1683.425 1878.035 1683.595 ;
        RECT 1878.785 1586.865 1878.955 1587.035 ;
        RECT 1877.405 1393.405 1877.575 1393.575 ;
        RECT 1877.865 1303.985 1878.035 1304.155 ;
        RECT 1877.865 305.405 1878.035 305.575 ;
        RECT 1877.405 207.825 1877.575 207.995 ;
      LAYER met1 ;
        RECT 1877.805 1683.580 1878.095 1683.625 ;
        RECT 1878.710 1683.580 1879.030 1683.640 ;
        RECT 1877.805 1683.440 1879.030 1683.580 ;
        RECT 1877.805 1683.395 1878.095 1683.440 ;
        RECT 1878.710 1683.380 1879.030 1683.440 ;
        RECT 1877.790 1635.640 1878.110 1635.700 ;
        RECT 1877.595 1635.500 1878.110 1635.640 ;
        RECT 1877.790 1635.440 1878.110 1635.500 ;
        RECT 1877.790 1593.820 1878.110 1593.880 ;
        RECT 1878.710 1593.820 1879.030 1593.880 ;
        RECT 1877.790 1593.680 1879.030 1593.820 ;
        RECT 1877.790 1593.620 1878.110 1593.680 ;
        RECT 1878.710 1593.620 1879.030 1593.680 ;
        RECT 1878.710 1587.020 1879.030 1587.080 ;
        RECT 1878.515 1586.880 1879.030 1587.020 ;
        RECT 1878.710 1586.820 1879.030 1586.880 ;
        RECT 1878.710 1545.540 1879.030 1545.600 ;
        RECT 1878.515 1545.400 1879.030 1545.540 ;
        RECT 1878.710 1545.340 1879.030 1545.400 ;
        RECT 1878.250 1497.600 1878.570 1497.660 ;
        RECT 1878.710 1497.600 1879.030 1497.660 ;
        RECT 1878.250 1497.460 1879.030 1497.600 ;
        RECT 1878.250 1497.400 1878.570 1497.460 ;
        RECT 1878.710 1497.400 1879.030 1497.460 ;
        RECT 1877.790 1448.980 1878.110 1449.040 ;
        RECT 1878.710 1448.980 1879.030 1449.040 ;
        RECT 1877.790 1448.840 1879.030 1448.980 ;
        RECT 1877.790 1448.780 1878.110 1448.840 ;
        RECT 1878.710 1448.780 1879.030 1448.840 ;
        RECT 1877.330 1400.700 1877.650 1400.760 ;
        RECT 1878.710 1400.700 1879.030 1400.760 ;
        RECT 1877.330 1400.560 1879.030 1400.700 ;
        RECT 1877.330 1400.500 1877.650 1400.560 ;
        RECT 1878.710 1400.500 1879.030 1400.560 ;
        RECT 1877.330 1393.560 1877.650 1393.620 ;
        RECT 1877.135 1393.420 1877.650 1393.560 ;
        RECT 1877.330 1393.360 1877.650 1393.420 ;
        RECT 1877.345 1317.400 1877.635 1317.445 ;
        RECT 1878.250 1317.400 1878.570 1317.460 ;
        RECT 1877.345 1317.260 1878.570 1317.400 ;
        RECT 1877.345 1317.215 1877.635 1317.260 ;
        RECT 1878.250 1317.200 1878.570 1317.260 ;
        RECT 1877.805 1304.140 1878.095 1304.185 ;
        RECT 1878.250 1304.140 1878.570 1304.200 ;
        RECT 1877.805 1304.000 1878.570 1304.140 ;
        RECT 1877.805 1303.955 1878.095 1304.000 ;
        RECT 1878.250 1303.940 1878.570 1304.000 ;
        RECT 1877.790 1256.200 1878.110 1256.260 ;
        RECT 1877.595 1256.060 1878.110 1256.200 ;
        RECT 1877.790 1256.000 1878.110 1256.060 ;
        RECT 1878.710 1207.580 1879.030 1207.640 ;
        RECT 1879.170 1207.580 1879.490 1207.640 ;
        RECT 1878.710 1207.440 1879.490 1207.580 ;
        RECT 1878.710 1207.380 1879.030 1207.440 ;
        RECT 1879.170 1207.380 1879.490 1207.440 ;
        RECT 1877.790 1159.300 1878.110 1159.360 ;
        RECT 1879.170 1159.300 1879.490 1159.360 ;
        RECT 1877.790 1159.160 1879.490 1159.300 ;
        RECT 1877.790 1159.100 1878.110 1159.160 ;
        RECT 1879.170 1159.100 1879.490 1159.160 ;
        RECT 1877.790 1062.740 1878.110 1062.800 ;
        RECT 1879.170 1062.740 1879.490 1062.800 ;
        RECT 1877.790 1062.600 1879.490 1062.740 ;
        RECT 1877.790 1062.540 1878.110 1062.600 ;
        RECT 1879.170 1062.540 1879.490 1062.600 ;
        RECT 1877.790 1007.320 1878.110 1007.380 ;
        RECT 1879.170 1007.320 1879.490 1007.380 ;
        RECT 1877.790 1007.180 1879.490 1007.320 ;
        RECT 1877.790 1007.120 1878.110 1007.180 ;
        RECT 1879.170 1007.120 1879.490 1007.180 ;
        RECT 1877.330 959.040 1877.650 959.100 ;
        RECT 1877.790 959.040 1878.110 959.100 ;
        RECT 1877.330 958.900 1878.110 959.040 ;
        RECT 1877.330 958.840 1877.650 958.900 ;
        RECT 1877.790 958.840 1878.110 958.900 ;
        RECT 1875.950 821.000 1876.270 821.060 ;
        RECT 1877.790 821.000 1878.110 821.060 ;
        RECT 1875.950 820.860 1878.110 821.000 ;
        RECT 1875.950 820.800 1876.270 820.860 ;
        RECT 1877.790 820.800 1878.110 820.860 ;
        RECT 1877.790 772.720 1878.110 772.780 ;
        RECT 1878.710 772.720 1879.030 772.780 ;
        RECT 1877.790 772.580 1879.030 772.720 ;
        RECT 1877.790 772.520 1878.110 772.580 ;
        RECT 1878.710 772.520 1879.030 772.580 ;
        RECT 1877.790 675.960 1878.110 676.220 ;
        RECT 1877.880 675.820 1878.020 675.960 ;
        RECT 1878.710 675.820 1879.030 675.880 ;
        RECT 1877.880 675.680 1879.030 675.820 ;
        RECT 1878.710 675.620 1879.030 675.680 ;
        RECT 1877.330 603.740 1877.650 603.800 ;
        RECT 1878.710 603.740 1879.030 603.800 ;
        RECT 1877.330 603.600 1879.030 603.740 ;
        RECT 1877.330 603.540 1877.650 603.600 ;
        RECT 1878.710 603.540 1879.030 603.600 ;
        RECT 1877.330 579.600 1877.650 579.660 ;
        RECT 1878.710 579.600 1879.030 579.660 ;
        RECT 1877.330 579.460 1879.030 579.600 ;
        RECT 1877.330 579.400 1877.650 579.460 ;
        RECT 1878.710 579.400 1879.030 579.460 ;
        RECT 1877.790 305.560 1878.110 305.620 ;
        RECT 1877.595 305.420 1878.110 305.560 ;
        RECT 1877.790 305.360 1878.110 305.420 ;
        RECT 1877.805 241.640 1878.095 241.685 ;
        RECT 1878.250 241.640 1878.570 241.700 ;
        RECT 1877.805 241.500 1878.570 241.640 ;
        RECT 1877.805 241.455 1878.095 241.500 ;
        RECT 1878.250 241.440 1878.570 241.500 ;
        RECT 1877.345 207.980 1877.635 208.025 ;
        RECT 1878.250 207.980 1878.570 208.040 ;
        RECT 1877.345 207.840 1878.570 207.980 ;
        RECT 1877.345 207.795 1877.635 207.840 ;
        RECT 1878.250 207.780 1878.570 207.840 ;
        RECT 1877.330 186.560 1877.650 186.620 ;
        RECT 1877.135 186.420 1877.650 186.560 ;
        RECT 1877.330 186.360 1877.650 186.420 ;
        RECT 1877.790 96.800 1878.110 96.860 ;
        RECT 1878.710 96.800 1879.030 96.860 ;
        RECT 1877.790 96.660 1879.030 96.800 ;
        RECT 1877.790 96.600 1878.110 96.660 ;
        RECT 1878.710 96.600 1879.030 96.660 ;
        RECT 1423.770 36.960 1424.090 37.020 ;
        RECT 1877.790 36.960 1878.110 37.020 ;
        RECT 1423.770 36.820 1878.110 36.960 ;
        RECT 1423.770 36.760 1424.090 36.820 ;
        RECT 1877.790 36.760 1878.110 36.820 ;
      LAYER via ;
        RECT 1878.740 1683.380 1879.000 1683.640 ;
        RECT 1877.820 1635.440 1878.080 1635.700 ;
        RECT 1877.820 1593.620 1878.080 1593.880 ;
        RECT 1878.740 1593.620 1879.000 1593.880 ;
        RECT 1878.740 1586.820 1879.000 1587.080 ;
        RECT 1878.740 1545.340 1879.000 1545.600 ;
        RECT 1878.280 1497.400 1878.540 1497.660 ;
        RECT 1878.740 1497.400 1879.000 1497.660 ;
        RECT 1877.820 1448.780 1878.080 1449.040 ;
        RECT 1878.740 1448.780 1879.000 1449.040 ;
        RECT 1877.360 1400.500 1877.620 1400.760 ;
        RECT 1878.740 1400.500 1879.000 1400.760 ;
        RECT 1877.360 1393.360 1877.620 1393.620 ;
        RECT 1878.280 1317.200 1878.540 1317.460 ;
        RECT 1878.280 1303.940 1878.540 1304.200 ;
        RECT 1877.820 1256.000 1878.080 1256.260 ;
        RECT 1878.740 1207.380 1879.000 1207.640 ;
        RECT 1879.200 1207.380 1879.460 1207.640 ;
        RECT 1877.820 1159.100 1878.080 1159.360 ;
        RECT 1879.200 1159.100 1879.460 1159.360 ;
        RECT 1877.820 1062.540 1878.080 1062.800 ;
        RECT 1879.200 1062.540 1879.460 1062.800 ;
        RECT 1877.820 1007.120 1878.080 1007.380 ;
        RECT 1879.200 1007.120 1879.460 1007.380 ;
        RECT 1877.360 958.840 1877.620 959.100 ;
        RECT 1877.820 958.840 1878.080 959.100 ;
        RECT 1875.980 820.800 1876.240 821.060 ;
        RECT 1877.820 820.800 1878.080 821.060 ;
        RECT 1877.820 772.520 1878.080 772.780 ;
        RECT 1878.740 772.520 1879.000 772.780 ;
        RECT 1877.820 675.960 1878.080 676.220 ;
        RECT 1878.740 675.620 1879.000 675.880 ;
        RECT 1877.360 603.540 1877.620 603.800 ;
        RECT 1878.740 603.540 1879.000 603.800 ;
        RECT 1877.360 579.400 1877.620 579.660 ;
        RECT 1878.740 579.400 1879.000 579.660 ;
        RECT 1877.820 305.360 1878.080 305.620 ;
        RECT 1878.280 241.440 1878.540 241.700 ;
        RECT 1878.280 207.780 1878.540 208.040 ;
        RECT 1877.360 186.360 1877.620 186.620 ;
        RECT 1877.820 96.600 1878.080 96.860 ;
        RECT 1878.740 96.600 1879.000 96.860 ;
        RECT 1423.800 36.760 1424.060 37.020 ;
        RECT 1877.820 36.760 1878.080 37.020 ;
      LAYER met2 ;
        RECT 1881.420 1701.090 1881.700 1702.400 ;
        RECT 1878.800 1700.950 1881.700 1701.090 ;
        RECT 1878.800 1683.670 1878.940 1700.950 ;
        RECT 1881.420 1700.000 1881.700 1700.950 ;
        RECT 1878.740 1683.350 1879.000 1683.670 ;
        RECT 1877.820 1635.410 1878.080 1635.730 ;
        RECT 1877.880 1593.910 1878.020 1635.410 ;
        RECT 1877.820 1593.590 1878.080 1593.910 ;
        RECT 1878.740 1593.590 1879.000 1593.910 ;
        RECT 1878.800 1587.110 1878.940 1593.590 ;
        RECT 1878.740 1586.790 1879.000 1587.110 ;
        RECT 1878.740 1545.310 1879.000 1545.630 ;
        RECT 1878.800 1497.690 1878.940 1545.310 ;
        RECT 1878.280 1497.370 1878.540 1497.690 ;
        RECT 1878.740 1497.370 1879.000 1497.690 ;
        RECT 1878.340 1463.090 1878.480 1497.370 ;
        RECT 1877.880 1462.950 1878.480 1463.090 ;
        RECT 1877.880 1449.070 1878.020 1462.950 ;
        RECT 1877.820 1448.750 1878.080 1449.070 ;
        RECT 1878.740 1448.750 1879.000 1449.070 ;
        RECT 1878.800 1400.790 1878.940 1448.750 ;
        RECT 1877.360 1400.470 1877.620 1400.790 ;
        RECT 1878.740 1400.470 1879.000 1400.790 ;
        RECT 1877.420 1393.650 1877.560 1400.470 ;
        RECT 1877.360 1393.330 1877.620 1393.650 ;
        RECT 1878.280 1317.170 1878.540 1317.490 ;
        RECT 1878.340 1304.230 1878.480 1317.170 ;
        RECT 1878.280 1303.910 1878.540 1304.230 ;
        RECT 1877.820 1255.970 1878.080 1256.290 ;
        RECT 1877.880 1255.805 1878.020 1255.970 ;
        RECT 1877.810 1255.435 1878.090 1255.805 ;
        RECT 1878.730 1255.435 1879.010 1255.805 ;
        RECT 1878.800 1207.670 1878.940 1255.435 ;
        RECT 1878.740 1207.350 1879.000 1207.670 ;
        RECT 1879.200 1207.350 1879.460 1207.670 ;
        RECT 1879.260 1159.390 1879.400 1207.350 ;
        RECT 1877.820 1159.245 1878.080 1159.390 ;
        RECT 1879.200 1159.245 1879.460 1159.390 ;
        RECT 1877.810 1158.875 1878.090 1159.245 ;
        RECT 1879.190 1158.875 1879.470 1159.245 ;
        RECT 1879.260 1062.830 1879.400 1158.875 ;
        RECT 1877.820 1062.685 1878.080 1062.830 ;
        RECT 1879.200 1062.685 1879.460 1062.830 ;
        RECT 1877.810 1062.315 1878.090 1062.685 ;
        RECT 1879.190 1062.315 1879.470 1062.685 ;
        RECT 1879.260 1007.410 1879.400 1062.315 ;
        RECT 1877.820 1007.090 1878.080 1007.410 ;
        RECT 1879.200 1007.090 1879.460 1007.410 ;
        RECT 1877.880 960.005 1878.020 1007.090 ;
        RECT 1877.810 959.635 1878.090 960.005 ;
        RECT 1877.360 958.810 1877.620 959.130 ;
        RECT 1877.810 958.955 1878.090 959.325 ;
        RECT 1877.820 958.810 1878.080 958.955 ;
        RECT 1877.420 911.045 1877.560 958.810 ;
        RECT 1877.350 910.675 1877.630 911.045 ;
        RECT 1878.730 910.675 1879.010 911.045 ;
        RECT 1878.800 862.765 1878.940 910.675 ;
        RECT 1877.810 862.395 1878.090 862.765 ;
        RECT 1878.730 862.395 1879.010 862.765 ;
        RECT 1877.880 821.090 1878.020 862.395 ;
        RECT 1875.980 820.770 1876.240 821.090 ;
        RECT 1877.820 820.770 1878.080 821.090 ;
        RECT 1876.040 773.005 1876.180 820.770 ;
        RECT 1875.970 772.635 1876.250 773.005 ;
        RECT 1877.810 772.635 1878.090 773.005 ;
        RECT 1877.820 772.490 1878.080 772.635 ;
        RECT 1878.740 772.490 1879.000 772.810 ;
        RECT 1878.800 677.125 1878.940 772.490 ;
        RECT 1878.730 676.755 1879.010 677.125 ;
        RECT 1877.810 676.075 1878.090 676.445 ;
        RECT 1877.820 675.930 1878.080 676.075 ;
        RECT 1878.740 675.590 1879.000 675.910 ;
        RECT 1878.800 603.830 1878.940 675.590 ;
        RECT 1877.360 603.510 1877.620 603.830 ;
        RECT 1878.740 603.510 1879.000 603.830 ;
        RECT 1877.420 579.690 1877.560 603.510 ;
        RECT 1877.360 579.370 1877.620 579.690 ;
        RECT 1878.740 579.370 1879.000 579.690 ;
        RECT 1878.800 484.005 1878.940 579.370 ;
        RECT 1878.730 483.635 1879.010 484.005 ;
        RECT 1877.810 482.955 1878.090 483.325 ;
        RECT 1877.880 305.650 1878.020 482.955 ;
        RECT 1877.820 305.330 1878.080 305.650 ;
        RECT 1878.280 241.410 1878.540 241.730 ;
        RECT 1878.340 208.070 1878.480 241.410 ;
        RECT 1878.280 207.750 1878.540 208.070 ;
        RECT 1877.360 186.330 1877.620 186.650 ;
        RECT 1877.420 169.050 1877.560 186.330 ;
        RECT 1877.420 168.910 1878.940 169.050 ;
        RECT 1878.800 96.890 1878.940 168.910 ;
        RECT 1877.820 96.570 1878.080 96.890 ;
        RECT 1878.740 96.570 1879.000 96.890 ;
        RECT 1877.880 37.050 1878.020 96.570 ;
        RECT 1423.800 36.730 1424.060 37.050 ;
        RECT 1877.820 36.730 1878.080 37.050 ;
        RECT 1423.860 2.400 1424.000 36.730 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
      LAYER via2 ;
        RECT 1877.810 1255.480 1878.090 1255.760 ;
        RECT 1878.730 1255.480 1879.010 1255.760 ;
        RECT 1877.810 1158.920 1878.090 1159.200 ;
        RECT 1879.190 1158.920 1879.470 1159.200 ;
        RECT 1877.810 1062.360 1878.090 1062.640 ;
        RECT 1879.190 1062.360 1879.470 1062.640 ;
        RECT 1877.810 959.680 1878.090 959.960 ;
        RECT 1877.810 959.000 1878.090 959.280 ;
        RECT 1877.350 910.720 1877.630 911.000 ;
        RECT 1878.730 910.720 1879.010 911.000 ;
        RECT 1877.810 862.440 1878.090 862.720 ;
        RECT 1878.730 862.440 1879.010 862.720 ;
        RECT 1875.970 772.680 1876.250 772.960 ;
        RECT 1877.810 772.680 1878.090 772.960 ;
        RECT 1878.730 676.800 1879.010 677.080 ;
        RECT 1877.810 676.120 1878.090 676.400 ;
        RECT 1878.730 483.680 1879.010 483.960 ;
        RECT 1877.810 483.000 1878.090 483.280 ;
      LAYER met3 ;
        RECT 1877.785 1255.770 1878.115 1255.785 ;
        RECT 1878.705 1255.770 1879.035 1255.785 ;
        RECT 1877.785 1255.470 1879.035 1255.770 ;
        RECT 1877.785 1255.455 1878.115 1255.470 ;
        RECT 1878.705 1255.455 1879.035 1255.470 ;
        RECT 1877.785 1159.210 1878.115 1159.225 ;
        RECT 1879.165 1159.210 1879.495 1159.225 ;
        RECT 1877.785 1158.910 1879.495 1159.210 ;
        RECT 1877.785 1158.895 1878.115 1158.910 ;
        RECT 1879.165 1158.895 1879.495 1158.910 ;
        RECT 1877.785 1062.650 1878.115 1062.665 ;
        RECT 1879.165 1062.650 1879.495 1062.665 ;
        RECT 1877.785 1062.350 1879.495 1062.650 ;
        RECT 1877.785 1062.335 1878.115 1062.350 ;
        RECT 1879.165 1062.335 1879.495 1062.350 ;
        RECT 1877.785 959.970 1878.115 959.985 ;
        RECT 1877.110 959.670 1878.115 959.970 ;
        RECT 1877.110 959.290 1877.410 959.670 ;
        RECT 1877.785 959.655 1878.115 959.670 ;
        RECT 1877.785 959.290 1878.115 959.305 ;
        RECT 1877.110 958.990 1878.115 959.290 ;
        RECT 1877.785 958.975 1878.115 958.990 ;
        RECT 1877.325 911.010 1877.655 911.025 ;
        RECT 1878.705 911.010 1879.035 911.025 ;
        RECT 1877.325 910.710 1879.035 911.010 ;
        RECT 1877.325 910.695 1877.655 910.710 ;
        RECT 1878.705 910.695 1879.035 910.710 ;
        RECT 1877.785 862.730 1878.115 862.745 ;
        RECT 1878.705 862.730 1879.035 862.745 ;
        RECT 1877.785 862.430 1879.035 862.730 ;
        RECT 1877.785 862.415 1878.115 862.430 ;
        RECT 1878.705 862.415 1879.035 862.430 ;
        RECT 1875.945 772.970 1876.275 772.985 ;
        RECT 1877.785 772.970 1878.115 772.985 ;
        RECT 1875.945 772.670 1878.115 772.970 ;
        RECT 1875.945 772.655 1876.275 772.670 ;
        RECT 1877.785 772.655 1878.115 772.670 ;
        RECT 1878.705 677.090 1879.035 677.105 ;
        RECT 1877.110 676.790 1879.035 677.090 ;
        RECT 1877.110 676.410 1877.410 676.790 ;
        RECT 1878.705 676.775 1879.035 676.790 ;
        RECT 1877.785 676.410 1878.115 676.425 ;
        RECT 1877.110 676.110 1878.115 676.410 ;
        RECT 1877.785 676.095 1878.115 676.110 ;
        RECT 1878.705 483.970 1879.035 483.985 ;
        RECT 1877.110 483.670 1879.035 483.970 ;
        RECT 1877.110 483.290 1877.410 483.670 ;
        RECT 1878.705 483.655 1879.035 483.670 ;
        RECT 1877.785 483.290 1878.115 483.305 ;
        RECT 1877.110 482.990 1878.115 483.290 ;
        RECT 1877.785 482.975 1878.115 482.990 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1464.710 51.580 1465.030 51.640 ;
        RECT 1891.590 51.580 1891.910 51.640 ;
        RECT 1464.710 51.440 1891.910 51.580 ;
        RECT 1464.710 51.380 1465.030 51.440 ;
        RECT 1891.590 51.380 1891.910 51.440 ;
        RECT 1441.710 16.220 1442.030 16.280 ;
        RECT 1464.710 16.220 1465.030 16.280 ;
        RECT 1441.710 16.080 1465.030 16.220 ;
        RECT 1441.710 16.020 1442.030 16.080 ;
        RECT 1464.710 16.020 1465.030 16.080 ;
      LAYER via ;
        RECT 1464.740 51.380 1465.000 51.640 ;
        RECT 1891.620 51.380 1891.880 51.640 ;
        RECT 1441.740 16.020 1442.000 16.280 ;
        RECT 1464.740 16.020 1465.000 16.280 ;
      LAYER met2 ;
        RECT 1890.620 1700.410 1890.900 1702.400 ;
        RECT 1890.620 1700.270 1891.820 1700.410 ;
        RECT 1890.620 1700.000 1890.900 1700.270 ;
        RECT 1891.680 51.670 1891.820 1700.270 ;
        RECT 1464.740 51.350 1465.000 51.670 ;
        RECT 1891.620 51.350 1891.880 51.670 ;
        RECT 1464.800 16.310 1464.940 51.350 ;
        RECT 1441.740 15.990 1442.000 16.310 ;
        RECT 1464.740 15.990 1465.000 16.310 ;
        RECT 1441.800 2.400 1441.940 15.990 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1498.290 52.260 1498.610 52.320 ;
        RECT 1898.030 52.260 1898.350 52.320 ;
        RECT 1498.290 52.120 1898.350 52.260 ;
        RECT 1498.290 52.060 1498.610 52.120 ;
        RECT 1898.030 52.060 1898.350 52.120 ;
        RECT 1459.650 18.260 1459.970 18.320 ;
        RECT 1498.290 18.260 1498.610 18.320 ;
        RECT 1459.650 18.120 1498.610 18.260 ;
        RECT 1459.650 18.060 1459.970 18.120 ;
        RECT 1498.290 18.060 1498.610 18.120 ;
      LAYER via ;
        RECT 1498.320 52.060 1498.580 52.320 ;
        RECT 1898.060 52.060 1898.320 52.320 ;
        RECT 1459.680 18.060 1459.940 18.320 ;
        RECT 1498.320 18.060 1498.580 18.320 ;
      LAYER met2 ;
        RECT 1899.820 1700.410 1900.100 1702.400 ;
        RECT 1898.120 1700.270 1900.100 1700.410 ;
        RECT 1898.120 52.350 1898.260 1700.270 ;
        RECT 1899.820 1700.000 1900.100 1700.270 ;
        RECT 1498.320 52.030 1498.580 52.350 ;
        RECT 1898.060 52.030 1898.320 52.350 ;
        RECT 1498.380 18.350 1498.520 52.030 ;
        RECT 1459.680 18.030 1459.940 18.350 ;
        RECT 1498.320 18.030 1498.580 18.350 ;
        RECT 1459.740 2.400 1459.880 18.030 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1906.385 1538.925 1906.555 1587.035 ;
        RECT 1905.465 1304.325 1905.635 1352.095 ;
        RECT 1905.465 1207.425 1905.635 1255.535 ;
        RECT 1905.465 1159.145 1905.635 1173.595 ;
        RECT 1905.925 1110.865 1906.095 1124.975 ;
        RECT 1905.465 1062.585 1905.635 1077.035 ;
        RECT 1905.005 737.885 1905.175 814.215 ;
        RECT 1905.005 41.565 1905.175 89.675 ;
      LAYER mcon ;
        RECT 1906.385 1586.865 1906.555 1587.035 ;
        RECT 1905.465 1351.925 1905.635 1352.095 ;
        RECT 1905.465 1255.365 1905.635 1255.535 ;
        RECT 1905.465 1173.425 1905.635 1173.595 ;
        RECT 1905.925 1124.805 1906.095 1124.975 ;
        RECT 1905.465 1076.865 1905.635 1077.035 ;
        RECT 1905.005 814.045 1905.175 814.215 ;
        RECT 1905.005 89.505 1905.175 89.675 ;
      LAYER met1 ;
        RECT 1904.930 1683.580 1905.250 1683.640 ;
        RECT 1906.770 1683.580 1907.090 1683.640 ;
        RECT 1904.930 1683.440 1907.090 1683.580 ;
        RECT 1904.930 1683.380 1905.250 1683.440 ;
        RECT 1906.770 1683.380 1907.090 1683.440 ;
        RECT 1905.390 1593.820 1905.710 1593.880 ;
        RECT 1906.310 1593.820 1906.630 1593.880 ;
        RECT 1905.390 1593.680 1906.630 1593.820 ;
        RECT 1905.390 1593.620 1905.710 1593.680 ;
        RECT 1906.310 1593.620 1906.630 1593.680 ;
        RECT 1906.310 1587.020 1906.630 1587.080 ;
        RECT 1906.115 1586.880 1906.630 1587.020 ;
        RECT 1906.310 1586.820 1906.630 1586.880 ;
        RECT 1906.310 1539.080 1906.630 1539.140 ;
        RECT 1906.115 1538.940 1906.630 1539.080 ;
        RECT 1906.310 1538.880 1906.630 1538.940 ;
        RECT 1905.390 1449.320 1905.710 1449.380 ;
        RECT 1906.770 1449.320 1907.090 1449.380 ;
        RECT 1905.390 1449.180 1907.090 1449.320 ;
        RECT 1905.390 1449.120 1905.710 1449.180 ;
        RECT 1906.770 1449.120 1907.090 1449.180 ;
        RECT 1905.390 1414.440 1905.710 1414.700 ;
        RECT 1905.480 1413.960 1905.620 1414.440 ;
        RECT 1905.850 1413.960 1906.170 1414.020 ;
        RECT 1905.480 1413.820 1906.170 1413.960 ;
        RECT 1905.850 1413.760 1906.170 1413.820 ;
        RECT 1904.930 1352.760 1905.250 1352.820 ;
        RECT 1905.390 1352.760 1905.710 1352.820 ;
        RECT 1904.930 1352.620 1905.710 1352.760 ;
        RECT 1904.930 1352.560 1905.250 1352.620 ;
        RECT 1905.390 1352.560 1905.710 1352.620 ;
        RECT 1905.390 1352.080 1905.710 1352.140 ;
        RECT 1905.195 1351.940 1905.710 1352.080 ;
        RECT 1905.390 1351.880 1905.710 1351.940 ;
        RECT 1905.405 1304.480 1905.695 1304.525 ;
        RECT 1905.850 1304.480 1906.170 1304.540 ;
        RECT 1905.405 1304.340 1906.170 1304.480 ;
        RECT 1905.405 1304.295 1905.695 1304.340 ;
        RECT 1905.850 1304.280 1906.170 1304.340 ;
        RECT 1905.390 1256.200 1905.710 1256.260 ;
        RECT 1906.770 1256.200 1907.090 1256.260 ;
        RECT 1905.390 1256.060 1907.090 1256.200 ;
        RECT 1905.390 1256.000 1905.710 1256.060 ;
        RECT 1906.770 1256.000 1907.090 1256.060 ;
        RECT 1905.390 1255.520 1905.710 1255.580 ;
        RECT 1905.195 1255.380 1905.710 1255.520 ;
        RECT 1905.390 1255.320 1905.710 1255.380 ;
        RECT 1905.405 1207.580 1905.695 1207.625 ;
        RECT 1905.850 1207.580 1906.170 1207.640 ;
        RECT 1905.405 1207.440 1906.170 1207.580 ;
        RECT 1905.405 1207.395 1905.695 1207.440 ;
        RECT 1905.850 1207.380 1906.170 1207.440 ;
        RECT 1905.390 1173.580 1905.710 1173.640 ;
        RECT 1905.195 1173.440 1905.710 1173.580 ;
        RECT 1905.390 1173.380 1905.710 1173.440 ;
        RECT 1905.405 1159.300 1905.695 1159.345 ;
        RECT 1905.850 1159.300 1906.170 1159.360 ;
        RECT 1905.405 1159.160 1906.170 1159.300 ;
        RECT 1905.405 1159.115 1905.695 1159.160 ;
        RECT 1905.850 1159.100 1906.170 1159.160 ;
        RECT 1905.850 1124.960 1906.170 1125.020 ;
        RECT 1905.655 1124.820 1906.170 1124.960 ;
        RECT 1905.850 1124.760 1906.170 1124.820 ;
        RECT 1905.850 1111.020 1906.170 1111.080 ;
        RECT 1905.655 1110.880 1906.170 1111.020 ;
        RECT 1905.850 1110.820 1906.170 1110.880 ;
        RECT 1905.390 1077.020 1905.710 1077.080 ;
        RECT 1905.195 1076.880 1905.710 1077.020 ;
        RECT 1905.390 1076.820 1905.710 1076.880 ;
        RECT 1905.405 1062.740 1905.695 1062.785 ;
        RECT 1905.850 1062.740 1906.170 1062.800 ;
        RECT 1905.405 1062.600 1906.170 1062.740 ;
        RECT 1905.405 1062.555 1905.695 1062.600 ;
        RECT 1905.850 1062.540 1906.170 1062.600 ;
        RECT 1905.850 1028.200 1906.170 1028.460 ;
        RECT 1905.940 1027.780 1906.080 1028.200 ;
        RECT 1905.850 1027.520 1906.170 1027.780 ;
        RECT 1905.390 1007.320 1905.710 1007.380 ;
        RECT 1906.770 1007.320 1907.090 1007.380 ;
        RECT 1905.390 1007.180 1907.090 1007.320 ;
        RECT 1905.390 1007.120 1905.710 1007.180 ;
        RECT 1906.770 1007.120 1907.090 1007.180 ;
        RECT 1905.850 917.900 1906.170 917.960 ;
        RECT 1906.770 917.900 1907.090 917.960 ;
        RECT 1905.850 917.760 1907.090 917.900 ;
        RECT 1905.850 917.700 1906.170 917.760 ;
        RECT 1906.770 917.700 1907.090 917.760 ;
        RECT 1904.010 869.620 1904.330 869.680 ;
        RECT 1904.930 869.620 1905.250 869.680 ;
        RECT 1904.010 869.480 1905.250 869.620 ;
        RECT 1904.010 869.420 1904.330 869.480 ;
        RECT 1904.930 869.420 1905.250 869.480 ;
        RECT 1904.930 820.660 1905.250 820.720 ;
        RECT 1905.390 820.660 1905.710 820.720 ;
        RECT 1904.930 820.520 1905.710 820.660 ;
        RECT 1904.930 820.460 1905.250 820.520 ;
        RECT 1905.390 820.460 1905.710 820.520 ;
        RECT 1904.930 814.200 1905.250 814.260 ;
        RECT 1904.735 814.060 1905.250 814.200 ;
        RECT 1904.930 814.000 1905.250 814.060 ;
        RECT 1904.945 738.040 1905.235 738.085 ;
        RECT 1905.390 738.040 1905.710 738.100 ;
        RECT 1904.945 737.900 1905.710 738.040 ;
        RECT 1904.945 737.855 1905.235 737.900 ;
        RECT 1905.390 737.840 1905.710 737.900 ;
        RECT 1905.390 676.500 1905.710 676.560 ;
        RECT 1906.310 676.500 1906.630 676.560 ;
        RECT 1905.390 676.360 1906.630 676.500 ;
        RECT 1905.390 676.300 1905.710 676.360 ;
        RECT 1906.310 676.300 1906.630 676.360 ;
        RECT 1905.390 641.620 1905.710 641.880 ;
        RECT 1905.480 641.480 1905.620 641.620 ;
        RECT 1905.850 641.480 1906.170 641.540 ;
        RECT 1905.480 641.340 1906.170 641.480 ;
        RECT 1905.850 641.280 1906.170 641.340 ;
        RECT 1905.390 579.600 1905.710 579.660 ;
        RECT 1906.310 579.600 1906.630 579.660 ;
        RECT 1905.390 579.460 1906.630 579.600 ;
        RECT 1905.390 579.400 1905.710 579.460 ;
        RECT 1906.310 579.400 1906.630 579.460 ;
        RECT 1905.390 386.480 1905.710 386.540 ;
        RECT 1905.850 386.480 1906.170 386.540 ;
        RECT 1905.390 386.340 1906.170 386.480 ;
        RECT 1905.390 386.280 1905.710 386.340 ;
        RECT 1905.850 386.280 1906.170 386.340 ;
        RECT 1905.850 241.300 1906.170 241.360 ;
        RECT 1906.310 241.300 1906.630 241.360 ;
        RECT 1905.850 241.160 1906.630 241.300 ;
        RECT 1905.850 241.100 1906.170 241.160 ;
        RECT 1906.310 241.100 1906.630 241.160 ;
        RECT 1905.850 145.080 1906.170 145.140 ;
        RECT 1906.310 145.080 1906.630 145.140 ;
        RECT 1905.850 144.940 1906.630 145.080 ;
        RECT 1905.850 144.880 1906.170 144.940 ;
        RECT 1906.310 144.880 1906.630 144.940 ;
        RECT 1905.390 96.800 1905.710 96.860 ;
        RECT 1906.310 96.800 1906.630 96.860 ;
        RECT 1905.390 96.660 1906.630 96.800 ;
        RECT 1905.390 96.600 1905.710 96.660 ;
        RECT 1906.310 96.600 1906.630 96.660 ;
        RECT 1904.945 89.660 1905.235 89.705 ;
        RECT 1905.390 89.660 1905.710 89.720 ;
        RECT 1904.945 89.520 1905.710 89.660 ;
        RECT 1904.945 89.475 1905.235 89.520 ;
        RECT 1905.390 89.460 1905.710 89.520 ;
        RECT 1904.930 41.720 1905.250 41.780 ;
        RECT 1904.735 41.580 1905.250 41.720 ;
        RECT 1904.930 41.520 1905.250 41.580 ;
        RECT 1593.970 33.560 1594.290 33.620 ;
        RECT 1904.930 33.560 1905.250 33.620 ;
        RECT 1593.970 33.420 1905.250 33.560 ;
        RECT 1593.970 33.360 1594.290 33.420 ;
        RECT 1904.930 33.360 1905.250 33.420 ;
        RECT 1477.590 16.900 1477.910 16.960 ;
        RECT 1593.970 16.900 1594.290 16.960 ;
        RECT 1477.590 16.760 1594.290 16.900 ;
        RECT 1477.590 16.700 1477.910 16.760 ;
        RECT 1593.970 16.700 1594.290 16.760 ;
      LAYER via ;
        RECT 1904.960 1683.380 1905.220 1683.640 ;
        RECT 1906.800 1683.380 1907.060 1683.640 ;
        RECT 1905.420 1593.620 1905.680 1593.880 ;
        RECT 1906.340 1593.620 1906.600 1593.880 ;
        RECT 1906.340 1586.820 1906.600 1587.080 ;
        RECT 1906.340 1538.880 1906.600 1539.140 ;
        RECT 1905.420 1449.120 1905.680 1449.380 ;
        RECT 1906.800 1449.120 1907.060 1449.380 ;
        RECT 1905.420 1414.440 1905.680 1414.700 ;
        RECT 1905.880 1413.760 1906.140 1414.020 ;
        RECT 1904.960 1352.560 1905.220 1352.820 ;
        RECT 1905.420 1352.560 1905.680 1352.820 ;
        RECT 1905.420 1351.880 1905.680 1352.140 ;
        RECT 1905.880 1304.280 1906.140 1304.540 ;
        RECT 1905.420 1256.000 1905.680 1256.260 ;
        RECT 1906.800 1256.000 1907.060 1256.260 ;
        RECT 1905.420 1255.320 1905.680 1255.580 ;
        RECT 1905.880 1207.380 1906.140 1207.640 ;
        RECT 1905.420 1173.380 1905.680 1173.640 ;
        RECT 1905.880 1159.100 1906.140 1159.360 ;
        RECT 1905.880 1124.760 1906.140 1125.020 ;
        RECT 1905.880 1110.820 1906.140 1111.080 ;
        RECT 1905.420 1076.820 1905.680 1077.080 ;
        RECT 1905.880 1062.540 1906.140 1062.800 ;
        RECT 1905.880 1028.200 1906.140 1028.460 ;
        RECT 1905.880 1027.520 1906.140 1027.780 ;
        RECT 1905.420 1007.120 1905.680 1007.380 ;
        RECT 1906.800 1007.120 1907.060 1007.380 ;
        RECT 1905.880 917.700 1906.140 917.960 ;
        RECT 1906.800 917.700 1907.060 917.960 ;
        RECT 1904.040 869.420 1904.300 869.680 ;
        RECT 1904.960 869.420 1905.220 869.680 ;
        RECT 1904.960 820.460 1905.220 820.720 ;
        RECT 1905.420 820.460 1905.680 820.720 ;
        RECT 1904.960 814.000 1905.220 814.260 ;
        RECT 1905.420 737.840 1905.680 738.100 ;
        RECT 1905.420 676.300 1905.680 676.560 ;
        RECT 1906.340 676.300 1906.600 676.560 ;
        RECT 1905.420 641.620 1905.680 641.880 ;
        RECT 1905.880 641.280 1906.140 641.540 ;
        RECT 1905.420 579.400 1905.680 579.660 ;
        RECT 1906.340 579.400 1906.600 579.660 ;
        RECT 1905.420 386.280 1905.680 386.540 ;
        RECT 1905.880 386.280 1906.140 386.540 ;
        RECT 1905.880 241.100 1906.140 241.360 ;
        RECT 1906.340 241.100 1906.600 241.360 ;
        RECT 1905.880 144.880 1906.140 145.140 ;
        RECT 1906.340 144.880 1906.600 145.140 ;
        RECT 1905.420 96.600 1905.680 96.860 ;
        RECT 1906.340 96.600 1906.600 96.860 ;
        RECT 1905.420 89.460 1905.680 89.720 ;
        RECT 1904.960 41.520 1905.220 41.780 ;
        RECT 1594.000 33.360 1594.260 33.620 ;
        RECT 1904.960 33.360 1905.220 33.620 ;
        RECT 1477.620 16.700 1477.880 16.960 ;
        RECT 1594.000 16.700 1594.260 16.960 ;
      LAYER met2 ;
        RECT 1909.020 1700.410 1909.300 1702.400 ;
        RECT 1906.860 1700.270 1909.300 1700.410 ;
        RECT 1906.860 1683.670 1907.000 1700.270 ;
        RECT 1909.020 1700.000 1909.300 1700.270 ;
        RECT 1904.960 1683.350 1905.220 1683.670 ;
        RECT 1906.800 1683.350 1907.060 1683.670 ;
        RECT 1905.020 1641.930 1905.160 1683.350 ;
        RECT 1905.020 1641.790 1905.620 1641.930 ;
        RECT 1905.480 1593.910 1905.620 1641.790 ;
        RECT 1905.420 1593.590 1905.680 1593.910 ;
        RECT 1906.340 1593.590 1906.600 1593.910 ;
        RECT 1906.400 1587.110 1906.540 1593.590 ;
        RECT 1906.340 1586.790 1906.600 1587.110 ;
        RECT 1906.340 1538.850 1906.600 1539.170 ;
        RECT 1906.400 1521.570 1906.540 1538.850 ;
        RECT 1906.400 1521.430 1907.000 1521.570 ;
        RECT 1906.860 1449.410 1907.000 1521.430 ;
        RECT 1905.420 1449.090 1905.680 1449.410 ;
        RECT 1906.800 1449.090 1907.060 1449.410 ;
        RECT 1905.480 1414.730 1905.620 1449.090 ;
        RECT 1905.420 1414.410 1905.680 1414.730 ;
        RECT 1905.880 1413.730 1906.140 1414.050 ;
        RECT 1905.940 1400.530 1906.080 1413.730 ;
        RECT 1905.020 1400.390 1906.080 1400.530 ;
        RECT 1905.020 1352.850 1905.160 1400.390 ;
        RECT 1904.960 1352.530 1905.220 1352.850 ;
        RECT 1905.420 1352.530 1905.680 1352.850 ;
        RECT 1905.480 1352.170 1905.620 1352.530 ;
        RECT 1905.420 1351.850 1905.680 1352.170 ;
        RECT 1905.880 1304.250 1906.140 1304.570 ;
        RECT 1905.940 1304.085 1906.080 1304.250 ;
        RECT 1905.870 1303.715 1906.150 1304.085 ;
        RECT 1906.790 1303.715 1907.070 1304.085 ;
        RECT 1906.860 1256.290 1907.000 1303.715 ;
        RECT 1905.420 1255.970 1905.680 1256.290 ;
        RECT 1906.800 1255.970 1907.060 1256.290 ;
        RECT 1905.480 1255.610 1905.620 1255.970 ;
        RECT 1905.420 1255.290 1905.680 1255.610 ;
        RECT 1905.940 1207.670 1906.080 1207.825 ;
        RECT 1905.880 1207.410 1906.140 1207.670 ;
        RECT 1905.480 1207.350 1906.140 1207.410 ;
        RECT 1905.480 1207.270 1906.080 1207.350 ;
        RECT 1905.480 1173.670 1905.620 1207.270 ;
        RECT 1905.420 1173.350 1905.680 1173.670 ;
        RECT 1905.880 1159.070 1906.140 1159.390 ;
        RECT 1905.940 1125.050 1906.080 1159.070 ;
        RECT 1905.880 1124.730 1906.140 1125.050 ;
        RECT 1905.940 1111.110 1906.080 1111.265 ;
        RECT 1905.880 1110.850 1906.140 1111.110 ;
        RECT 1905.480 1110.790 1906.140 1110.850 ;
        RECT 1905.480 1110.710 1906.080 1110.790 ;
        RECT 1905.480 1077.110 1905.620 1110.710 ;
        RECT 1905.420 1076.790 1905.680 1077.110 ;
        RECT 1905.880 1062.510 1906.140 1062.830 ;
        RECT 1905.940 1028.490 1906.080 1062.510 ;
        RECT 1905.880 1028.170 1906.140 1028.490 ;
        RECT 1905.880 1027.490 1906.140 1027.810 ;
        RECT 1905.940 1014.290 1906.080 1027.490 ;
        RECT 1905.480 1014.150 1906.080 1014.290 ;
        RECT 1905.480 1007.410 1905.620 1014.150 ;
        RECT 1905.420 1007.090 1905.680 1007.410 ;
        RECT 1906.800 1007.090 1907.060 1007.410 ;
        RECT 1905.940 917.990 1906.080 918.145 ;
        RECT 1906.860 917.990 1907.000 1007.090 ;
        RECT 1904.030 917.475 1904.310 917.845 ;
        RECT 1905.410 917.730 1905.690 917.845 ;
        RECT 1905.880 917.730 1906.140 917.990 ;
        RECT 1905.410 917.670 1906.140 917.730 ;
        RECT 1906.800 917.670 1907.060 917.990 ;
        RECT 1905.410 917.590 1906.080 917.670 ;
        RECT 1905.410 917.475 1905.690 917.590 ;
        RECT 1904.100 869.710 1904.240 917.475 ;
        RECT 1904.040 869.390 1904.300 869.710 ;
        RECT 1904.960 869.390 1905.220 869.710 ;
        RECT 1905.020 856.530 1905.160 869.390 ;
        RECT 1905.020 856.390 1905.620 856.530 ;
        RECT 1905.480 820.750 1905.620 856.390 ;
        RECT 1904.960 820.430 1905.220 820.750 ;
        RECT 1905.420 820.430 1905.680 820.750 ;
        RECT 1905.020 814.290 1905.160 820.430 ;
        RECT 1904.960 813.970 1905.220 814.290 ;
        RECT 1905.420 737.810 1905.680 738.130 ;
        RECT 1905.480 724.610 1905.620 737.810 ;
        RECT 1905.480 724.470 1906.080 724.610 ;
        RECT 1905.940 724.440 1906.080 724.470 ;
        RECT 1905.940 724.300 1906.540 724.440 ;
        RECT 1906.400 676.590 1906.540 724.300 ;
        RECT 1905.420 676.270 1905.680 676.590 ;
        RECT 1906.340 676.270 1906.600 676.590 ;
        RECT 1905.480 641.910 1905.620 676.270 ;
        RECT 1905.420 641.590 1905.680 641.910 ;
        RECT 1905.880 641.250 1906.140 641.570 ;
        RECT 1905.940 627.880 1906.080 641.250 ;
        RECT 1905.940 627.740 1906.540 627.880 ;
        RECT 1906.400 580.565 1906.540 627.740 ;
        RECT 1906.330 580.195 1906.610 580.565 ;
        RECT 1905.410 579.515 1905.690 579.885 ;
        RECT 1905.420 579.370 1905.680 579.515 ;
        RECT 1906.340 579.370 1906.600 579.690 ;
        RECT 1906.400 483.210 1906.540 579.370 ;
        RECT 1905.940 483.070 1906.540 483.210 ;
        RECT 1905.940 386.570 1906.080 483.070 ;
        RECT 1905.420 386.250 1905.680 386.570 ;
        RECT 1905.880 386.250 1906.140 386.570 ;
        RECT 1905.480 254.730 1905.620 386.250 ;
        RECT 1905.480 254.590 1906.080 254.730 ;
        RECT 1905.940 241.390 1906.080 254.590 ;
        RECT 1905.880 241.070 1906.140 241.390 ;
        RECT 1906.340 241.070 1906.600 241.390 ;
        RECT 1906.400 145.170 1906.540 241.070 ;
        RECT 1905.880 144.850 1906.140 145.170 ;
        RECT 1906.340 144.850 1906.600 145.170 ;
        RECT 1905.940 98.330 1906.080 144.850 ;
        RECT 1905.940 98.190 1906.540 98.330 ;
        RECT 1906.400 96.890 1906.540 98.190 ;
        RECT 1905.420 96.570 1905.680 96.890 ;
        RECT 1906.340 96.570 1906.600 96.890 ;
        RECT 1905.480 89.750 1905.620 96.570 ;
        RECT 1905.420 89.430 1905.680 89.750 ;
        RECT 1904.960 41.490 1905.220 41.810 ;
        RECT 1905.020 33.650 1905.160 41.490 ;
        RECT 1594.000 33.330 1594.260 33.650 ;
        RECT 1904.960 33.330 1905.220 33.650 ;
        RECT 1594.060 16.990 1594.200 33.330 ;
        RECT 1477.620 16.670 1477.880 16.990 ;
        RECT 1594.000 16.670 1594.260 16.990 ;
        RECT 1477.680 2.400 1477.820 16.670 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
      LAYER via2 ;
        RECT 1905.870 1303.760 1906.150 1304.040 ;
        RECT 1906.790 1303.760 1907.070 1304.040 ;
        RECT 1904.030 917.520 1904.310 917.800 ;
        RECT 1905.410 917.520 1905.690 917.800 ;
        RECT 1906.330 580.240 1906.610 580.520 ;
        RECT 1905.410 579.560 1905.690 579.840 ;
      LAYER met3 ;
        RECT 1905.845 1304.050 1906.175 1304.065 ;
        RECT 1906.765 1304.050 1907.095 1304.065 ;
        RECT 1905.845 1303.750 1907.095 1304.050 ;
        RECT 1905.845 1303.735 1906.175 1303.750 ;
        RECT 1906.765 1303.735 1907.095 1303.750 ;
        RECT 1904.005 917.810 1904.335 917.825 ;
        RECT 1905.385 917.810 1905.715 917.825 ;
        RECT 1904.005 917.510 1905.715 917.810 ;
        RECT 1904.005 917.495 1904.335 917.510 ;
        RECT 1905.385 917.495 1905.715 917.510 ;
        RECT 1906.305 580.530 1906.635 580.545 ;
        RECT 1905.630 580.230 1906.635 580.530 ;
        RECT 1905.630 579.865 1905.930 580.230 ;
        RECT 1906.305 580.215 1906.635 580.230 ;
        RECT 1905.385 579.550 1905.930 579.865 ;
        RECT 1905.385 579.535 1905.715 579.550 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1504.730 51.920 1505.050 51.980 ;
        RECT 1918.730 51.920 1919.050 51.980 ;
        RECT 1504.730 51.780 1919.050 51.920 ;
        RECT 1504.730 51.720 1505.050 51.780 ;
        RECT 1918.730 51.720 1919.050 51.780 ;
        RECT 1495.530 18.600 1495.850 18.660 ;
        RECT 1504.730 18.600 1505.050 18.660 ;
        RECT 1495.530 18.460 1505.050 18.600 ;
        RECT 1495.530 18.400 1495.850 18.460 ;
        RECT 1504.730 18.400 1505.050 18.460 ;
      LAYER via ;
        RECT 1504.760 51.720 1505.020 51.980 ;
        RECT 1918.760 51.720 1919.020 51.980 ;
        RECT 1495.560 18.400 1495.820 18.660 ;
        RECT 1504.760 18.400 1505.020 18.660 ;
      LAYER met2 ;
        RECT 1918.220 1700.410 1918.500 1702.400 ;
        RECT 1918.220 1700.270 1918.960 1700.410 ;
        RECT 1918.220 1700.000 1918.500 1700.270 ;
        RECT 1918.820 52.010 1918.960 1700.270 ;
        RECT 1504.760 51.690 1505.020 52.010 ;
        RECT 1918.760 51.690 1919.020 52.010 ;
        RECT 1504.820 18.690 1504.960 51.690 ;
        RECT 1495.560 18.370 1495.820 18.690 ;
        RECT 1504.760 18.370 1505.020 18.690 ;
        RECT 1495.620 2.400 1495.760 18.370 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1600.870 33.220 1601.190 33.280 ;
        RECT 1925.630 33.220 1925.950 33.280 ;
        RECT 1600.870 33.080 1925.950 33.220 ;
        RECT 1600.870 33.020 1601.190 33.080 ;
        RECT 1925.630 33.020 1925.950 33.080 ;
        RECT 1513.010 16.220 1513.330 16.280 ;
        RECT 1600.870 16.220 1601.190 16.280 ;
        RECT 1513.010 16.080 1601.190 16.220 ;
        RECT 1513.010 16.020 1513.330 16.080 ;
        RECT 1600.870 16.020 1601.190 16.080 ;
      LAYER via ;
        RECT 1600.900 33.020 1601.160 33.280 ;
        RECT 1925.660 33.020 1925.920 33.280 ;
        RECT 1513.040 16.020 1513.300 16.280 ;
        RECT 1600.900 16.020 1601.160 16.280 ;
      LAYER met2 ;
        RECT 1927.420 1700.410 1927.700 1702.400 ;
        RECT 1925.720 1700.270 1927.700 1700.410 ;
        RECT 1925.720 33.310 1925.860 1700.270 ;
        RECT 1927.420 1700.000 1927.700 1700.270 ;
        RECT 1600.900 32.990 1601.160 33.310 ;
        RECT 1925.660 32.990 1925.920 33.310 ;
        RECT 1600.960 16.310 1601.100 32.990 ;
        RECT 1513.040 15.990 1513.300 16.310 ;
        RECT 1600.900 15.990 1601.160 16.310 ;
        RECT 1513.100 2.400 1513.240 15.990 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 709.850 36.280 710.170 36.340 ;
        RECT 1512.550 36.280 1512.870 36.340 ;
        RECT 709.850 36.140 1512.870 36.280 ;
        RECT 709.850 36.080 710.170 36.140 ;
        RECT 1512.550 36.080 1512.870 36.140 ;
      LAYER via ;
        RECT 709.880 36.080 710.140 36.340 ;
        RECT 1512.580 36.080 1512.840 36.340 ;
      LAYER met2 ;
        RECT 1513.880 1700.410 1514.160 1702.400 ;
        RECT 1512.640 1700.270 1514.160 1700.410 ;
        RECT 1512.640 36.370 1512.780 1700.270 ;
        RECT 1513.880 1700.000 1514.160 1700.270 ;
        RECT 709.880 36.050 710.140 36.370 ;
        RECT 1512.580 36.050 1512.840 36.370 ;
        RECT 709.940 17.410 710.080 36.050 ;
        RECT 709.940 17.270 710.540 17.410 ;
        RECT 710.400 2.400 710.540 17.270 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1933.065 855.525 1933.235 903.975 ;
        RECT 1933.065 386.325 1933.235 434.435 ;
      LAYER mcon ;
        RECT 1933.065 903.805 1933.235 903.975 ;
        RECT 1933.065 434.265 1933.235 434.435 ;
      LAYER met1 ;
        RECT 1933.450 1400.700 1933.770 1400.760 ;
        RECT 1933.910 1400.700 1934.230 1400.760 ;
        RECT 1933.450 1400.560 1934.230 1400.700 ;
        RECT 1933.450 1400.500 1933.770 1400.560 ;
        RECT 1933.910 1400.500 1934.230 1400.560 ;
        RECT 1932.990 1249.400 1933.310 1249.460 ;
        RECT 1933.450 1249.400 1933.770 1249.460 ;
        RECT 1932.990 1249.260 1933.770 1249.400 ;
        RECT 1932.990 1249.200 1933.310 1249.260 ;
        RECT 1933.450 1249.200 1933.770 1249.260 ;
        RECT 1933.450 1221.520 1933.770 1221.580 ;
        RECT 1933.080 1221.380 1933.770 1221.520 ;
        RECT 1933.080 1221.240 1933.220 1221.380 ;
        RECT 1933.450 1221.320 1933.770 1221.380 ;
        RECT 1932.990 1220.980 1933.310 1221.240 ;
        RECT 1932.990 1124.760 1933.310 1125.020 ;
        RECT 1933.080 1124.280 1933.220 1124.760 ;
        RECT 1933.450 1124.280 1933.770 1124.340 ;
        RECT 1933.080 1124.140 1933.770 1124.280 ;
        RECT 1933.450 1124.080 1933.770 1124.140 ;
        RECT 1932.990 966.520 1933.310 966.580 ;
        RECT 1933.910 966.520 1934.230 966.580 ;
        RECT 1932.990 966.380 1934.230 966.520 ;
        RECT 1932.990 966.320 1933.310 966.380 ;
        RECT 1933.910 966.320 1934.230 966.380 ;
        RECT 1933.450 911.100 1933.770 911.160 ;
        RECT 1933.910 911.100 1934.230 911.160 ;
        RECT 1933.450 910.960 1934.230 911.100 ;
        RECT 1933.450 910.900 1933.770 910.960 ;
        RECT 1933.910 910.900 1934.230 910.960 ;
        RECT 1933.005 903.960 1933.295 904.005 ;
        RECT 1933.450 903.960 1933.770 904.020 ;
        RECT 1933.005 903.820 1933.770 903.960 ;
        RECT 1933.005 903.775 1933.295 903.820 ;
        RECT 1933.450 903.760 1933.770 903.820 ;
        RECT 1932.990 855.680 1933.310 855.740 ;
        RECT 1932.795 855.540 1933.310 855.680 ;
        RECT 1932.990 855.480 1933.310 855.540 ;
        RECT 1932.990 814.200 1933.310 814.260 ;
        RECT 1933.910 814.200 1934.230 814.260 ;
        RECT 1932.990 814.060 1934.230 814.200 ;
        RECT 1932.990 814.000 1933.310 814.060 ;
        RECT 1933.910 814.000 1934.230 814.060 ;
        RECT 1933.450 627.880 1933.770 627.940 ;
        RECT 1933.910 627.880 1934.230 627.940 ;
        RECT 1933.450 627.740 1934.230 627.880 ;
        RECT 1933.450 627.680 1933.770 627.740 ;
        RECT 1933.910 627.680 1934.230 627.740 ;
        RECT 1932.990 579.600 1933.310 579.660 ;
        RECT 1933.910 579.600 1934.230 579.660 ;
        RECT 1932.990 579.460 1934.230 579.600 ;
        RECT 1932.990 579.400 1933.310 579.460 ;
        RECT 1933.910 579.400 1934.230 579.460 ;
        RECT 1932.990 434.420 1933.310 434.480 ;
        RECT 1932.795 434.280 1933.310 434.420 ;
        RECT 1932.990 434.220 1933.310 434.280 ;
        RECT 1932.990 386.480 1933.310 386.540 ;
        RECT 1932.795 386.340 1933.310 386.480 ;
        RECT 1932.990 386.280 1933.310 386.340 ;
        RECT 1932.990 338.340 1933.310 338.600 ;
        RECT 1933.080 338.200 1933.220 338.340 ;
        RECT 1933.450 338.200 1933.770 338.260 ;
        RECT 1933.080 338.060 1933.770 338.200 ;
        RECT 1933.450 338.000 1933.770 338.060 ;
        RECT 1932.990 289.920 1933.310 289.980 ;
        RECT 1933.450 289.920 1933.770 289.980 ;
        RECT 1932.990 289.780 1933.770 289.920 ;
        RECT 1932.990 289.720 1933.310 289.780 ;
        RECT 1933.450 289.720 1933.770 289.780 ;
        RECT 1932.990 241.640 1933.310 241.700 ;
        RECT 1933.450 241.640 1933.770 241.700 ;
        RECT 1932.990 241.500 1933.770 241.640 ;
        RECT 1932.990 241.440 1933.310 241.500 ;
        RECT 1933.450 241.440 1933.770 241.500 ;
        RECT 1933.450 186.700 1933.770 186.960 ;
        RECT 1933.540 186.560 1933.680 186.700 ;
        RECT 1933.910 186.560 1934.230 186.620 ;
        RECT 1933.540 186.420 1934.230 186.560 ;
        RECT 1933.910 186.360 1934.230 186.420 ;
        RECT 1933.450 145.080 1933.770 145.140 ;
        RECT 1933.450 144.940 1934.140 145.080 ;
        RECT 1933.450 144.880 1933.770 144.940 ;
        RECT 1934.000 144.460 1934.140 144.940 ;
        RECT 1933.910 144.200 1934.230 144.460 ;
        RECT 1933.910 94.900 1934.230 95.160 ;
        RECT 1934.000 94.480 1934.140 94.900 ;
        RECT 1933.910 94.220 1934.230 94.480 ;
        RECT 1932.530 48.520 1932.850 48.580 ;
        RECT 1933.910 48.520 1934.230 48.580 ;
        RECT 1932.530 48.380 1934.230 48.520 ;
        RECT 1932.530 48.320 1932.850 48.380 ;
        RECT 1933.910 48.320 1934.230 48.380 ;
        RECT 1628.010 33.900 1628.330 33.960 ;
        RECT 1932.530 33.900 1932.850 33.960 ;
        RECT 1628.010 33.760 1932.850 33.900 ;
        RECT 1628.010 33.700 1628.330 33.760 ;
        RECT 1932.530 33.700 1932.850 33.760 ;
        RECT 1530.950 16.560 1531.270 16.620 ;
        RECT 1628.010 16.560 1628.330 16.620 ;
        RECT 1530.950 16.420 1628.330 16.560 ;
        RECT 1530.950 16.360 1531.270 16.420 ;
        RECT 1628.010 16.360 1628.330 16.420 ;
      LAYER via ;
        RECT 1933.480 1400.500 1933.740 1400.760 ;
        RECT 1933.940 1400.500 1934.200 1400.760 ;
        RECT 1933.020 1249.200 1933.280 1249.460 ;
        RECT 1933.480 1249.200 1933.740 1249.460 ;
        RECT 1933.480 1221.320 1933.740 1221.580 ;
        RECT 1933.020 1220.980 1933.280 1221.240 ;
        RECT 1933.020 1124.760 1933.280 1125.020 ;
        RECT 1933.480 1124.080 1933.740 1124.340 ;
        RECT 1933.020 966.320 1933.280 966.580 ;
        RECT 1933.940 966.320 1934.200 966.580 ;
        RECT 1933.480 910.900 1933.740 911.160 ;
        RECT 1933.940 910.900 1934.200 911.160 ;
        RECT 1933.480 903.760 1933.740 904.020 ;
        RECT 1933.020 855.480 1933.280 855.740 ;
        RECT 1933.020 814.000 1933.280 814.260 ;
        RECT 1933.940 814.000 1934.200 814.260 ;
        RECT 1933.480 627.680 1933.740 627.940 ;
        RECT 1933.940 627.680 1934.200 627.940 ;
        RECT 1933.020 579.400 1933.280 579.660 ;
        RECT 1933.940 579.400 1934.200 579.660 ;
        RECT 1933.020 434.220 1933.280 434.480 ;
        RECT 1933.020 386.280 1933.280 386.540 ;
        RECT 1933.020 338.340 1933.280 338.600 ;
        RECT 1933.480 338.000 1933.740 338.260 ;
        RECT 1933.020 289.720 1933.280 289.980 ;
        RECT 1933.480 289.720 1933.740 289.980 ;
        RECT 1933.020 241.440 1933.280 241.700 ;
        RECT 1933.480 241.440 1933.740 241.700 ;
        RECT 1933.480 186.700 1933.740 186.960 ;
        RECT 1933.940 186.360 1934.200 186.620 ;
        RECT 1933.480 144.880 1933.740 145.140 ;
        RECT 1933.940 144.200 1934.200 144.460 ;
        RECT 1933.940 94.900 1934.200 95.160 ;
        RECT 1933.940 94.220 1934.200 94.480 ;
        RECT 1932.560 48.320 1932.820 48.580 ;
        RECT 1933.940 48.320 1934.200 48.580 ;
        RECT 1628.040 33.700 1628.300 33.960 ;
        RECT 1932.560 33.700 1932.820 33.960 ;
        RECT 1530.980 16.360 1531.240 16.620 ;
        RECT 1628.040 16.360 1628.300 16.620 ;
      LAYER met2 ;
        RECT 1936.620 1700.410 1936.900 1702.400 ;
        RECT 1934.460 1700.270 1936.900 1700.410 ;
        RECT 1934.460 1656.210 1934.600 1700.270 ;
        RECT 1936.620 1700.000 1936.900 1700.270 ;
        RECT 1933.080 1656.070 1934.600 1656.210 ;
        RECT 1933.080 1655.530 1933.220 1656.070 ;
        RECT 1933.080 1655.390 1933.680 1655.530 ;
        RECT 1933.540 1606.570 1933.680 1655.390 ;
        RECT 1933.080 1606.430 1933.680 1606.570 ;
        RECT 1933.080 1593.650 1933.220 1606.430 ;
        RECT 1933.080 1593.510 1933.680 1593.650 ;
        RECT 1933.540 1463.090 1933.680 1593.510 ;
        RECT 1933.080 1462.950 1933.680 1463.090 ;
        RECT 1933.080 1425.010 1933.220 1462.950 ;
        RECT 1933.080 1424.870 1934.140 1425.010 ;
        RECT 1934.000 1414.130 1934.140 1424.870 ;
        RECT 1933.540 1413.990 1934.140 1414.130 ;
        RECT 1933.540 1400.790 1933.680 1413.990 ;
        RECT 1933.480 1400.470 1933.740 1400.790 ;
        RECT 1933.940 1400.470 1934.200 1400.790 ;
        RECT 1934.000 1353.045 1934.140 1400.470 ;
        RECT 1933.930 1352.675 1934.210 1353.045 ;
        RECT 1933.470 1351.995 1933.750 1352.365 ;
        RECT 1933.540 1249.490 1933.680 1351.995 ;
        RECT 1933.020 1249.170 1933.280 1249.490 ;
        RECT 1933.480 1249.170 1933.740 1249.490 ;
        RECT 1933.080 1248.890 1933.220 1249.170 ;
        RECT 1933.080 1248.750 1933.680 1248.890 ;
        RECT 1933.540 1221.610 1933.680 1248.750 ;
        RECT 1933.480 1221.290 1933.740 1221.610 ;
        RECT 1933.020 1220.950 1933.280 1221.270 ;
        RECT 1933.080 1125.050 1933.220 1220.950 ;
        RECT 1933.020 1124.730 1933.280 1125.050 ;
        RECT 1933.480 1124.050 1933.740 1124.370 ;
        RECT 1933.540 1087.050 1933.680 1124.050 ;
        RECT 1933.080 1086.910 1933.680 1087.050 ;
        RECT 1933.080 1062.685 1933.220 1086.910 ;
        RECT 1933.010 1062.315 1933.290 1062.685 ;
        RECT 1933.930 1062.315 1934.210 1062.685 ;
        RECT 1934.000 966.610 1934.140 1062.315 ;
        RECT 1933.020 966.290 1933.280 966.610 ;
        RECT 1933.940 966.290 1934.200 966.610 ;
        RECT 1933.080 966.125 1933.220 966.290 ;
        RECT 1933.010 965.755 1933.290 966.125 ;
        RECT 1933.930 965.755 1934.210 966.125 ;
        RECT 1934.000 911.190 1934.140 965.755 ;
        RECT 1933.480 910.870 1933.740 911.190 ;
        RECT 1933.940 910.870 1934.200 911.190 ;
        RECT 1933.540 904.050 1933.680 910.870 ;
        RECT 1933.480 903.730 1933.740 904.050 ;
        RECT 1933.020 855.450 1933.280 855.770 ;
        RECT 1933.080 814.290 1933.220 855.450 ;
        RECT 1933.020 813.970 1933.280 814.290 ;
        RECT 1933.940 813.970 1934.200 814.290 ;
        RECT 1934.000 676.445 1934.140 813.970 ;
        RECT 1933.010 676.075 1933.290 676.445 ;
        RECT 1933.930 676.075 1934.210 676.445 ;
        RECT 1933.080 651.850 1933.220 676.075 ;
        RECT 1933.080 651.710 1933.680 651.850 ;
        RECT 1933.540 627.970 1933.680 651.710 ;
        RECT 1933.480 627.650 1933.740 627.970 ;
        RECT 1933.940 627.650 1934.200 627.970 ;
        RECT 1934.000 579.885 1934.140 627.650 ;
        RECT 1933.010 579.515 1933.290 579.885 ;
        RECT 1933.930 579.515 1934.210 579.885 ;
        RECT 1933.020 579.370 1933.280 579.515 ;
        RECT 1933.940 579.370 1934.200 579.515 ;
        RECT 1934.000 483.325 1934.140 579.370 ;
        RECT 1933.010 482.955 1933.290 483.325 ;
        RECT 1933.930 482.955 1934.210 483.325 ;
        RECT 1933.080 434.510 1933.220 482.955 ;
        RECT 1933.020 434.190 1933.280 434.510 ;
        RECT 1933.020 386.250 1933.280 386.570 ;
        RECT 1933.080 338.630 1933.220 386.250 ;
        RECT 1933.020 338.310 1933.280 338.630 ;
        RECT 1933.480 337.970 1933.740 338.290 ;
        RECT 1933.540 290.010 1933.680 337.970 ;
        RECT 1933.020 289.690 1933.280 290.010 ;
        RECT 1933.480 289.690 1933.740 290.010 ;
        RECT 1933.080 241.730 1933.220 289.690 ;
        RECT 1933.020 241.410 1933.280 241.730 ;
        RECT 1933.480 241.410 1933.740 241.730 ;
        RECT 1933.540 186.990 1933.680 241.410 ;
        RECT 1933.480 186.670 1933.740 186.990 ;
        RECT 1933.940 186.330 1934.200 186.650 ;
        RECT 1934.000 186.050 1934.140 186.330 ;
        RECT 1933.540 185.910 1934.140 186.050 ;
        RECT 1933.540 145.170 1933.680 185.910 ;
        RECT 1933.480 144.850 1933.740 145.170 ;
        RECT 1933.940 144.170 1934.200 144.490 ;
        RECT 1934.000 95.190 1934.140 144.170 ;
        RECT 1933.940 94.870 1934.200 95.190 ;
        RECT 1933.940 94.190 1934.200 94.510 ;
        RECT 1934.000 48.610 1934.140 94.190 ;
        RECT 1932.560 48.290 1932.820 48.610 ;
        RECT 1933.940 48.290 1934.200 48.610 ;
        RECT 1932.620 33.990 1932.760 48.290 ;
        RECT 1628.040 33.670 1628.300 33.990 ;
        RECT 1932.560 33.670 1932.820 33.990 ;
        RECT 1628.100 16.650 1628.240 33.670 ;
        RECT 1530.980 16.330 1531.240 16.650 ;
        RECT 1628.040 16.330 1628.300 16.650 ;
        RECT 1531.040 2.400 1531.180 16.330 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
      LAYER via2 ;
        RECT 1933.930 1352.720 1934.210 1353.000 ;
        RECT 1933.470 1352.040 1933.750 1352.320 ;
        RECT 1933.010 1062.360 1933.290 1062.640 ;
        RECT 1933.930 1062.360 1934.210 1062.640 ;
        RECT 1933.010 965.800 1933.290 966.080 ;
        RECT 1933.930 965.800 1934.210 966.080 ;
        RECT 1933.010 676.120 1933.290 676.400 ;
        RECT 1933.930 676.120 1934.210 676.400 ;
        RECT 1933.010 579.560 1933.290 579.840 ;
        RECT 1933.930 579.560 1934.210 579.840 ;
        RECT 1933.010 483.000 1933.290 483.280 ;
        RECT 1933.930 483.000 1934.210 483.280 ;
      LAYER met3 ;
        RECT 1933.905 1353.010 1934.235 1353.025 ;
        RECT 1933.230 1352.710 1934.235 1353.010 ;
        RECT 1933.230 1352.345 1933.530 1352.710 ;
        RECT 1933.905 1352.695 1934.235 1352.710 ;
        RECT 1933.230 1352.030 1933.775 1352.345 ;
        RECT 1933.445 1352.015 1933.775 1352.030 ;
        RECT 1932.985 1062.650 1933.315 1062.665 ;
        RECT 1933.905 1062.650 1934.235 1062.665 ;
        RECT 1932.985 1062.350 1934.235 1062.650 ;
        RECT 1932.985 1062.335 1933.315 1062.350 ;
        RECT 1933.905 1062.335 1934.235 1062.350 ;
        RECT 1932.985 966.090 1933.315 966.105 ;
        RECT 1933.905 966.090 1934.235 966.105 ;
        RECT 1932.985 965.790 1934.235 966.090 ;
        RECT 1932.985 965.775 1933.315 965.790 ;
        RECT 1933.905 965.775 1934.235 965.790 ;
        RECT 1932.985 676.410 1933.315 676.425 ;
        RECT 1933.905 676.410 1934.235 676.425 ;
        RECT 1932.985 676.110 1934.235 676.410 ;
        RECT 1932.985 676.095 1933.315 676.110 ;
        RECT 1933.905 676.095 1934.235 676.110 ;
        RECT 1932.985 579.850 1933.315 579.865 ;
        RECT 1933.905 579.850 1934.235 579.865 ;
        RECT 1932.985 579.550 1934.235 579.850 ;
        RECT 1932.985 579.535 1933.315 579.550 ;
        RECT 1933.905 579.535 1934.235 579.550 ;
        RECT 1932.985 483.290 1933.315 483.305 ;
        RECT 1933.905 483.290 1934.235 483.305 ;
        RECT 1932.985 482.990 1934.235 483.290 ;
        RECT 1932.985 482.975 1933.315 482.990 ;
        RECT 1933.905 482.975 1934.235 482.990 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1617.890 45.120 1618.210 45.180 ;
        RECT 1946.330 45.120 1946.650 45.180 ;
        RECT 1617.890 44.980 1946.650 45.120 ;
        RECT 1617.890 44.920 1618.210 44.980 ;
        RECT 1946.330 44.920 1946.650 44.980 ;
        RECT 1548.890 15.880 1549.210 15.940 ;
        RECT 1617.890 15.880 1618.210 15.940 ;
        RECT 1548.890 15.740 1618.210 15.880 ;
        RECT 1548.890 15.680 1549.210 15.740 ;
        RECT 1617.890 15.680 1618.210 15.740 ;
      LAYER via ;
        RECT 1617.920 44.920 1618.180 45.180 ;
        RECT 1946.360 44.920 1946.620 45.180 ;
        RECT 1548.920 15.680 1549.180 15.940 ;
        RECT 1617.920 15.680 1618.180 15.940 ;
      LAYER met2 ;
        RECT 1945.820 1700.410 1946.100 1702.400 ;
        RECT 1945.820 1700.270 1946.560 1700.410 ;
        RECT 1945.820 1700.000 1946.100 1700.270 ;
        RECT 1946.420 45.210 1946.560 1700.270 ;
        RECT 1617.920 44.890 1618.180 45.210 ;
        RECT 1946.360 44.890 1946.620 45.210 ;
        RECT 1617.980 15.970 1618.120 44.890 ;
        RECT 1548.920 15.650 1549.180 15.970 ;
        RECT 1617.920 15.650 1618.180 15.970 ;
        RECT 1548.980 2.400 1549.120 15.650 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1627.550 45.800 1627.870 45.860 ;
        RECT 1953.230 45.800 1953.550 45.860 ;
        RECT 1627.550 45.660 1953.550 45.800 ;
        RECT 1627.550 45.600 1627.870 45.660 ;
        RECT 1953.230 45.600 1953.550 45.660 ;
        RECT 1566.830 15.540 1567.150 15.600 ;
        RECT 1627.550 15.540 1627.870 15.600 ;
        RECT 1566.830 15.400 1627.870 15.540 ;
        RECT 1566.830 15.340 1567.150 15.400 ;
        RECT 1627.550 15.340 1627.870 15.400 ;
      LAYER via ;
        RECT 1627.580 45.600 1627.840 45.860 ;
        RECT 1953.260 45.600 1953.520 45.860 ;
        RECT 1566.860 15.340 1567.120 15.600 ;
        RECT 1627.580 15.340 1627.840 15.600 ;
      LAYER met2 ;
        RECT 1955.020 1700.410 1955.300 1702.400 ;
        RECT 1953.320 1700.270 1955.300 1700.410 ;
        RECT 1953.320 45.890 1953.460 1700.270 ;
        RECT 1955.020 1700.000 1955.300 1700.270 ;
        RECT 1627.580 45.570 1627.840 45.890 ;
        RECT 1953.260 45.570 1953.520 45.890 ;
        RECT 1627.640 15.630 1627.780 45.570 ;
        RECT 1566.860 15.310 1567.120 15.630 ;
        RECT 1627.580 15.310 1627.840 15.630 ;
        RECT 1566.920 2.400 1567.060 15.310 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1960.665 1594.005 1960.835 1608.115 ;
        RECT 1960.665 1321.325 1960.835 1352.435 ;
        RECT 1960.665 1110.865 1960.835 1183.795 ;
        RECT 1960.665 855.525 1960.835 903.975 ;
        RECT 1960.665 676.345 1960.835 741.795 ;
        RECT 1960.665 386.325 1960.835 434.435 ;
        RECT 1960.665 235.025 1960.835 282.795 ;
      LAYER mcon ;
        RECT 1960.665 1607.945 1960.835 1608.115 ;
        RECT 1960.665 1352.265 1960.835 1352.435 ;
        RECT 1960.665 1183.625 1960.835 1183.795 ;
        RECT 1960.665 903.805 1960.835 903.975 ;
        RECT 1960.665 741.625 1960.835 741.795 ;
        RECT 1960.665 434.265 1960.835 434.435 ;
        RECT 1960.665 282.625 1960.835 282.795 ;
      LAYER met1 ;
        RECT 1960.605 1608.100 1960.895 1608.145 ;
        RECT 1961.050 1608.100 1961.370 1608.160 ;
        RECT 1960.605 1607.960 1961.370 1608.100 ;
        RECT 1960.605 1607.915 1960.895 1607.960 ;
        RECT 1961.050 1607.900 1961.370 1607.960 ;
        RECT 1960.590 1594.160 1960.910 1594.220 ;
        RECT 1960.395 1594.020 1960.910 1594.160 ;
        RECT 1960.590 1593.960 1960.910 1594.020 ;
        RECT 1960.590 1448.980 1960.910 1449.040 ;
        RECT 1961.050 1448.980 1961.370 1449.040 ;
        RECT 1960.590 1448.840 1961.370 1448.980 ;
        RECT 1960.590 1448.780 1960.910 1448.840 ;
        RECT 1961.050 1448.780 1961.370 1448.840 ;
        RECT 1960.590 1393.900 1960.910 1393.960 ;
        RECT 1961.050 1393.900 1961.370 1393.960 ;
        RECT 1960.590 1393.760 1961.370 1393.900 ;
        RECT 1960.590 1393.700 1960.910 1393.760 ;
        RECT 1961.050 1393.700 1961.370 1393.760 ;
        RECT 1960.590 1352.420 1960.910 1352.480 ;
        RECT 1960.395 1352.280 1960.910 1352.420 ;
        RECT 1960.590 1352.220 1960.910 1352.280 ;
        RECT 1960.605 1321.480 1960.895 1321.525 ;
        RECT 1961.050 1321.480 1961.370 1321.540 ;
        RECT 1960.605 1321.340 1961.370 1321.480 ;
        RECT 1960.605 1321.295 1960.895 1321.340 ;
        RECT 1961.050 1321.280 1961.370 1321.340 ;
        RECT 1960.590 1249.400 1960.910 1249.460 ;
        RECT 1961.050 1249.400 1961.370 1249.460 ;
        RECT 1960.590 1249.260 1961.370 1249.400 ;
        RECT 1960.590 1249.200 1960.910 1249.260 ;
        RECT 1961.050 1249.200 1961.370 1249.260 ;
        RECT 1961.050 1200.780 1961.370 1200.840 ;
        RECT 1961.970 1200.780 1962.290 1200.840 ;
        RECT 1961.050 1200.640 1962.290 1200.780 ;
        RECT 1961.050 1200.580 1961.370 1200.640 ;
        RECT 1961.970 1200.580 1962.290 1200.640 ;
        RECT 1960.605 1183.780 1960.895 1183.825 ;
        RECT 1961.050 1183.780 1961.370 1183.840 ;
        RECT 1960.605 1183.640 1961.370 1183.780 ;
        RECT 1960.605 1183.595 1960.895 1183.640 ;
        RECT 1961.050 1183.580 1961.370 1183.640 ;
        RECT 1960.605 1111.020 1960.895 1111.065 ;
        RECT 1961.050 1111.020 1961.370 1111.080 ;
        RECT 1960.605 1110.880 1961.370 1111.020 ;
        RECT 1960.605 1110.835 1960.895 1110.880 ;
        RECT 1961.050 1110.820 1961.370 1110.880 ;
        RECT 1960.130 976.380 1960.450 976.440 ;
        RECT 1961.510 976.380 1961.830 976.440 ;
        RECT 1960.130 976.240 1961.830 976.380 ;
        RECT 1960.130 976.180 1960.450 976.240 ;
        RECT 1961.510 976.180 1961.830 976.240 ;
        RECT 1960.605 903.960 1960.895 904.005 ;
        RECT 1961.050 903.960 1961.370 904.020 ;
        RECT 1960.605 903.820 1961.370 903.960 ;
        RECT 1960.605 903.775 1960.895 903.820 ;
        RECT 1961.050 903.760 1961.370 903.820 ;
        RECT 1960.590 855.680 1960.910 855.740 ;
        RECT 1960.395 855.540 1960.910 855.680 ;
        RECT 1960.590 855.480 1960.910 855.540 ;
        RECT 1960.590 814.200 1960.910 814.260 ;
        RECT 1961.510 814.200 1961.830 814.260 ;
        RECT 1960.590 814.060 1961.830 814.200 ;
        RECT 1960.590 814.000 1960.910 814.060 ;
        RECT 1961.510 814.000 1961.830 814.060 ;
        RECT 1960.605 741.780 1960.895 741.825 ;
        RECT 1961.510 741.780 1961.830 741.840 ;
        RECT 1960.605 741.640 1961.830 741.780 ;
        RECT 1960.605 741.595 1960.895 741.640 ;
        RECT 1961.510 741.580 1961.830 741.640 ;
        RECT 1960.590 676.500 1960.910 676.560 ;
        RECT 1960.395 676.360 1960.910 676.500 ;
        RECT 1960.590 676.300 1960.910 676.360 ;
        RECT 1961.050 627.880 1961.370 627.940 ;
        RECT 1961.510 627.880 1961.830 627.940 ;
        RECT 1961.050 627.740 1961.830 627.880 ;
        RECT 1961.050 627.680 1961.370 627.740 ;
        RECT 1961.510 627.680 1961.830 627.740 ;
        RECT 1960.590 579.600 1960.910 579.660 ;
        RECT 1961.510 579.600 1961.830 579.660 ;
        RECT 1960.590 579.460 1961.830 579.600 ;
        RECT 1960.590 579.400 1960.910 579.460 ;
        RECT 1961.510 579.400 1961.830 579.460 ;
        RECT 1960.590 434.420 1960.910 434.480 ;
        RECT 1960.395 434.280 1960.910 434.420 ;
        RECT 1960.590 434.220 1960.910 434.280 ;
        RECT 1960.590 386.480 1960.910 386.540 ;
        RECT 1960.395 386.340 1960.910 386.480 ;
        RECT 1960.590 386.280 1960.910 386.340 ;
        RECT 1960.590 338.340 1960.910 338.600 ;
        RECT 1960.680 338.200 1960.820 338.340 ;
        RECT 1961.050 338.200 1961.370 338.260 ;
        RECT 1960.680 338.060 1961.370 338.200 ;
        RECT 1961.050 338.000 1961.370 338.060 ;
        RECT 1961.050 308.620 1961.370 308.680 ;
        RECT 1961.970 308.620 1962.290 308.680 ;
        RECT 1961.050 308.480 1962.290 308.620 ;
        RECT 1961.050 308.420 1961.370 308.480 ;
        RECT 1961.970 308.420 1962.290 308.480 ;
        RECT 1960.605 282.780 1960.895 282.825 ;
        RECT 1961.510 282.780 1961.830 282.840 ;
        RECT 1960.605 282.640 1961.830 282.780 ;
        RECT 1960.605 282.595 1960.895 282.640 ;
        RECT 1961.510 282.580 1961.830 282.640 ;
        RECT 1960.590 235.180 1960.910 235.240 ;
        RECT 1960.395 235.040 1960.910 235.180 ;
        RECT 1960.590 234.980 1960.910 235.040 ;
        RECT 1960.590 234.300 1960.910 234.560 ;
        RECT 1960.680 233.880 1960.820 234.300 ;
        RECT 1960.590 233.620 1960.910 233.880 ;
        RECT 1960.130 144.740 1960.450 144.800 ;
        RECT 1961.050 144.740 1961.370 144.800 ;
        RECT 1960.130 144.600 1961.370 144.740 ;
        RECT 1960.130 144.540 1960.450 144.600 ;
        RECT 1961.050 144.540 1961.370 144.600 ;
        RECT 1635.370 46.140 1635.690 46.200 ;
        RECT 1960.130 46.140 1960.450 46.200 ;
        RECT 1635.370 46.000 1960.450 46.140 ;
        RECT 1635.370 45.940 1635.690 46.000 ;
        RECT 1960.130 45.940 1960.450 46.000 ;
        RECT 1584.770 19.280 1585.090 19.340 ;
        RECT 1635.370 19.280 1635.690 19.340 ;
        RECT 1584.770 19.140 1635.690 19.280 ;
        RECT 1584.770 19.080 1585.090 19.140 ;
        RECT 1635.370 19.080 1635.690 19.140 ;
      LAYER via ;
        RECT 1961.080 1607.900 1961.340 1608.160 ;
        RECT 1960.620 1593.960 1960.880 1594.220 ;
        RECT 1960.620 1448.780 1960.880 1449.040 ;
        RECT 1961.080 1448.780 1961.340 1449.040 ;
        RECT 1960.620 1393.700 1960.880 1393.960 ;
        RECT 1961.080 1393.700 1961.340 1393.960 ;
        RECT 1960.620 1352.220 1960.880 1352.480 ;
        RECT 1961.080 1321.280 1961.340 1321.540 ;
        RECT 1960.620 1249.200 1960.880 1249.460 ;
        RECT 1961.080 1249.200 1961.340 1249.460 ;
        RECT 1961.080 1200.580 1961.340 1200.840 ;
        RECT 1962.000 1200.580 1962.260 1200.840 ;
        RECT 1961.080 1183.580 1961.340 1183.840 ;
        RECT 1961.080 1110.820 1961.340 1111.080 ;
        RECT 1960.160 976.180 1960.420 976.440 ;
        RECT 1961.540 976.180 1961.800 976.440 ;
        RECT 1961.080 903.760 1961.340 904.020 ;
        RECT 1960.620 855.480 1960.880 855.740 ;
        RECT 1960.620 814.000 1960.880 814.260 ;
        RECT 1961.540 814.000 1961.800 814.260 ;
        RECT 1961.540 741.580 1961.800 741.840 ;
        RECT 1960.620 676.300 1960.880 676.560 ;
        RECT 1961.080 627.680 1961.340 627.940 ;
        RECT 1961.540 627.680 1961.800 627.940 ;
        RECT 1960.620 579.400 1960.880 579.660 ;
        RECT 1961.540 579.400 1961.800 579.660 ;
        RECT 1960.620 434.220 1960.880 434.480 ;
        RECT 1960.620 386.280 1960.880 386.540 ;
        RECT 1960.620 338.340 1960.880 338.600 ;
        RECT 1961.080 338.000 1961.340 338.260 ;
        RECT 1961.080 308.420 1961.340 308.680 ;
        RECT 1962.000 308.420 1962.260 308.680 ;
        RECT 1961.540 282.580 1961.800 282.840 ;
        RECT 1960.620 234.980 1960.880 235.240 ;
        RECT 1960.620 234.300 1960.880 234.560 ;
        RECT 1960.620 233.620 1960.880 233.880 ;
        RECT 1960.160 144.540 1960.420 144.800 ;
        RECT 1961.080 144.540 1961.340 144.800 ;
        RECT 1635.400 45.940 1635.660 46.200 ;
        RECT 1960.160 45.940 1960.420 46.200 ;
        RECT 1584.800 19.080 1585.060 19.340 ;
        RECT 1635.400 19.080 1635.660 19.340 ;
      LAYER met2 ;
        RECT 1964.220 1700.410 1964.500 1702.400 ;
        RECT 1962.060 1700.270 1964.500 1700.410 ;
        RECT 1962.060 1677.970 1962.200 1700.270 ;
        RECT 1964.220 1700.000 1964.500 1700.270 ;
        RECT 1960.680 1677.830 1962.200 1677.970 ;
        RECT 1960.680 1655.530 1960.820 1677.830 ;
        RECT 1960.680 1655.390 1961.280 1655.530 ;
        RECT 1961.140 1608.190 1961.280 1655.390 ;
        RECT 1961.080 1607.870 1961.340 1608.190 ;
        RECT 1960.620 1593.930 1960.880 1594.250 ;
        RECT 1960.680 1593.650 1960.820 1593.930 ;
        RECT 1960.680 1593.510 1961.280 1593.650 ;
        RECT 1961.140 1463.090 1961.280 1593.510 ;
        RECT 1960.680 1462.950 1961.280 1463.090 ;
        RECT 1960.680 1449.070 1960.820 1462.950 ;
        RECT 1960.620 1448.750 1960.880 1449.070 ;
        RECT 1961.080 1448.750 1961.340 1449.070 ;
        RECT 1961.140 1393.990 1961.280 1448.750 ;
        RECT 1960.620 1393.670 1960.880 1393.990 ;
        RECT 1961.080 1393.670 1961.340 1393.990 ;
        RECT 1960.680 1352.510 1960.820 1393.670 ;
        RECT 1960.620 1352.190 1960.880 1352.510 ;
        RECT 1961.080 1321.250 1961.340 1321.570 ;
        RECT 1961.140 1249.490 1961.280 1321.250 ;
        RECT 1960.620 1249.170 1960.880 1249.490 ;
        RECT 1961.080 1249.170 1961.340 1249.490 ;
        RECT 1960.680 1249.005 1960.820 1249.170 ;
        RECT 1960.610 1248.635 1960.890 1249.005 ;
        RECT 1961.990 1248.635 1962.270 1249.005 ;
        RECT 1962.060 1200.870 1962.200 1248.635 ;
        RECT 1961.080 1200.550 1961.340 1200.870 ;
        RECT 1962.000 1200.550 1962.260 1200.870 ;
        RECT 1961.140 1183.870 1961.280 1200.550 ;
        RECT 1961.080 1183.550 1961.340 1183.870 ;
        RECT 1961.080 1110.790 1961.340 1111.110 ;
        RECT 1961.140 1087.050 1961.280 1110.790 ;
        RECT 1960.680 1086.910 1961.280 1087.050 ;
        RECT 1960.680 1062.685 1960.820 1086.910 ;
        RECT 1960.610 1062.315 1960.890 1062.685 ;
        RECT 1961.530 1062.315 1961.810 1062.685 ;
        RECT 1961.600 976.470 1961.740 1062.315 ;
        RECT 1960.160 976.150 1960.420 976.470 ;
        RECT 1961.540 976.150 1961.800 976.470 ;
        RECT 1960.220 952.525 1960.360 976.150 ;
        RECT 1960.150 952.155 1960.430 952.525 ;
        RECT 1961.070 952.155 1961.350 952.525 ;
        RECT 1961.140 911.610 1961.280 952.155 ;
        RECT 1960.680 911.470 1961.280 911.610 ;
        RECT 1960.680 910.930 1960.820 911.470 ;
        RECT 1960.680 910.790 1961.280 910.930 ;
        RECT 1961.140 904.050 1961.280 910.790 ;
        RECT 1961.080 903.730 1961.340 904.050 ;
        RECT 1960.620 855.450 1960.880 855.770 ;
        RECT 1960.680 814.290 1960.820 855.450 ;
        RECT 1960.620 813.970 1960.880 814.290 ;
        RECT 1961.540 813.970 1961.800 814.290 ;
        RECT 1961.600 741.870 1961.740 813.970 ;
        RECT 1961.540 741.550 1961.800 741.870 ;
        RECT 1960.620 676.270 1960.880 676.590 ;
        RECT 1960.680 651.850 1960.820 676.270 ;
        RECT 1960.680 651.710 1961.280 651.850 ;
        RECT 1961.140 627.970 1961.280 651.710 ;
        RECT 1961.080 627.650 1961.340 627.970 ;
        RECT 1961.540 627.650 1961.800 627.970 ;
        RECT 1961.600 579.885 1961.740 627.650 ;
        RECT 1960.610 579.515 1960.890 579.885 ;
        RECT 1961.530 579.515 1961.810 579.885 ;
        RECT 1960.620 579.370 1960.880 579.515 ;
        RECT 1961.540 579.370 1961.800 579.515 ;
        RECT 1961.600 483.325 1961.740 579.370 ;
        RECT 1960.610 482.955 1960.890 483.325 ;
        RECT 1961.530 482.955 1961.810 483.325 ;
        RECT 1960.680 434.510 1960.820 482.955 ;
        RECT 1960.620 434.190 1960.880 434.510 ;
        RECT 1960.620 386.250 1960.880 386.570 ;
        RECT 1960.680 338.630 1960.820 386.250 ;
        RECT 1960.620 338.310 1960.880 338.630 ;
        RECT 1961.080 337.970 1961.340 338.290 ;
        RECT 1961.140 308.710 1961.280 337.970 ;
        RECT 1961.080 308.390 1961.340 308.710 ;
        RECT 1962.000 308.390 1962.260 308.710 ;
        RECT 1962.060 283.290 1962.200 308.390 ;
        RECT 1961.600 283.150 1962.200 283.290 ;
        RECT 1961.600 282.870 1961.740 283.150 ;
        RECT 1961.540 282.550 1961.800 282.870 ;
        RECT 1960.620 234.950 1960.880 235.270 ;
        RECT 1960.680 234.590 1960.820 234.950 ;
        RECT 1960.620 234.270 1960.880 234.590 ;
        RECT 1960.620 233.590 1960.880 233.910 ;
        RECT 1960.680 169.050 1960.820 233.590 ;
        RECT 1960.220 168.910 1960.820 169.050 ;
        RECT 1960.220 158.170 1960.360 168.910 ;
        RECT 1960.220 158.030 1961.280 158.170 ;
        RECT 1961.140 144.830 1961.280 158.030 ;
        RECT 1960.160 144.510 1960.420 144.830 ;
        RECT 1961.080 144.510 1961.340 144.830 ;
        RECT 1960.220 96.970 1960.360 144.510 ;
        RECT 1960.220 96.830 1960.820 96.970 ;
        RECT 1960.680 72.490 1960.820 96.830 ;
        RECT 1960.220 72.350 1960.820 72.490 ;
        RECT 1960.220 46.230 1960.360 72.350 ;
        RECT 1635.400 45.910 1635.660 46.230 ;
        RECT 1960.160 45.910 1960.420 46.230 ;
        RECT 1635.460 19.370 1635.600 45.910 ;
        RECT 1584.800 19.050 1585.060 19.370 ;
        RECT 1635.400 19.050 1635.660 19.370 ;
        RECT 1584.860 2.400 1585.000 19.050 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
      LAYER via2 ;
        RECT 1960.610 1248.680 1960.890 1248.960 ;
        RECT 1961.990 1248.680 1962.270 1248.960 ;
        RECT 1960.610 1062.360 1960.890 1062.640 ;
        RECT 1961.530 1062.360 1961.810 1062.640 ;
        RECT 1960.150 952.200 1960.430 952.480 ;
        RECT 1961.070 952.200 1961.350 952.480 ;
        RECT 1960.610 579.560 1960.890 579.840 ;
        RECT 1961.530 579.560 1961.810 579.840 ;
        RECT 1960.610 483.000 1960.890 483.280 ;
        RECT 1961.530 483.000 1961.810 483.280 ;
      LAYER met3 ;
        RECT 1960.585 1248.970 1960.915 1248.985 ;
        RECT 1961.965 1248.970 1962.295 1248.985 ;
        RECT 1960.585 1248.670 1962.295 1248.970 ;
        RECT 1960.585 1248.655 1960.915 1248.670 ;
        RECT 1961.965 1248.655 1962.295 1248.670 ;
        RECT 1960.585 1062.650 1960.915 1062.665 ;
        RECT 1961.505 1062.650 1961.835 1062.665 ;
        RECT 1960.585 1062.350 1961.835 1062.650 ;
        RECT 1960.585 1062.335 1960.915 1062.350 ;
        RECT 1961.505 1062.335 1961.835 1062.350 ;
        RECT 1960.125 952.490 1960.455 952.505 ;
        RECT 1961.045 952.490 1961.375 952.505 ;
        RECT 1960.125 952.190 1961.375 952.490 ;
        RECT 1960.125 952.175 1960.455 952.190 ;
        RECT 1961.045 952.175 1961.375 952.190 ;
        RECT 1960.585 579.850 1960.915 579.865 ;
        RECT 1961.505 579.850 1961.835 579.865 ;
        RECT 1960.585 579.550 1961.835 579.850 ;
        RECT 1960.585 579.535 1960.915 579.550 ;
        RECT 1961.505 579.535 1961.835 579.550 ;
        RECT 1960.585 483.290 1960.915 483.305 ;
        RECT 1961.505 483.290 1961.835 483.305 ;
        RECT 1960.585 482.990 1961.835 483.290 ;
        RECT 1960.585 482.975 1960.915 482.990 ;
        RECT 1961.505 482.975 1961.835 482.990 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1642.730 45.460 1643.050 45.520 ;
        RECT 1973.930 45.460 1974.250 45.520 ;
        RECT 1642.730 45.320 1974.250 45.460 ;
        RECT 1642.730 45.260 1643.050 45.320 ;
        RECT 1973.930 45.260 1974.250 45.320 ;
        RECT 1602.250 15.200 1602.570 15.260 ;
        RECT 1642.730 15.200 1643.050 15.260 ;
        RECT 1602.250 15.060 1643.050 15.200 ;
        RECT 1602.250 15.000 1602.570 15.060 ;
        RECT 1642.730 15.000 1643.050 15.060 ;
      LAYER via ;
        RECT 1642.760 45.260 1643.020 45.520 ;
        RECT 1973.960 45.260 1974.220 45.520 ;
        RECT 1602.280 15.000 1602.540 15.260 ;
        RECT 1642.760 15.000 1643.020 15.260 ;
      LAYER met2 ;
        RECT 1973.420 1700.410 1973.700 1702.400 ;
        RECT 1973.420 1700.270 1974.160 1700.410 ;
        RECT 1973.420 1700.000 1973.700 1700.270 ;
        RECT 1974.020 45.550 1974.160 1700.270 ;
        RECT 1642.760 45.230 1643.020 45.550 ;
        RECT 1973.960 45.230 1974.220 45.550 ;
        RECT 1642.820 15.290 1642.960 45.230 ;
        RECT 1602.280 14.970 1602.540 15.290 ;
        RECT 1642.760 14.970 1643.020 15.290 ;
        RECT 1602.340 2.400 1602.480 14.970 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1732.430 36.280 1732.750 36.340 ;
        RECT 1980.830 36.280 1981.150 36.340 ;
        RECT 1732.430 36.140 1981.150 36.280 ;
        RECT 1732.430 36.080 1732.750 36.140 ;
        RECT 1980.830 36.080 1981.150 36.140 ;
        RECT 1620.190 16.900 1620.510 16.960 ;
        RECT 1732.430 16.900 1732.750 16.960 ;
        RECT 1620.190 16.760 1732.750 16.900 ;
        RECT 1620.190 16.700 1620.510 16.760 ;
        RECT 1732.430 16.700 1732.750 16.760 ;
      LAYER via ;
        RECT 1732.460 36.080 1732.720 36.340 ;
        RECT 1980.860 36.080 1981.120 36.340 ;
        RECT 1620.220 16.700 1620.480 16.960 ;
        RECT 1732.460 16.700 1732.720 16.960 ;
      LAYER met2 ;
        RECT 1982.620 1700.410 1982.900 1702.400 ;
        RECT 1980.920 1700.270 1982.900 1700.410 ;
        RECT 1980.920 36.370 1981.060 1700.270 ;
        RECT 1982.620 1700.000 1982.900 1700.270 ;
        RECT 1732.460 36.050 1732.720 36.370 ;
        RECT 1980.860 36.050 1981.120 36.370 ;
        RECT 1732.520 16.990 1732.660 36.050 ;
        RECT 1620.220 16.670 1620.480 16.990 ;
        RECT 1732.460 16.670 1732.720 16.990 ;
        RECT 1620.280 2.400 1620.420 16.670 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1988.725 1560.685 1988.895 1593.835 ;
        RECT 1988.265 1062.585 1988.435 1076.695 ;
        RECT 1988.265 966.025 1988.435 980.135 ;
        RECT 1988.725 689.605 1988.895 717.655 ;
        RECT 1988.265 386.325 1988.435 434.775 ;
        RECT 1988.265 289.765 1988.435 337.875 ;
        RECT 1675.925 15.725 1676.095 16.575 ;
      LAYER mcon ;
        RECT 1988.725 1593.665 1988.895 1593.835 ;
        RECT 1988.265 1076.525 1988.435 1076.695 ;
        RECT 1988.265 979.965 1988.435 980.135 ;
        RECT 1988.725 717.485 1988.895 717.655 ;
        RECT 1988.265 434.605 1988.435 434.775 ;
        RECT 1988.265 337.705 1988.435 337.875 ;
        RECT 1675.925 16.405 1676.095 16.575 ;
      LAYER met1 ;
        RECT 1988.650 1642.440 1988.970 1642.500 ;
        RECT 1989.570 1642.440 1989.890 1642.500 ;
        RECT 1988.650 1642.300 1989.890 1642.440 ;
        RECT 1988.650 1642.240 1988.970 1642.300 ;
        RECT 1989.570 1642.240 1989.890 1642.300 ;
        RECT 1988.650 1593.820 1988.970 1593.880 ;
        RECT 1988.455 1593.680 1988.970 1593.820 ;
        RECT 1988.650 1593.620 1988.970 1593.680 ;
        RECT 1988.650 1560.840 1988.970 1560.900 ;
        RECT 1988.455 1560.700 1988.970 1560.840 ;
        RECT 1988.650 1560.640 1988.970 1560.700 ;
        RECT 1986.810 1317.400 1987.130 1317.460 ;
        RECT 1988.650 1317.400 1988.970 1317.460 ;
        RECT 1986.810 1317.260 1988.970 1317.400 ;
        RECT 1986.810 1317.200 1987.130 1317.260 ;
        RECT 1988.650 1317.200 1988.970 1317.260 ;
        RECT 1986.810 1303.800 1987.130 1303.860 ;
        RECT 1988.650 1303.800 1988.970 1303.860 ;
        RECT 1986.810 1303.660 1988.970 1303.800 ;
        RECT 1986.810 1303.600 1987.130 1303.660 ;
        RECT 1988.650 1303.600 1988.970 1303.660 ;
        RECT 1988.650 1159.300 1988.970 1159.360 ;
        RECT 1989.570 1159.300 1989.890 1159.360 ;
        RECT 1988.650 1159.160 1989.890 1159.300 ;
        RECT 1988.650 1159.100 1988.970 1159.160 ;
        RECT 1989.570 1159.100 1989.890 1159.160 ;
        RECT 1988.650 1124.760 1988.970 1125.020 ;
        RECT 1988.740 1124.340 1988.880 1124.760 ;
        RECT 1988.650 1124.080 1988.970 1124.340 ;
        RECT 1988.190 1076.680 1988.510 1076.740 ;
        RECT 1987.995 1076.540 1988.510 1076.680 ;
        RECT 1988.190 1076.480 1988.510 1076.540 ;
        RECT 1987.730 1062.740 1988.050 1062.800 ;
        RECT 1988.205 1062.740 1988.495 1062.785 ;
        RECT 1987.730 1062.600 1988.495 1062.740 ;
        RECT 1987.730 1062.540 1988.050 1062.600 ;
        RECT 1988.205 1062.555 1988.495 1062.600 ;
        RECT 1986.810 1014.460 1987.130 1014.520 ;
        RECT 1988.650 1014.460 1988.970 1014.520 ;
        RECT 1986.810 1014.320 1988.970 1014.460 ;
        RECT 1986.810 1014.260 1987.130 1014.320 ;
        RECT 1988.650 1014.260 1988.970 1014.320 ;
        RECT 1988.190 980.120 1988.510 980.180 ;
        RECT 1987.995 979.980 1988.510 980.120 ;
        RECT 1988.190 979.920 1988.510 979.980 ;
        RECT 1987.730 966.180 1988.050 966.240 ;
        RECT 1988.205 966.180 1988.495 966.225 ;
        RECT 1987.730 966.040 1988.495 966.180 ;
        RECT 1987.730 965.980 1988.050 966.040 ;
        RECT 1988.205 965.995 1988.495 966.040 ;
        RECT 1988.650 931.640 1988.970 931.900 ;
        RECT 1988.740 931.220 1988.880 931.640 ;
        RECT 1988.650 930.960 1988.970 931.220 ;
        RECT 1986.810 910.760 1987.130 910.820 ;
        RECT 1988.650 910.760 1988.970 910.820 ;
        RECT 1986.810 910.620 1988.970 910.760 ;
        RECT 1986.810 910.560 1987.130 910.620 ;
        RECT 1988.650 910.560 1988.970 910.620 ;
        RECT 1988.650 717.640 1988.970 717.700 ;
        RECT 1988.455 717.500 1988.970 717.640 ;
        RECT 1988.650 717.440 1988.970 717.500 ;
        RECT 1988.650 689.760 1988.970 689.820 ;
        RECT 1988.455 689.620 1988.970 689.760 ;
        RECT 1988.650 689.560 1988.970 689.620 ;
        RECT 1988.190 545.400 1988.510 545.660 ;
        RECT 1988.280 544.980 1988.420 545.400 ;
        RECT 1988.190 544.720 1988.510 544.980 ;
        RECT 1988.190 434.760 1988.510 434.820 ;
        RECT 1987.995 434.620 1988.510 434.760 ;
        RECT 1988.190 434.560 1988.510 434.620 ;
        RECT 1988.190 386.480 1988.510 386.540 ;
        RECT 1987.995 386.340 1988.510 386.480 ;
        RECT 1988.190 386.280 1988.510 386.340 ;
        RECT 1988.190 337.860 1988.510 337.920 ;
        RECT 1987.995 337.720 1988.510 337.860 ;
        RECT 1988.190 337.660 1988.510 337.720 ;
        RECT 1988.205 289.920 1988.495 289.965 ;
        RECT 1988.650 289.920 1988.970 289.980 ;
        RECT 1988.205 289.780 1988.970 289.920 ;
        RECT 1988.205 289.735 1988.495 289.780 ;
        RECT 1988.650 289.720 1988.970 289.780 ;
        RECT 1988.190 62.460 1988.510 62.520 ;
        RECT 1987.820 62.320 1988.510 62.460 ;
        RECT 1987.820 62.180 1987.960 62.320 ;
        RECT 1988.190 62.260 1988.510 62.320 ;
        RECT 1987.730 61.920 1988.050 62.180 ;
        RECT 1739.790 36.620 1740.110 36.680 ;
        RECT 1987.730 36.620 1988.050 36.680 ;
        RECT 1739.790 36.480 1988.050 36.620 ;
        RECT 1739.790 36.420 1740.110 36.480 ;
        RECT 1987.730 36.420 1988.050 36.480 ;
        RECT 1675.865 16.560 1676.155 16.605 ;
        RECT 1739.790 16.560 1740.110 16.620 ;
        RECT 1675.865 16.420 1740.110 16.560 ;
        RECT 1675.865 16.375 1676.155 16.420 ;
        RECT 1739.790 16.360 1740.110 16.420 ;
        RECT 1638.130 15.880 1638.450 15.940 ;
        RECT 1675.865 15.880 1676.155 15.925 ;
        RECT 1638.130 15.740 1676.155 15.880 ;
        RECT 1638.130 15.680 1638.450 15.740 ;
        RECT 1675.865 15.695 1676.155 15.740 ;
      LAYER via ;
        RECT 1988.680 1642.240 1988.940 1642.500 ;
        RECT 1989.600 1642.240 1989.860 1642.500 ;
        RECT 1988.680 1593.620 1988.940 1593.880 ;
        RECT 1988.680 1560.640 1988.940 1560.900 ;
        RECT 1986.840 1317.200 1987.100 1317.460 ;
        RECT 1988.680 1317.200 1988.940 1317.460 ;
        RECT 1986.840 1303.600 1987.100 1303.860 ;
        RECT 1988.680 1303.600 1988.940 1303.860 ;
        RECT 1988.680 1159.100 1988.940 1159.360 ;
        RECT 1989.600 1159.100 1989.860 1159.360 ;
        RECT 1988.680 1124.760 1988.940 1125.020 ;
        RECT 1988.680 1124.080 1988.940 1124.340 ;
        RECT 1988.220 1076.480 1988.480 1076.740 ;
        RECT 1987.760 1062.540 1988.020 1062.800 ;
        RECT 1986.840 1014.260 1987.100 1014.520 ;
        RECT 1988.680 1014.260 1988.940 1014.520 ;
        RECT 1988.220 979.920 1988.480 980.180 ;
        RECT 1987.760 965.980 1988.020 966.240 ;
        RECT 1988.680 931.640 1988.940 931.900 ;
        RECT 1988.680 930.960 1988.940 931.220 ;
        RECT 1986.840 910.560 1987.100 910.820 ;
        RECT 1988.680 910.560 1988.940 910.820 ;
        RECT 1988.680 717.440 1988.940 717.700 ;
        RECT 1988.680 689.560 1988.940 689.820 ;
        RECT 1988.220 545.400 1988.480 545.660 ;
        RECT 1988.220 544.720 1988.480 544.980 ;
        RECT 1988.220 434.560 1988.480 434.820 ;
        RECT 1988.220 386.280 1988.480 386.540 ;
        RECT 1988.220 337.660 1988.480 337.920 ;
        RECT 1988.680 289.720 1988.940 289.980 ;
        RECT 1988.220 62.260 1988.480 62.520 ;
        RECT 1987.760 61.920 1988.020 62.180 ;
        RECT 1739.820 36.420 1740.080 36.680 ;
        RECT 1987.760 36.420 1988.020 36.680 ;
        RECT 1739.820 16.360 1740.080 16.620 ;
        RECT 1638.160 15.680 1638.420 15.940 ;
      LAYER met2 ;
        RECT 1991.820 1700.410 1992.100 1702.400 ;
        RECT 1989.660 1700.270 1992.100 1700.410 ;
        RECT 1989.660 1642.530 1989.800 1700.270 ;
        RECT 1991.820 1700.000 1992.100 1700.270 ;
        RECT 1988.680 1642.210 1988.940 1642.530 ;
        RECT 1989.600 1642.210 1989.860 1642.530 ;
        RECT 1988.740 1593.910 1988.880 1642.210 ;
        RECT 1988.680 1593.590 1988.940 1593.910 ;
        RECT 1988.680 1560.610 1988.940 1560.930 ;
        RECT 1988.740 1463.090 1988.880 1560.610 ;
        RECT 1988.280 1462.950 1988.880 1463.090 ;
        RECT 1988.280 1414.130 1988.420 1462.950 ;
        RECT 1988.280 1413.990 1988.880 1414.130 ;
        RECT 1988.740 1400.645 1988.880 1413.990 ;
        RECT 1988.670 1400.275 1988.950 1400.645 ;
        RECT 1986.830 1399.595 1987.110 1399.965 ;
        RECT 1986.900 1317.490 1987.040 1399.595 ;
        RECT 1986.840 1317.170 1987.100 1317.490 ;
        RECT 1988.680 1317.170 1988.940 1317.490 ;
        RECT 1988.740 1303.890 1988.880 1317.170 ;
        RECT 1986.840 1303.570 1987.100 1303.890 ;
        RECT 1988.680 1303.570 1988.940 1303.890 ;
        RECT 1986.900 1297.285 1987.040 1303.570 ;
        RECT 1986.830 1296.915 1987.110 1297.285 ;
        RECT 1989.590 1296.915 1989.870 1297.285 ;
        RECT 1989.660 1159.390 1989.800 1296.915 ;
        RECT 1988.680 1159.070 1988.940 1159.390 ;
        RECT 1989.600 1159.070 1989.860 1159.390 ;
        RECT 1988.740 1125.050 1988.880 1159.070 ;
        RECT 1988.680 1124.730 1988.940 1125.050 ;
        RECT 1988.680 1124.050 1988.940 1124.370 ;
        RECT 1988.740 1110.850 1988.880 1124.050 ;
        RECT 1988.280 1110.710 1988.880 1110.850 ;
        RECT 1988.280 1076.770 1988.420 1110.710 ;
        RECT 1988.220 1076.450 1988.480 1076.770 ;
        RECT 1987.760 1062.685 1988.020 1062.830 ;
        RECT 1986.830 1062.315 1987.110 1062.685 ;
        RECT 1987.750 1062.315 1988.030 1062.685 ;
        RECT 1986.900 1014.550 1987.040 1062.315 ;
        RECT 1988.740 1014.550 1988.880 1014.705 ;
        RECT 1986.840 1014.230 1987.100 1014.550 ;
        RECT 1988.680 1014.290 1988.940 1014.550 ;
        RECT 1988.280 1014.230 1988.940 1014.290 ;
        RECT 1988.280 1014.150 1988.880 1014.230 ;
        RECT 1988.280 980.210 1988.420 1014.150 ;
        RECT 1988.220 979.890 1988.480 980.210 ;
        RECT 1987.760 966.125 1988.020 966.270 ;
        RECT 1987.750 965.755 1988.030 966.125 ;
        RECT 1988.670 965.755 1988.950 966.125 ;
        RECT 1988.740 931.930 1988.880 965.755 ;
        RECT 1988.680 931.610 1988.940 931.930 ;
        RECT 1988.680 930.930 1988.940 931.250 ;
        RECT 1988.740 910.850 1988.880 930.930 ;
        RECT 1986.840 910.530 1987.100 910.850 ;
        RECT 1988.680 910.530 1988.940 910.850 ;
        RECT 1986.900 862.765 1987.040 910.530 ;
        RECT 1986.830 862.395 1987.110 862.765 ;
        RECT 1987.750 862.395 1988.030 862.765 ;
        RECT 1987.820 844.970 1987.960 862.395 ;
        RECT 1987.820 844.830 1988.420 844.970 ;
        RECT 1988.280 821.170 1988.420 844.830 ;
        RECT 1988.280 821.030 1988.880 821.170 ;
        RECT 1988.740 717.730 1988.880 821.030 ;
        RECT 1988.680 717.410 1988.940 717.730 ;
        RECT 1988.680 689.530 1988.940 689.850 ;
        RECT 1988.740 594.050 1988.880 689.530 ;
        RECT 1988.280 593.910 1988.880 594.050 ;
        RECT 1988.280 545.690 1988.420 593.910 ;
        RECT 1988.220 545.370 1988.480 545.690 ;
        RECT 1988.220 544.690 1988.480 545.010 ;
        RECT 1988.280 434.850 1988.420 544.690 ;
        RECT 1988.220 434.530 1988.480 434.850 ;
        RECT 1988.220 386.250 1988.480 386.570 ;
        RECT 1988.280 337.950 1988.420 386.250 ;
        RECT 1988.220 337.630 1988.480 337.950 ;
        RECT 1988.680 289.690 1988.940 290.010 ;
        RECT 1988.740 207.130 1988.880 289.690 ;
        RECT 1988.280 206.990 1988.880 207.130 ;
        RECT 1988.280 206.450 1988.420 206.990 ;
        RECT 1988.280 206.310 1988.880 206.450 ;
        RECT 1988.740 110.570 1988.880 206.310 ;
        RECT 1988.280 110.430 1988.880 110.570 ;
        RECT 1988.280 62.550 1988.420 110.430 ;
        RECT 1988.220 62.230 1988.480 62.550 ;
        RECT 1987.760 61.890 1988.020 62.210 ;
        RECT 1987.820 36.710 1987.960 61.890 ;
        RECT 1739.820 36.390 1740.080 36.710 ;
        RECT 1987.760 36.390 1988.020 36.710 ;
        RECT 1739.880 16.650 1740.020 36.390 ;
        RECT 1739.820 16.330 1740.080 16.650 ;
        RECT 1638.160 15.650 1638.420 15.970 ;
        RECT 1638.220 2.400 1638.360 15.650 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
      LAYER via2 ;
        RECT 1988.670 1400.320 1988.950 1400.600 ;
        RECT 1986.830 1399.640 1987.110 1399.920 ;
        RECT 1986.830 1296.960 1987.110 1297.240 ;
        RECT 1989.590 1296.960 1989.870 1297.240 ;
        RECT 1986.830 1062.360 1987.110 1062.640 ;
        RECT 1987.750 1062.360 1988.030 1062.640 ;
        RECT 1987.750 965.800 1988.030 966.080 ;
        RECT 1988.670 965.800 1988.950 966.080 ;
        RECT 1986.830 862.440 1987.110 862.720 ;
        RECT 1987.750 862.440 1988.030 862.720 ;
      LAYER met3 ;
        RECT 1988.645 1400.610 1988.975 1400.625 ;
        RECT 1988.645 1400.310 1989.650 1400.610 ;
        RECT 1988.645 1400.295 1988.975 1400.310 ;
        RECT 1986.805 1399.930 1987.135 1399.945 ;
        RECT 1989.350 1399.930 1989.650 1400.310 ;
        RECT 1986.805 1399.630 1989.650 1399.930 ;
        RECT 1986.805 1399.615 1987.135 1399.630 ;
        RECT 1986.805 1297.250 1987.135 1297.265 ;
        RECT 1989.565 1297.250 1989.895 1297.265 ;
        RECT 1986.805 1296.950 1989.895 1297.250 ;
        RECT 1986.805 1296.935 1987.135 1296.950 ;
        RECT 1989.565 1296.935 1989.895 1296.950 ;
        RECT 1986.805 1062.650 1987.135 1062.665 ;
        RECT 1987.725 1062.650 1988.055 1062.665 ;
        RECT 1986.805 1062.350 1988.055 1062.650 ;
        RECT 1986.805 1062.335 1987.135 1062.350 ;
        RECT 1987.725 1062.335 1988.055 1062.350 ;
        RECT 1987.725 966.090 1988.055 966.105 ;
        RECT 1988.645 966.090 1988.975 966.105 ;
        RECT 1987.725 965.790 1988.975 966.090 ;
        RECT 1987.725 965.775 1988.055 965.790 ;
        RECT 1988.645 965.775 1988.975 965.790 ;
        RECT 1986.805 862.730 1987.135 862.745 ;
        RECT 1987.725 862.730 1988.055 862.745 ;
        RECT 1986.805 862.430 1988.055 862.730 ;
        RECT 1986.805 862.415 1987.135 862.430 ;
        RECT 1987.725 862.415 1988.055 862.430 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 1690.380 1662.830 1690.440 ;
        RECT 2001.070 1690.380 2001.390 1690.440 ;
        RECT 1662.510 1690.240 2001.390 1690.380 ;
        RECT 1662.510 1690.180 1662.830 1690.240 ;
        RECT 2001.070 1690.180 2001.390 1690.240 ;
        RECT 1656.070 20.640 1656.390 20.700 ;
        RECT 1662.510 20.640 1662.830 20.700 ;
        RECT 1656.070 20.500 1662.830 20.640 ;
        RECT 1656.070 20.440 1656.390 20.500 ;
        RECT 1662.510 20.440 1662.830 20.500 ;
      LAYER via ;
        RECT 1662.540 1690.180 1662.800 1690.440 ;
        RECT 2001.100 1690.180 2001.360 1690.440 ;
        RECT 1656.100 20.440 1656.360 20.700 ;
        RECT 1662.540 20.440 1662.800 20.700 ;
      LAYER met2 ;
        RECT 2001.020 1700.000 2001.300 1702.400 ;
        RECT 2001.160 1690.470 2001.300 1700.000 ;
        RECT 1662.540 1690.150 1662.800 1690.470 ;
        RECT 2001.100 1690.150 2001.360 1690.470 ;
        RECT 1662.600 20.730 1662.740 1690.150 ;
        RECT 1656.100 20.410 1656.360 20.730 ;
        RECT 1662.540 20.410 1662.800 20.730 ;
        RECT 1656.160 2.400 1656.300 20.410 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1673.550 44.780 1673.870 44.840 ;
        RECT 2008.430 44.780 2008.750 44.840 ;
        RECT 1673.550 44.640 2008.750 44.780 ;
        RECT 1673.550 44.580 1673.870 44.640 ;
        RECT 2008.430 44.580 2008.750 44.640 ;
      LAYER via ;
        RECT 1673.580 44.580 1673.840 44.840 ;
        RECT 2008.460 44.580 2008.720 44.840 ;
      LAYER met2 ;
        RECT 2010.220 1700.410 2010.500 1702.400 ;
        RECT 2008.520 1700.270 2010.500 1700.410 ;
        RECT 2008.520 44.870 2008.660 1700.270 ;
        RECT 2010.220 1700.000 2010.500 1700.270 ;
        RECT 1673.580 44.550 1673.840 44.870 ;
        RECT 2008.460 44.550 2008.720 44.870 ;
        RECT 1673.640 2.400 1673.780 44.550 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1779.885 1685.465 1780.055 1686.655 ;
        RECT 1925.245 1686.485 1925.415 1690.735 ;
        RECT 1977.225 1689.545 1977.395 1690.735 ;
        RECT 1993.785 1686.485 1993.955 1689.715 ;
      LAYER mcon ;
        RECT 1925.245 1690.565 1925.415 1690.735 ;
        RECT 1977.225 1690.565 1977.395 1690.735 ;
        RECT 1993.785 1689.545 1993.955 1689.715 ;
        RECT 1779.885 1686.485 1780.055 1686.655 ;
      LAYER met1 ;
        RECT 1925.185 1690.720 1925.475 1690.765 ;
        RECT 1977.165 1690.720 1977.455 1690.765 ;
        RECT 1925.185 1690.580 1977.455 1690.720 ;
        RECT 1925.185 1690.535 1925.475 1690.580 ;
        RECT 1977.165 1690.535 1977.455 1690.580 ;
        RECT 1977.165 1689.700 1977.455 1689.745 ;
        RECT 1993.725 1689.700 1994.015 1689.745 ;
        RECT 1977.165 1689.560 1994.015 1689.700 ;
        RECT 1977.165 1689.515 1977.455 1689.560 ;
        RECT 1993.725 1689.515 1994.015 1689.560 ;
        RECT 1779.825 1686.640 1780.115 1686.685 ;
        RECT 1828.570 1686.640 1828.890 1686.700 ;
        RECT 1779.825 1686.500 1828.890 1686.640 ;
        RECT 1779.825 1686.455 1780.115 1686.500 ;
        RECT 1828.570 1686.440 1828.890 1686.500 ;
        RECT 1892.510 1686.640 1892.830 1686.700 ;
        RECT 1925.185 1686.640 1925.475 1686.685 ;
        RECT 1892.510 1686.500 1925.475 1686.640 ;
        RECT 1892.510 1686.440 1892.830 1686.500 ;
        RECT 1925.185 1686.455 1925.475 1686.500 ;
        RECT 1993.725 1686.640 1994.015 1686.685 ;
        RECT 2019.470 1686.640 2019.790 1686.700 ;
        RECT 1993.725 1686.500 2019.790 1686.640 ;
        RECT 1993.725 1686.455 1994.015 1686.500 ;
        RECT 2019.470 1686.440 2019.790 1686.500 ;
        RECT 1697.010 1686.300 1697.330 1686.360 ;
        RECT 1697.010 1686.160 1728.520 1686.300 ;
        RECT 1697.010 1686.100 1697.330 1686.160 ;
        RECT 1728.380 1685.960 1728.520 1686.160 ;
        RECT 1728.380 1685.820 1739.560 1685.960 ;
        RECT 1739.420 1685.620 1739.560 1685.820 ;
        RECT 1779.825 1685.620 1780.115 1685.665 ;
        RECT 1739.420 1685.480 1780.115 1685.620 ;
        RECT 1779.825 1685.435 1780.115 1685.480 ;
        RECT 1691.490 15.200 1691.810 15.260 ;
        RECT 1697.010 15.200 1697.330 15.260 ;
        RECT 1691.490 15.060 1697.330 15.200 ;
        RECT 1691.490 15.000 1691.810 15.060 ;
        RECT 1697.010 15.000 1697.330 15.060 ;
      LAYER via ;
        RECT 1828.600 1686.440 1828.860 1686.700 ;
        RECT 1892.540 1686.440 1892.800 1686.700 ;
        RECT 2019.500 1686.440 2019.760 1686.700 ;
        RECT 1697.040 1686.100 1697.300 1686.360 ;
        RECT 1691.520 15.000 1691.780 15.260 ;
        RECT 1697.040 15.000 1697.300 15.260 ;
      LAYER met2 ;
        RECT 2019.420 1700.000 2019.700 1702.400 ;
        RECT 1829.050 1687.235 1829.330 1687.605 ;
        RECT 1892.530 1687.235 1892.810 1687.605 ;
        RECT 1828.600 1686.410 1828.860 1686.730 ;
        RECT 1697.040 1686.070 1697.300 1686.390 ;
        RECT 1828.660 1686.130 1828.800 1686.410 ;
        RECT 1829.120 1686.130 1829.260 1687.235 ;
        RECT 1892.600 1686.730 1892.740 1687.235 ;
        RECT 2019.560 1686.730 2019.700 1700.000 ;
        RECT 1892.540 1686.410 1892.800 1686.730 ;
        RECT 2019.500 1686.410 2019.760 1686.730 ;
        RECT 1697.100 15.290 1697.240 1686.070 ;
        RECT 1828.660 1685.990 1829.260 1686.130 ;
        RECT 1691.520 14.970 1691.780 15.290 ;
        RECT 1697.040 14.970 1697.300 15.290 ;
        RECT 1691.580 2.400 1691.720 14.970 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
      LAYER via2 ;
        RECT 1829.050 1687.280 1829.330 1687.560 ;
        RECT 1892.530 1687.280 1892.810 1687.560 ;
      LAYER met3 ;
        RECT 1829.025 1687.570 1829.355 1687.585 ;
        RECT 1892.505 1687.570 1892.835 1687.585 ;
        RECT 1829.025 1687.270 1892.835 1687.570 ;
        RECT 1829.025 1687.255 1829.355 1687.270 ;
        RECT 1892.505 1687.255 1892.835 1687.270 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1518.070 1678.140 1518.390 1678.200 ;
        RECT 1521.750 1678.140 1522.070 1678.200 ;
        RECT 1518.070 1678.000 1522.070 1678.140 ;
        RECT 1518.070 1677.940 1518.390 1678.000 ;
        RECT 1521.750 1677.940 1522.070 1678.000 ;
        RECT 731.010 66.540 731.330 66.600 ;
        RECT 1518.070 66.540 1518.390 66.600 ;
        RECT 731.010 66.400 1518.390 66.540 ;
        RECT 731.010 66.340 731.330 66.400 ;
        RECT 1518.070 66.340 1518.390 66.400 ;
      LAYER via ;
        RECT 1518.100 1677.940 1518.360 1678.200 ;
        RECT 1521.780 1677.940 1522.040 1678.200 ;
        RECT 731.040 66.340 731.300 66.600 ;
        RECT 1518.100 66.340 1518.360 66.600 ;
      LAYER met2 ;
        RECT 1523.080 1700.410 1523.360 1702.400 ;
        RECT 1521.840 1700.270 1523.360 1700.410 ;
        RECT 1521.840 1678.230 1521.980 1700.270 ;
        RECT 1523.080 1700.000 1523.360 1700.270 ;
        RECT 1518.100 1677.910 1518.360 1678.230 ;
        RECT 1521.780 1677.910 1522.040 1678.230 ;
        RECT 1518.160 66.630 1518.300 1677.910 ;
        RECT 731.040 66.310 731.300 66.630 ;
        RECT 1518.100 66.310 1518.360 66.630 ;
        RECT 731.100 16.730 731.240 66.310 ;
        RECT 728.340 16.590 731.240 16.730 ;
        RECT 728.340 2.400 728.480 16.590 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1759.110 37.980 1759.430 38.040 ;
        RECT 2029.130 37.980 2029.450 38.040 ;
        RECT 1759.110 37.840 2029.450 37.980 ;
        RECT 1759.110 37.780 1759.430 37.840 ;
        RECT 2029.130 37.780 2029.450 37.840 ;
        RECT 1709.430 14.860 1709.750 14.920 ;
        RECT 1759.110 14.860 1759.430 14.920 ;
        RECT 1709.430 14.720 1759.430 14.860 ;
        RECT 1709.430 14.660 1709.750 14.720 ;
        RECT 1759.110 14.660 1759.430 14.720 ;
      LAYER via ;
        RECT 1759.140 37.780 1759.400 38.040 ;
        RECT 2029.160 37.780 2029.420 38.040 ;
        RECT 1709.460 14.660 1709.720 14.920 ;
        RECT 1759.140 14.660 1759.400 14.920 ;
      LAYER met2 ;
        RECT 2028.620 1700.410 2028.900 1702.400 ;
        RECT 2028.620 1700.270 2029.360 1700.410 ;
        RECT 2028.620 1700.000 2028.900 1700.270 ;
        RECT 2029.220 38.070 2029.360 1700.270 ;
        RECT 1759.140 37.750 1759.400 38.070 ;
        RECT 2029.160 37.750 2029.420 38.070 ;
        RECT 1759.200 14.950 1759.340 37.750 ;
        RECT 1709.460 14.630 1709.720 14.950 ;
        RECT 1759.140 14.630 1759.400 14.950 ;
        RECT 1709.520 2.400 1709.660 14.630 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1731.510 1686.300 1731.830 1686.360 ;
        RECT 2037.410 1686.300 2037.730 1686.360 ;
        RECT 1731.510 1686.160 2037.730 1686.300 ;
        RECT 1731.510 1686.100 1731.830 1686.160 ;
        RECT 2037.410 1686.100 2037.730 1686.160 ;
        RECT 1727.370 3.640 1727.690 3.700 ;
        RECT 1731.510 3.640 1731.830 3.700 ;
        RECT 1727.370 3.500 1731.830 3.640 ;
        RECT 1727.370 3.440 1727.690 3.500 ;
        RECT 1731.510 3.440 1731.830 3.500 ;
      LAYER via ;
        RECT 1731.540 1686.100 1731.800 1686.360 ;
        RECT 2037.440 1686.100 2037.700 1686.360 ;
        RECT 1727.400 3.440 1727.660 3.700 ;
        RECT 1731.540 3.440 1731.800 3.700 ;
      LAYER met2 ;
        RECT 2037.360 1700.000 2037.640 1702.400 ;
        RECT 2037.500 1686.390 2037.640 1700.000 ;
        RECT 1731.540 1686.070 1731.800 1686.390 ;
        RECT 2037.440 1686.070 2037.700 1686.390 ;
        RECT 1731.600 3.730 1731.740 1686.070 ;
        RECT 1727.400 3.410 1727.660 3.730 ;
        RECT 1731.540 3.410 1731.800 3.730 ;
        RECT 1727.460 2.400 1727.600 3.410 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2043.925 1490.645 2044.095 1511.215 ;
        RECT 2043.925 1413.805 2044.095 1465.315 ;
        RECT 2043.925 1317.245 2044.095 1393.575 ;
        RECT 2043.465 1110.865 2043.635 1158.975 ;
        RECT 2043.465 1014.305 2043.635 1062.415 ;
        RECT 2043.465 737.885 2043.635 772.735 ;
        RECT 2043.465 641.325 2043.635 676.175 ;
        RECT 2043.465 476.085 2043.635 524.195 ;
        RECT 2043.925 386.325 2044.095 410.635 ;
        RECT 2043.925 338.045 2044.095 352.155 ;
        RECT 2043.925 289.765 2044.095 314.075 ;
        RECT 2043.925 241.825 2044.095 255.935 ;
        RECT 2043.925 192.525 2044.095 234.515 ;
      LAYER mcon ;
        RECT 2043.925 1511.045 2044.095 1511.215 ;
        RECT 2043.925 1465.145 2044.095 1465.315 ;
        RECT 2043.925 1393.405 2044.095 1393.575 ;
        RECT 2043.465 1158.805 2043.635 1158.975 ;
        RECT 2043.465 1062.245 2043.635 1062.415 ;
        RECT 2043.465 772.565 2043.635 772.735 ;
        RECT 2043.465 676.005 2043.635 676.175 ;
        RECT 2043.465 524.025 2043.635 524.195 ;
        RECT 2043.925 410.465 2044.095 410.635 ;
        RECT 2043.925 351.985 2044.095 352.155 ;
        RECT 2043.925 313.905 2044.095 314.075 ;
        RECT 2043.925 255.765 2044.095 255.935 ;
        RECT 2043.925 234.345 2044.095 234.515 ;
      LAYER met1 ;
        RECT 2043.390 1607.900 2043.710 1608.160 ;
        RECT 2043.480 1607.420 2043.620 1607.900 ;
        RECT 2043.850 1607.420 2044.170 1607.480 ;
        RECT 2043.480 1607.280 2044.170 1607.420 ;
        RECT 2043.850 1607.220 2044.170 1607.280 ;
        RECT 2043.850 1511.200 2044.170 1511.260 ;
        RECT 2043.655 1511.060 2044.170 1511.200 ;
        RECT 2043.850 1511.000 2044.170 1511.060 ;
        RECT 2043.850 1490.800 2044.170 1490.860 ;
        RECT 2043.655 1490.660 2044.170 1490.800 ;
        RECT 2043.850 1490.600 2044.170 1490.660 ;
        RECT 2043.850 1465.300 2044.170 1465.360 ;
        RECT 2043.655 1465.160 2044.170 1465.300 ;
        RECT 2043.850 1465.100 2044.170 1465.160 ;
        RECT 2043.850 1413.960 2044.170 1414.020 ;
        RECT 2043.655 1413.820 2044.170 1413.960 ;
        RECT 2043.850 1413.760 2044.170 1413.820 ;
        RECT 2043.850 1393.560 2044.170 1393.620 ;
        RECT 2043.655 1393.420 2044.170 1393.560 ;
        RECT 2043.850 1393.360 2044.170 1393.420 ;
        RECT 2043.850 1317.400 2044.170 1317.460 ;
        RECT 2043.655 1317.260 2044.170 1317.400 ;
        RECT 2043.850 1317.200 2044.170 1317.260 ;
        RECT 2043.850 1220.840 2044.170 1220.900 ;
        RECT 2044.770 1220.840 2045.090 1220.900 ;
        RECT 2043.850 1220.700 2045.090 1220.840 ;
        RECT 2043.850 1220.640 2044.170 1220.700 ;
        RECT 2044.770 1220.640 2045.090 1220.700 ;
        RECT 2043.850 1173.580 2044.170 1173.640 ;
        RECT 2043.480 1173.440 2044.170 1173.580 ;
        RECT 2043.480 1172.960 2043.620 1173.440 ;
        RECT 2043.850 1173.380 2044.170 1173.440 ;
        RECT 2043.390 1172.700 2043.710 1172.960 ;
        RECT 2043.390 1158.960 2043.710 1159.020 ;
        RECT 2043.195 1158.820 2043.710 1158.960 ;
        RECT 2043.390 1158.760 2043.710 1158.820 ;
        RECT 2043.405 1111.020 2043.695 1111.065 ;
        RECT 2043.850 1111.020 2044.170 1111.080 ;
        RECT 2043.405 1110.880 2044.170 1111.020 ;
        RECT 2043.405 1110.835 2043.695 1110.880 ;
        RECT 2043.850 1110.820 2044.170 1110.880 ;
        RECT 2043.850 1077.020 2044.170 1077.080 ;
        RECT 2043.480 1076.880 2044.170 1077.020 ;
        RECT 2043.480 1076.400 2043.620 1076.880 ;
        RECT 2043.850 1076.820 2044.170 1076.880 ;
        RECT 2043.390 1076.140 2043.710 1076.400 ;
        RECT 2043.390 1062.400 2043.710 1062.460 ;
        RECT 2043.195 1062.260 2043.710 1062.400 ;
        RECT 2043.390 1062.200 2043.710 1062.260 ;
        RECT 2043.405 1014.460 2043.695 1014.505 ;
        RECT 2043.850 1014.460 2044.170 1014.520 ;
        RECT 2043.405 1014.320 2044.170 1014.460 ;
        RECT 2043.405 1014.275 2043.695 1014.320 ;
        RECT 2043.850 1014.260 2044.170 1014.320 ;
        RECT 2043.850 980.460 2044.170 980.520 ;
        RECT 2043.480 980.320 2044.170 980.460 ;
        RECT 2043.480 979.840 2043.620 980.320 ;
        RECT 2043.850 980.260 2044.170 980.320 ;
        RECT 2043.390 979.580 2043.710 979.840 ;
        RECT 2043.850 917.900 2044.170 917.960 ;
        RECT 2044.770 917.900 2045.090 917.960 ;
        RECT 2043.850 917.760 2045.090 917.900 ;
        RECT 2043.850 917.700 2044.170 917.760 ;
        RECT 2044.770 917.700 2045.090 917.760 ;
        RECT 2043.850 883.700 2044.170 883.960 ;
        RECT 2043.940 882.940 2044.080 883.700 ;
        RECT 2043.850 882.680 2044.170 882.940 ;
        RECT 2042.930 786.800 2043.250 787.060 ;
        RECT 2043.020 786.320 2043.160 786.800 ;
        RECT 2043.390 786.320 2043.710 786.380 ;
        RECT 2043.020 786.180 2043.710 786.320 ;
        RECT 2043.390 786.120 2043.710 786.180 ;
        RECT 2043.390 772.720 2043.710 772.780 ;
        RECT 2043.195 772.580 2043.710 772.720 ;
        RECT 2043.390 772.520 2043.710 772.580 ;
        RECT 2043.390 738.040 2043.710 738.100 ;
        RECT 2043.195 737.900 2043.710 738.040 ;
        RECT 2043.390 737.840 2043.710 737.900 ;
        RECT 2043.850 690.440 2044.170 690.500 ;
        RECT 2043.480 690.300 2044.170 690.440 ;
        RECT 2043.480 689.820 2043.620 690.300 ;
        RECT 2043.850 690.240 2044.170 690.300 ;
        RECT 2043.390 689.560 2043.710 689.820 ;
        RECT 2043.390 676.160 2043.710 676.220 ;
        RECT 2043.195 676.020 2043.710 676.160 ;
        RECT 2043.390 675.960 2043.710 676.020 ;
        RECT 2043.390 641.480 2043.710 641.540 ;
        RECT 2043.195 641.340 2043.710 641.480 ;
        RECT 2043.390 641.280 2043.710 641.340 ;
        RECT 2043.850 593.880 2044.170 593.940 ;
        RECT 2043.480 593.740 2044.170 593.880 ;
        RECT 2043.480 593.260 2043.620 593.740 ;
        RECT 2043.850 593.680 2044.170 593.740 ;
        RECT 2043.390 593.000 2043.710 593.260 ;
        RECT 2043.390 545.060 2043.710 545.320 ;
        RECT 2043.480 544.920 2043.620 545.060 ;
        RECT 2043.850 544.920 2044.170 544.980 ;
        RECT 2043.480 544.780 2044.170 544.920 ;
        RECT 2043.850 544.720 2044.170 544.780 ;
        RECT 2043.405 524.180 2043.695 524.225 ;
        RECT 2043.850 524.180 2044.170 524.240 ;
        RECT 2043.405 524.040 2044.170 524.180 ;
        RECT 2043.405 523.995 2043.695 524.040 ;
        RECT 2043.850 523.980 2044.170 524.040 ;
        RECT 2043.390 476.240 2043.710 476.300 ;
        RECT 2043.195 476.100 2043.710 476.240 ;
        RECT 2043.390 476.040 2043.710 476.100 ;
        RECT 2043.390 448.500 2043.710 448.760 ;
        RECT 2043.480 448.020 2043.620 448.500 ;
        RECT 2043.850 448.020 2044.170 448.080 ;
        RECT 2043.480 447.880 2044.170 448.020 ;
        RECT 2043.850 447.820 2044.170 447.880 ;
        RECT 2043.850 410.620 2044.170 410.680 ;
        RECT 2043.655 410.480 2044.170 410.620 ;
        RECT 2043.850 410.420 2044.170 410.480 ;
        RECT 2043.850 386.480 2044.170 386.540 ;
        RECT 2043.655 386.340 2044.170 386.480 ;
        RECT 2043.850 386.280 2044.170 386.340 ;
        RECT 2043.850 352.140 2044.170 352.200 ;
        RECT 2043.655 352.000 2044.170 352.140 ;
        RECT 2043.850 351.940 2044.170 352.000 ;
        RECT 2043.850 338.200 2044.170 338.260 ;
        RECT 2043.655 338.060 2044.170 338.200 ;
        RECT 2043.850 338.000 2044.170 338.060 ;
        RECT 2043.850 314.060 2044.170 314.120 ;
        RECT 2043.655 313.920 2044.170 314.060 ;
        RECT 2043.850 313.860 2044.170 313.920 ;
        RECT 2043.850 289.920 2044.170 289.980 ;
        RECT 2043.655 289.780 2044.170 289.920 ;
        RECT 2043.850 289.720 2044.170 289.780 ;
        RECT 2043.850 255.920 2044.170 255.980 ;
        RECT 2043.655 255.780 2044.170 255.920 ;
        RECT 2043.850 255.720 2044.170 255.780 ;
        RECT 2043.390 241.980 2043.710 242.040 ;
        RECT 2043.865 241.980 2044.155 242.025 ;
        RECT 2043.390 241.840 2044.155 241.980 ;
        RECT 2043.390 241.780 2043.710 241.840 ;
        RECT 2043.865 241.795 2044.155 241.840 ;
        RECT 2043.850 234.500 2044.170 234.560 ;
        RECT 2043.655 234.360 2044.170 234.500 ;
        RECT 2043.850 234.300 2044.170 234.360 ;
        RECT 2043.865 192.680 2044.155 192.725 ;
        RECT 2044.310 192.680 2044.630 192.740 ;
        RECT 2043.865 192.540 2044.630 192.680 ;
        RECT 2043.865 192.495 2044.155 192.540 ;
        RECT 2044.310 192.480 2044.630 192.540 ;
        RECT 2043.850 110.740 2044.170 110.800 ;
        RECT 2043.480 110.600 2044.170 110.740 ;
        RECT 2043.480 110.460 2043.620 110.600 ;
        RECT 2043.850 110.540 2044.170 110.600 ;
        RECT 2043.390 110.200 2043.710 110.460 ;
        RECT 1745.310 34.240 1745.630 34.300 ;
        RECT 2043.850 34.240 2044.170 34.300 ;
        RECT 1745.310 34.100 2044.170 34.240 ;
        RECT 1745.310 34.040 1745.630 34.100 ;
        RECT 2043.850 34.040 2044.170 34.100 ;
      LAYER via ;
        RECT 2043.420 1607.900 2043.680 1608.160 ;
        RECT 2043.880 1607.220 2044.140 1607.480 ;
        RECT 2043.880 1511.000 2044.140 1511.260 ;
        RECT 2043.880 1490.600 2044.140 1490.860 ;
        RECT 2043.880 1465.100 2044.140 1465.360 ;
        RECT 2043.880 1413.760 2044.140 1414.020 ;
        RECT 2043.880 1393.360 2044.140 1393.620 ;
        RECT 2043.880 1317.200 2044.140 1317.460 ;
        RECT 2043.880 1220.640 2044.140 1220.900 ;
        RECT 2044.800 1220.640 2045.060 1220.900 ;
        RECT 2043.880 1173.380 2044.140 1173.640 ;
        RECT 2043.420 1172.700 2043.680 1172.960 ;
        RECT 2043.420 1158.760 2043.680 1159.020 ;
        RECT 2043.880 1110.820 2044.140 1111.080 ;
        RECT 2043.880 1076.820 2044.140 1077.080 ;
        RECT 2043.420 1076.140 2043.680 1076.400 ;
        RECT 2043.420 1062.200 2043.680 1062.460 ;
        RECT 2043.880 1014.260 2044.140 1014.520 ;
        RECT 2043.880 980.260 2044.140 980.520 ;
        RECT 2043.420 979.580 2043.680 979.840 ;
        RECT 2043.880 917.700 2044.140 917.960 ;
        RECT 2044.800 917.700 2045.060 917.960 ;
        RECT 2043.880 883.700 2044.140 883.960 ;
        RECT 2043.880 882.680 2044.140 882.940 ;
        RECT 2042.960 786.800 2043.220 787.060 ;
        RECT 2043.420 786.120 2043.680 786.380 ;
        RECT 2043.420 772.520 2043.680 772.780 ;
        RECT 2043.420 737.840 2043.680 738.100 ;
        RECT 2043.880 690.240 2044.140 690.500 ;
        RECT 2043.420 689.560 2043.680 689.820 ;
        RECT 2043.420 675.960 2043.680 676.220 ;
        RECT 2043.420 641.280 2043.680 641.540 ;
        RECT 2043.880 593.680 2044.140 593.940 ;
        RECT 2043.420 593.000 2043.680 593.260 ;
        RECT 2043.420 545.060 2043.680 545.320 ;
        RECT 2043.880 544.720 2044.140 544.980 ;
        RECT 2043.880 523.980 2044.140 524.240 ;
        RECT 2043.420 476.040 2043.680 476.300 ;
        RECT 2043.420 448.500 2043.680 448.760 ;
        RECT 2043.880 447.820 2044.140 448.080 ;
        RECT 2043.880 410.420 2044.140 410.680 ;
        RECT 2043.880 386.280 2044.140 386.540 ;
        RECT 2043.880 351.940 2044.140 352.200 ;
        RECT 2043.880 338.000 2044.140 338.260 ;
        RECT 2043.880 313.860 2044.140 314.120 ;
        RECT 2043.880 289.720 2044.140 289.980 ;
        RECT 2043.880 255.720 2044.140 255.980 ;
        RECT 2043.420 241.780 2043.680 242.040 ;
        RECT 2043.880 234.300 2044.140 234.560 ;
        RECT 2044.340 192.480 2044.600 192.740 ;
        RECT 2043.880 110.540 2044.140 110.800 ;
        RECT 2043.420 110.200 2043.680 110.460 ;
        RECT 1745.340 34.040 1745.600 34.300 ;
        RECT 2043.880 34.040 2044.140 34.300 ;
      LAYER met2 ;
        RECT 2046.560 1701.090 2046.840 1702.400 ;
        RECT 2044.400 1700.950 2046.840 1701.090 ;
        RECT 2044.400 1656.210 2044.540 1700.950 ;
        RECT 2046.560 1700.000 2046.840 1700.950 ;
        RECT 2043.480 1656.070 2044.540 1656.210 ;
        RECT 2043.480 1608.190 2043.620 1656.070 ;
        RECT 2043.420 1607.870 2043.680 1608.190 ;
        RECT 2043.880 1607.190 2044.140 1607.510 ;
        RECT 2043.940 1560.330 2044.080 1607.190 ;
        RECT 2043.940 1560.190 2044.540 1560.330 ;
        RECT 2044.400 1539.250 2044.540 1560.190 ;
        RECT 2043.940 1539.110 2044.540 1539.250 ;
        RECT 2043.940 1511.290 2044.080 1539.110 ;
        RECT 2043.880 1510.970 2044.140 1511.290 ;
        RECT 2043.880 1490.570 2044.140 1490.890 ;
        RECT 2043.940 1465.390 2044.080 1490.570 ;
        RECT 2043.880 1465.070 2044.140 1465.390 ;
        RECT 2043.880 1413.730 2044.140 1414.050 ;
        RECT 2043.940 1393.650 2044.080 1413.730 ;
        RECT 2043.880 1393.330 2044.140 1393.650 ;
        RECT 2043.880 1317.170 2044.140 1317.490 ;
        RECT 2043.940 1297.285 2044.080 1317.170 ;
        RECT 2043.870 1296.915 2044.150 1297.285 ;
        RECT 2044.790 1296.915 2045.070 1297.285 ;
        RECT 2044.860 1220.930 2045.000 1296.915 ;
        RECT 2043.880 1220.610 2044.140 1220.930 ;
        RECT 2044.800 1220.610 2045.060 1220.930 ;
        RECT 2043.940 1173.670 2044.080 1220.610 ;
        RECT 2043.880 1173.350 2044.140 1173.670 ;
        RECT 2043.420 1172.670 2043.680 1172.990 ;
        RECT 2043.480 1159.050 2043.620 1172.670 ;
        RECT 2043.420 1158.730 2043.680 1159.050 ;
        RECT 2043.880 1110.790 2044.140 1111.110 ;
        RECT 2043.940 1077.110 2044.080 1110.790 ;
        RECT 2043.880 1076.790 2044.140 1077.110 ;
        RECT 2043.420 1076.110 2043.680 1076.430 ;
        RECT 2043.480 1062.490 2043.620 1076.110 ;
        RECT 2043.420 1062.170 2043.680 1062.490 ;
        RECT 2043.880 1014.230 2044.140 1014.550 ;
        RECT 2043.940 980.550 2044.080 1014.230 ;
        RECT 2043.880 980.230 2044.140 980.550 ;
        RECT 2043.420 979.550 2043.680 979.870 ;
        RECT 2043.480 966.125 2043.620 979.550 ;
        RECT 2043.410 965.755 2043.690 966.125 ;
        RECT 2044.790 965.755 2045.070 966.125 ;
        RECT 2044.860 917.990 2045.000 965.755 ;
        RECT 2043.880 917.670 2044.140 917.990 ;
        RECT 2044.800 917.670 2045.060 917.990 ;
        RECT 2043.940 883.990 2044.080 917.670 ;
        RECT 2043.880 883.670 2044.140 883.990 ;
        RECT 2043.880 882.650 2044.140 882.970 ;
        RECT 2043.940 834.770 2044.080 882.650 ;
        RECT 2043.020 834.630 2044.080 834.770 ;
        RECT 2043.020 787.090 2043.160 834.630 ;
        RECT 2042.960 786.770 2043.220 787.090 ;
        RECT 2043.420 786.090 2043.680 786.410 ;
        RECT 2043.480 772.810 2043.620 786.090 ;
        RECT 2043.420 772.490 2043.680 772.810 ;
        RECT 2043.420 737.810 2043.680 738.130 ;
        RECT 2043.480 724.610 2043.620 737.810 ;
        RECT 2043.480 724.470 2044.080 724.610 ;
        RECT 2043.940 690.530 2044.080 724.470 ;
        RECT 2043.880 690.210 2044.140 690.530 ;
        RECT 2043.420 689.530 2043.680 689.850 ;
        RECT 2043.480 676.250 2043.620 689.530 ;
        RECT 2043.420 675.930 2043.680 676.250 ;
        RECT 2043.420 641.250 2043.680 641.570 ;
        RECT 2043.480 628.050 2043.620 641.250 ;
        RECT 2043.480 627.910 2044.080 628.050 ;
        RECT 2043.940 593.970 2044.080 627.910 ;
        RECT 2043.880 593.650 2044.140 593.970 ;
        RECT 2043.420 592.970 2043.680 593.290 ;
        RECT 2043.480 545.350 2043.620 592.970 ;
        RECT 2043.420 545.030 2043.680 545.350 ;
        RECT 2043.880 544.690 2044.140 545.010 ;
        RECT 2043.940 524.270 2044.080 544.690 ;
        RECT 2043.880 523.950 2044.140 524.270 ;
        RECT 2043.420 476.010 2043.680 476.330 ;
        RECT 2043.480 448.790 2043.620 476.010 ;
        RECT 2043.420 448.470 2043.680 448.790 ;
        RECT 2043.880 447.790 2044.140 448.110 ;
        RECT 2043.940 410.710 2044.080 447.790 ;
        RECT 2043.880 410.390 2044.140 410.710 ;
        RECT 2043.880 386.250 2044.140 386.570 ;
        RECT 2043.940 352.230 2044.080 386.250 ;
        RECT 2043.880 351.910 2044.140 352.230 ;
        RECT 2043.880 337.970 2044.140 338.290 ;
        RECT 2043.940 314.150 2044.080 337.970 ;
        RECT 2043.880 313.830 2044.140 314.150 ;
        RECT 2043.880 289.690 2044.140 290.010 ;
        RECT 2043.940 256.010 2044.080 289.690 ;
        RECT 2043.880 255.690 2044.140 256.010 ;
        RECT 2043.420 241.810 2043.680 242.070 ;
        RECT 2043.420 241.750 2044.080 241.810 ;
        RECT 2043.480 241.670 2044.080 241.750 ;
        RECT 2043.940 234.590 2044.080 241.670 ;
        RECT 2043.880 234.270 2044.140 234.590 ;
        RECT 2044.340 192.450 2044.600 192.770 ;
        RECT 2044.400 158.170 2044.540 192.450 ;
        RECT 2043.940 158.030 2044.540 158.170 ;
        RECT 2043.940 110.830 2044.080 158.030 ;
        RECT 2043.880 110.510 2044.140 110.830 ;
        RECT 2043.420 110.170 2043.680 110.490 ;
        RECT 2043.480 62.290 2043.620 110.170 ;
        RECT 2043.480 62.150 2044.080 62.290 ;
        RECT 2043.940 34.330 2044.080 62.150 ;
        RECT 1745.340 34.010 1745.600 34.330 ;
        RECT 2043.880 34.010 2044.140 34.330 ;
        RECT 1745.400 2.400 1745.540 34.010 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
      LAYER via2 ;
        RECT 2043.870 1296.960 2044.150 1297.240 ;
        RECT 2044.790 1296.960 2045.070 1297.240 ;
        RECT 2043.410 965.800 2043.690 966.080 ;
        RECT 2044.790 965.800 2045.070 966.080 ;
      LAYER met3 ;
        RECT 2043.845 1297.250 2044.175 1297.265 ;
        RECT 2044.765 1297.250 2045.095 1297.265 ;
        RECT 2043.845 1296.950 2045.095 1297.250 ;
        RECT 2043.845 1296.935 2044.175 1296.950 ;
        RECT 2044.765 1296.935 2045.095 1296.950 ;
        RECT 2043.385 966.090 2043.715 966.105 ;
        RECT 2044.765 966.090 2045.095 966.105 ;
        RECT 2043.385 965.790 2045.095 966.090 ;
        RECT 2043.385 965.775 2043.715 965.790 ;
        RECT 2044.765 965.775 2045.095 965.790 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1766.010 1685.960 1766.330 1686.020 ;
        RECT 2055.810 1685.960 2056.130 1686.020 ;
        RECT 1766.010 1685.820 2056.130 1685.960 ;
        RECT 1766.010 1685.760 1766.330 1685.820 ;
        RECT 2055.810 1685.760 2056.130 1685.820 ;
        RECT 1762.790 18.600 1763.110 18.660 ;
        RECT 1766.010 18.600 1766.330 18.660 ;
        RECT 1762.790 18.460 1766.330 18.600 ;
        RECT 1762.790 18.400 1763.110 18.460 ;
        RECT 1766.010 18.400 1766.330 18.460 ;
      LAYER via ;
        RECT 1766.040 1685.760 1766.300 1686.020 ;
        RECT 2055.840 1685.760 2056.100 1686.020 ;
        RECT 1762.820 18.400 1763.080 18.660 ;
        RECT 1766.040 18.400 1766.300 18.660 ;
      LAYER met2 ;
        RECT 2055.760 1700.000 2056.040 1702.400 ;
        RECT 2055.900 1686.050 2056.040 1700.000 ;
        RECT 1766.040 1685.730 1766.300 1686.050 ;
        RECT 2055.840 1685.730 2056.100 1686.050 ;
        RECT 1766.100 18.690 1766.240 1685.730 ;
        RECT 1762.820 18.370 1763.080 18.690 ;
        RECT 1766.040 18.370 1766.300 18.690 ;
        RECT 1762.880 2.400 1763.020 18.370 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2053.050 1683.920 2053.370 1683.980 ;
        RECT 2065.010 1683.920 2065.330 1683.980 ;
        RECT 2053.050 1683.780 2065.330 1683.920 ;
        RECT 2053.050 1683.720 2053.370 1683.780 ;
        RECT 2065.010 1683.720 2065.330 1683.780 ;
      LAYER via ;
        RECT 2053.080 1683.720 2053.340 1683.980 ;
        RECT 2065.040 1683.720 2065.300 1683.980 ;
      LAYER met2 ;
        RECT 2064.960 1700.000 2065.240 1702.400 ;
        RECT 2065.100 1684.010 2065.240 1700.000 ;
        RECT 2053.080 1683.690 2053.340 1684.010 ;
        RECT 2065.040 1683.690 2065.300 1684.010 ;
        RECT 2053.140 16.845 2053.280 1683.690 ;
        RECT 1780.750 16.475 1781.030 16.845 ;
        RECT 2053.070 16.475 2053.350 16.845 ;
        RECT 1780.820 2.400 1780.960 16.475 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
      LAYER via2 ;
        RECT 1780.750 16.520 1781.030 16.800 ;
        RECT 2053.070 16.520 2053.350 16.800 ;
      LAYER met3 ;
        RECT 1780.725 16.810 1781.055 16.825 ;
        RECT 2053.045 16.810 2053.375 16.825 ;
        RECT 1780.725 16.510 2053.375 16.810 ;
        RECT 1780.725 16.495 1781.055 16.510 ;
        RECT 2053.045 16.495 2053.375 16.510 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1800.510 1685.280 1800.830 1685.340 ;
        RECT 2074.210 1685.280 2074.530 1685.340 ;
        RECT 1800.510 1685.140 2074.530 1685.280 ;
        RECT 1800.510 1685.080 1800.830 1685.140 ;
        RECT 2074.210 1685.080 2074.530 1685.140 ;
      LAYER via ;
        RECT 1800.540 1685.080 1800.800 1685.340 ;
        RECT 2074.240 1685.080 2074.500 1685.340 ;
      LAYER met2 ;
        RECT 2074.160 1700.000 2074.440 1702.400 ;
        RECT 2074.300 1685.370 2074.440 1700.000 ;
        RECT 1800.540 1685.050 1800.800 1685.370 ;
        RECT 2074.240 1685.050 2074.500 1685.370 ;
        RECT 1800.600 3.130 1800.740 1685.050 ;
        RECT 1798.760 2.990 1800.740 3.130 ;
        RECT 1798.760 2.400 1798.900 2.990 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2017.245 19.805 2018.795 19.975 ;
        RECT 2041.625 19.805 2041.795 20.995 ;
        RECT 2017.245 16.405 2017.415 19.805 ;
      LAYER mcon ;
        RECT 2041.625 20.825 2041.795 20.995 ;
        RECT 2018.625 19.805 2018.795 19.975 ;
      LAYER met1 ;
        RECT 2052.590 1684.940 2052.910 1685.000 ;
        RECT 2082.030 1684.940 2082.350 1685.000 ;
        RECT 2052.590 1684.800 2082.350 1684.940 ;
        RECT 2052.590 1684.740 2052.910 1684.800 ;
        RECT 2082.030 1684.740 2082.350 1684.800 ;
        RECT 2041.565 20.980 2041.855 21.025 ;
        RECT 2041.565 20.840 2042.700 20.980 ;
        RECT 2041.565 20.795 2041.855 20.840 ;
        RECT 2042.560 20.640 2042.700 20.840 ;
        RECT 2052.590 20.640 2052.910 20.700 ;
        RECT 2042.560 20.500 2052.910 20.640 ;
        RECT 2052.590 20.440 2052.910 20.500 ;
        RECT 2018.565 19.960 2018.855 20.005 ;
        RECT 2041.565 19.960 2041.855 20.005 ;
        RECT 2018.565 19.820 2041.855 19.960 ;
        RECT 2018.565 19.775 2018.855 19.820 ;
        RECT 2041.565 19.775 2041.855 19.820 ;
        RECT 2017.185 16.560 2017.475 16.605 ;
        RECT 1851.660 16.420 2017.475 16.560 ;
        RECT 1816.610 15.540 1816.930 15.600 ;
        RECT 1851.660 15.540 1851.800 16.420 ;
        RECT 2017.185 16.375 2017.475 16.420 ;
        RECT 1816.610 15.400 1851.800 15.540 ;
        RECT 1816.610 15.340 1816.930 15.400 ;
      LAYER via ;
        RECT 2052.620 1684.740 2052.880 1685.000 ;
        RECT 2082.060 1684.740 2082.320 1685.000 ;
        RECT 2052.620 20.440 2052.880 20.700 ;
        RECT 1816.640 15.340 1816.900 15.600 ;
      LAYER met2 ;
        RECT 2083.360 1700.410 2083.640 1702.400 ;
        RECT 2082.120 1700.270 2083.640 1700.410 ;
        RECT 2082.120 1685.030 2082.260 1700.270 ;
        RECT 2083.360 1700.000 2083.640 1700.270 ;
        RECT 2052.620 1684.710 2052.880 1685.030 ;
        RECT 2082.060 1684.710 2082.320 1685.030 ;
        RECT 2052.680 20.730 2052.820 1684.710 ;
        RECT 2052.620 20.410 2052.880 20.730 ;
        RECT 1816.640 15.310 1816.900 15.630 ;
        RECT 1816.700 2.400 1816.840 15.310 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1834.550 1688.340 1834.870 1688.400 ;
        RECT 2092.610 1688.340 2092.930 1688.400 ;
        RECT 1834.550 1688.200 2092.930 1688.340 ;
        RECT 1834.550 1688.140 1834.870 1688.200 ;
        RECT 2092.610 1688.140 2092.930 1688.200 ;
      LAYER via ;
        RECT 1834.580 1688.140 1834.840 1688.400 ;
        RECT 2092.640 1688.140 2092.900 1688.400 ;
      LAYER met2 ;
        RECT 2092.560 1700.000 2092.840 1702.400 ;
        RECT 2092.700 1688.430 2092.840 1700.000 ;
        RECT 1834.580 1688.110 1834.840 1688.430 ;
        RECT 2092.640 1688.110 2092.900 1688.430 ;
        RECT 1834.640 2.400 1834.780 1688.110 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1969.405 16.065 1969.575 20.655 ;
      LAYER mcon ;
        RECT 1969.405 20.485 1969.575 20.655 ;
      LAYER met1 ;
        RECT 2067.310 1687.320 2067.630 1687.380 ;
        RECT 2101.810 1687.320 2102.130 1687.380 ;
        RECT 2067.310 1687.180 2102.130 1687.320 ;
        RECT 2067.310 1687.120 2067.630 1687.180 ;
        RECT 2101.810 1687.120 2102.130 1687.180 ;
        RECT 1969.345 20.640 1969.635 20.685 ;
        RECT 1969.345 20.500 2000.840 20.640 ;
        RECT 1969.345 20.455 1969.635 20.500 ;
        RECT 2000.700 20.300 2000.840 20.500 ;
        RECT 2017.630 20.300 2017.950 20.360 ;
        RECT 2000.700 20.160 2017.950 20.300 ;
        RECT 2017.630 20.100 2017.950 20.160 ;
        RECT 2063.170 17.240 2063.490 17.300 ;
        RECT 2067.310 17.240 2067.630 17.300 ;
        RECT 2063.170 17.100 2067.630 17.240 ;
        RECT 2063.170 17.040 2063.490 17.100 ;
        RECT 2067.310 17.040 2067.630 17.100 ;
        RECT 1852.030 16.220 1852.350 16.280 ;
        RECT 1969.345 16.220 1969.635 16.265 ;
        RECT 1852.030 16.080 1969.635 16.220 ;
        RECT 1852.030 16.020 1852.350 16.080 ;
        RECT 1969.345 16.035 1969.635 16.080 ;
        RECT 2018.090 15.540 2018.410 15.600 ;
        RECT 2018.090 15.400 2047.300 15.540 ;
        RECT 2018.090 15.340 2018.410 15.400 ;
        RECT 2047.160 15.200 2047.300 15.400 ;
        RECT 2063.170 15.200 2063.490 15.260 ;
        RECT 2047.160 15.060 2063.490 15.200 ;
        RECT 2063.170 15.000 2063.490 15.060 ;
      LAYER via ;
        RECT 2067.340 1687.120 2067.600 1687.380 ;
        RECT 2101.840 1687.120 2102.100 1687.380 ;
        RECT 2017.660 20.100 2017.920 20.360 ;
        RECT 2063.200 17.040 2063.460 17.300 ;
        RECT 2067.340 17.040 2067.600 17.300 ;
        RECT 1852.060 16.020 1852.320 16.280 ;
        RECT 2018.120 15.340 2018.380 15.600 ;
        RECT 2063.200 15.000 2063.460 15.260 ;
      LAYER met2 ;
        RECT 2101.760 1700.000 2102.040 1702.400 ;
        RECT 2101.900 1687.410 2102.040 1700.000 ;
        RECT 2067.340 1687.090 2067.600 1687.410 ;
        RECT 2101.840 1687.090 2102.100 1687.410 ;
        RECT 2017.660 20.130 2017.920 20.390 ;
        RECT 2017.660 20.070 2018.320 20.130 ;
        RECT 2017.720 19.990 2018.320 20.070 ;
        RECT 1852.060 15.990 1852.320 16.310 ;
        RECT 1852.120 2.400 1852.260 15.990 ;
        RECT 2018.180 15.630 2018.320 19.990 ;
        RECT 2067.400 17.330 2067.540 1687.090 ;
        RECT 2063.200 17.010 2063.460 17.330 ;
        RECT 2067.340 17.010 2067.600 17.330 ;
        RECT 2018.120 15.310 2018.380 15.630 ;
        RECT 2063.260 15.290 2063.400 17.010 ;
        RECT 2063.200 14.970 2063.460 15.290 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1921.105 1687.165 1921.275 1689.035 ;
        RECT 2064.625 1684.445 2064.795 1687.335 ;
      LAYER mcon ;
        RECT 1921.105 1688.865 1921.275 1689.035 ;
        RECT 2064.625 1687.165 2064.795 1687.335 ;
      LAYER met1 ;
        RECT 1876.410 1689.020 1876.730 1689.080 ;
        RECT 1921.045 1689.020 1921.335 1689.065 ;
        RECT 1876.410 1688.880 1921.335 1689.020 ;
        RECT 1876.410 1688.820 1876.730 1688.880 ;
        RECT 1921.045 1688.835 1921.335 1688.880 ;
        RECT 1921.045 1687.320 1921.335 1687.365 ;
        RECT 2064.565 1687.320 2064.855 1687.365 ;
        RECT 1921.045 1687.180 2064.855 1687.320 ;
        RECT 1921.045 1687.135 1921.335 1687.180 ;
        RECT 2064.565 1687.135 2064.855 1687.180 ;
        RECT 2064.565 1684.600 2064.855 1684.645 ;
        RECT 2109.630 1684.600 2109.950 1684.660 ;
        RECT 2064.565 1684.460 2109.950 1684.600 ;
        RECT 2064.565 1684.415 2064.855 1684.460 ;
        RECT 2109.630 1684.400 2109.950 1684.460 ;
        RECT 1869.970 15.200 1870.290 15.260 ;
        RECT 1876.410 15.200 1876.730 15.260 ;
        RECT 1869.970 15.060 1876.730 15.200 ;
        RECT 1869.970 15.000 1870.290 15.060 ;
        RECT 1876.410 15.000 1876.730 15.060 ;
      LAYER via ;
        RECT 1876.440 1688.820 1876.700 1689.080 ;
        RECT 2109.660 1684.400 2109.920 1684.660 ;
        RECT 1870.000 15.000 1870.260 15.260 ;
        RECT 1876.440 15.000 1876.700 15.260 ;
      LAYER met2 ;
        RECT 2110.960 1700.410 2111.240 1702.400 ;
        RECT 2109.720 1700.270 2111.240 1700.410 ;
        RECT 1876.440 1688.790 1876.700 1689.110 ;
        RECT 1876.500 15.290 1876.640 1688.790 ;
        RECT 2109.720 1684.690 2109.860 1700.270 ;
        RECT 2110.960 1700.000 2111.240 1700.270 ;
        RECT 2109.660 1684.370 2109.920 1684.690 ;
        RECT 1870.000 14.970 1870.260 15.290 ;
        RECT 1876.440 14.970 1876.700 15.290 ;
        RECT 1870.060 2.400 1870.200 14.970 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 751.710 67.220 752.030 67.280 ;
        RECT 1532.330 67.220 1532.650 67.280 ;
        RECT 751.710 67.080 1532.650 67.220 ;
        RECT 751.710 67.020 752.030 67.080 ;
        RECT 1532.330 67.020 1532.650 67.080 ;
      LAYER via ;
        RECT 751.740 67.020 752.000 67.280 ;
        RECT 1532.360 67.020 1532.620 67.280 ;
      LAYER met2 ;
        RECT 1532.280 1700.000 1532.560 1702.400 ;
        RECT 1532.420 67.310 1532.560 1700.000 ;
        RECT 751.740 66.990 752.000 67.310 ;
        RECT 1532.360 66.990 1532.620 67.310 ;
        RECT 751.800 16.730 751.940 66.990 ;
        RECT 746.280 16.590 751.940 16.730 ;
        RECT 746.280 2.400 746.420 16.590 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2018.165 14.705 2018.335 16.235 ;
      LAYER mcon ;
        RECT 2018.165 16.065 2018.335 16.235 ;
      LAYER met1 ;
        RECT 2066.850 1686.300 2067.170 1686.360 ;
        RECT 2066.850 1686.160 2105.720 1686.300 ;
        RECT 2066.850 1686.100 2067.170 1686.160 ;
        RECT 2105.580 1685.960 2105.720 1686.160 ;
        RECT 2120.210 1685.960 2120.530 1686.020 ;
        RECT 2105.580 1685.820 2120.530 1685.960 ;
        RECT 2120.210 1685.760 2120.530 1685.820 ;
        RECT 2018.105 16.220 2018.395 16.265 ;
        RECT 2066.850 16.220 2067.170 16.280 ;
        RECT 2018.105 16.080 2067.170 16.220 ;
        RECT 2018.105 16.035 2018.395 16.080 ;
        RECT 2066.850 16.020 2067.170 16.080 ;
        RECT 1887.910 14.860 1888.230 14.920 ;
        RECT 2018.105 14.860 2018.395 14.905 ;
        RECT 1887.910 14.720 2018.395 14.860 ;
        RECT 1887.910 14.660 1888.230 14.720 ;
        RECT 2018.105 14.675 2018.395 14.720 ;
      LAYER via ;
        RECT 2066.880 1686.100 2067.140 1686.360 ;
        RECT 2120.240 1685.760 2120.500 1686.020 ;
        RECT 2066.880 16.020 2067.140 16.280 ;
        RECT 1887.940 14.660 1888.200 14.920 ;
      LAYER met2 ;
        RECT 2120.160 1700.000 2120.440 1702.400 ;
        RECT 2066.880 1686.070 2067.140 1686.390 ;
        RECT 2066.940 16.310 2067.080 1686.070 ;
        RECT 2120.300 1686.050 2120.440 1700.000 ;
        RECT 2120.240 1685.730 2120.500 1686.050 ;
        RECT 2066.880 15.990 2067.140 16.310 ;
        RECT 1887.940 14.630 1888.200 14.950 ;
        RECT 1888.000 2.400 1888.140 14.630 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2016.325 15.725 2017.875 15.895 ;
      LAYER mcon ;
        RECT 2017.705 15.725 2017.875 15.895 ;
      LAYER met1 ;
        RECT 2121.590 1683.920 2121.910 1683.980 ;
        RECT 2129.410 1683.920 2129.730 1683.980 ;
        RECT 2121.590 1683.780 2129.730 1683.920 ;
        RECT 2121.590 1683.720 2121.910 1683.780 ;
        RECT 2129.410 1683.720 2129.730 1683.780 ;
        RECT 1905.850 15.880 1906.170 15.940 ;
        RECT 2016.265 15.880 2016.555 15.925 ;
        RECT 1905.850 15.740 2016.555 15.880 ;
        RECT 1905.850 15.680 1906.170 15.740 ;
        RECT 2016.265 15.695 2016.555 15.740 ;
        RECT 2017.645 15.880 2017.935 15.925 ;
        RECT 2017.645 15.740 2092.840 15.880 ;
        RECT 2017.645 15.695 2017.935 15.740 ;
        RECT 2092.700 15.540 2092.840 15.740 ;
        RECT 2121.590 15.540 2121.910 15.600 ;
        RECT 2092.700 15.400 2121.910 15.540 ;
        RECT 2121.590 15.340 2121.910 15.400 ;
      LAYER via ;
        RECT 2121.620 1683.720 2121.880 1683.980 ;
        RECT 2129.440 1683.720 2129.700 1683.980 ;
        RECT 1905.880 15.680 1906.140 15.940 ;
        RECT 2121.620 15.340 2121.880 15.600 ;
      LAYER met2 ;
        RECT 2129.360 1700.000 2129.640 1702.400 ;
        RECT 2129.500 1684.010 2129.640 1700.000 ;
        RECT 2121.620 1683.690 2121.880 1684.010 ;
        RECT 2129.440 1683.690 2129.700 1684.010 ;
        RECT 1905.880 15.650 1906.140 15.970 ;
        RECT 1905.940 2.400 1906.080 15.650 ;
        RECT 2121.680 15.630 2121.820 1683.690 ;
        RECT 2121.620 15.310 2121.880 15.630 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2105.105 1685.805 2105.275 1690.395 ;
        RECT 2046.225 17.085 2049.615 17.255 ;
        RECT 2046.225 14.365 2046.395 17.085 ;
        RECT 2062.785 16.575 2062.955 17.255 ;
        RECT 2067.385 16.745 2068.015 16.915 ;
        RECT 2067.385 16.575 2067.555 16.745 ;
        RECT 2062.785 16.405 2067.555 16.575 ;
      LAYER mcon ;
        RECT 2105.105 1690.225 2105.275 1690.395 ;
        RECT 2049.445 17.085 2049.615 17.255 ;
        RECT 2062.785 17.085 2062.955 17.255 ;
        RECT 2067.845 16.745 2068.015 16.915 ;
      LAYER met1 ;
        RECT 2105.045 1690.380 2105.335 1690.425 ;
        RECT 2137.230 1690.380 2137.550 1690.440 ;
        RECT 2105.045 1690.240 2137.550 1690.380 ;
        RECT 2105.045 1690.195 2105.335 1690.240 ;
        RECT 2137.230 1690.180 2137.550 1690.240 ;
        RECT 2088.010 1685.960 2088.330 1686.020 ;
        RECT 2105.045 1685.960 2105.335 1686.005 ;
        RECT 2088.010 1685.820 2105.335 1685.960 ;
        RECT 2088.010 1685.760 2088.330 1685.820 ;
        RECT 2105.045 1685.775 2105.335 1685.820 ;
        RECT 2049.385 17.240 2049.675 17.285 ;
        RECT 2062.725 17.240 2063.015 17.285 ;
        RECT 2049.385 17.100 2063.015 17.240 ;
        RECT 2049.385 17.055 2049.675 17.100 ;
        RECT 2062.725 17.055 2063.015 17.100 ;
        RECT 2067.785 16.900 2068.075 16.945 ;
        RECT 2087.090 16.900 2087.410 16.960 ;
        RECT 2067.785 16.760 2087.410 16.900 ;
        RECT 2067.785 16.715 2068.075 16.760 ;
        RECT 2087.090 16.700 2087.410 16.760 ;
        RECT 1923.330 14.520 1923.650 14.580 ;
        RECT 2046.165 14.520 2046.455 14.565 ;
        RECT 1923.330 14.380 2046.455 14.520 ;
        RECT 1923.330 14.320 1923.650 14.380 ;
        RECT 2046.165 14.335 2046.455 14.380 ;
      LAYER via ;
        RECT 2137.260 1690.180 2137.520 1690.440 ;
        RECT 2088.040 1685.760 2088.300 1686.020 ;
        RECT 2087.120 16.700 2087.380 16.960 ;
        RECT 1923.360 14.320 1923.620 14.580 ;
      LAYER met2 ;
        RECT 2138.560 1700.410 2138.840 1702.400 ;
        RECT 2137.320 1700.270 2138.840 1700.410 ;
        RECT 2137.320 1690.470 2137.460 1700.270 ;
        RECT 2138.560 1700.000 2138.840 1700.270 ;
        RECT 2137.260 1690.150 2137.520 1690.470 ;
        RECT 2088.040 1685.730 2088.300 1686.050 ;
        RECT 2088.100 1671.170 2088.240 1685.730 ;
        RECT 2087.180 1671.030 2088.240 1671.170 ;
        RECT 2087.180 16.990 2087.320 1671.030 ;
        RECT 2087.120 16.670 2087.380 16.990 ;
        RECT 1923.360 14.290 1923.620 14.610 ;
        RECT 1923.420 2.400 1923.560 14.290 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1945.410 1687.660 1945.730 1687.720 ;
        RECT 1945.410 1687.520 2114.920 1687.660 ;
        RECT 1945.410 1687.460 1945.730 1687.520 ;
        RECT 2114.780 1686.980 2114.920 1687.520 ;
        RECT 2147.810 1686.980 2148.130 1687.040 ;
        RECT 2114.780 1686.840 2148.130 1686.980 ;
        RECT 2147.810 1686.780 2148.130 1686.840 ;
        RECT 1941.270 18.260 1941.590 18.320 ;
        RECT 1945.410 18.260 1945.730 18.320 ;
        RECT 1941.270 18.120 1945.730 18.260 ;
        RECT 1941.270 18.060 1941.590 18.120 ;
        RECT 1945.410 18.060 1945.730 18.120 ;
      LAYER via ;
        RECT 1945.440 1687.460 1945.700 1687.720 ;
        RECT 2147.840 1686.780 2148.100 1687.040 ;
        RECT 1941.300 18.060 1941.560 18.320 ;
        RECT 1945.440 18.060 1945.700 18.320 ;
      LAYER met2 ;
        RECT 2147.760 1700.000 2148.040 1702.400 ;
        RECT 1945.440 1687.430 1945.700 1687.750 ;
        RECT 1945.500 18.350 1945.640 1687.430 ;
        RECT 2147.900 1687.070 2148.040 1700.000 ;
        RECT 2147.840 1686.750 2148.100 1687.070 ;
        RECT 1941.300 18.030 1941.560 18.350 ;
        RECT 1945.440 18.030 1945.700 18.350 ;
        RECT 1941.360 2.400 1941.500 18.030 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2114.305 15.725 2114.475 18.275 ;
      LAYER mcon ;
        RECT 2114.305 18.105 2114.475 18.275 ;
      LAYER met1 ;
        RECT 2152.870 1678.140 2153.190 1678.200 ;
        RECT 2155.630 1678.140 2155.950 1678.200 ;
        RECT 2152.870 1678.000 2155.950 1678.140 ;
        RECT 2152.870 1677.940 2153.190 1678.000 ;
        RECT 2155.630 1677.940 2155.950 1678.000 ;
        RECT 1959.210 18.260 1959.530 18.320 ;
        RECT 2041.550 18.260 2041.870 18.320 ;
        RECT 1959.210 18.120 2041.870 18.260 ;
        RECT 1959.210 18.060 1959.530 18.120 ;
        RECT 2041.550 18.060 2041.870 18.120 ;
        RECT 2042.930 18.260 2043.250 18.320 ;
        RECT 2114.245 18.260 2114.535 18.305 ;
        RECT 2042.930 18.120 2114.535 18.260 ;
        RECT 2042.930 18.060 2043.250 18.120 ;
        RECT 2114.245 18.075 2114.535 18.120 ;
        RECT 2114.245 15.880 2114.535 15.925 ;
        RECT 2152.870 15.880 2153.190 15.940 ;
        RECT 2114.245 15.740 2153.190 15.880 ;
        RECT 2114.245 15.695 2114.535 15.740 ;
        RECT 2152.870 15.680 2153.190 15.740 ;
      LAYER via ;
        RECT 2152.900 1677.940 2153.160 1678.200 ;
        RECT 2155.660 1677.940 2155.920 1678.200 ;
        RECT 1959.240 18.060 1959.500 18.320 ;
        RECT 2041.580 18.060 2041.840 18.320 ;
        RECT 2042.960 18.060 2043.220 18.320 ;
        RECT 2152.900 15.680 2153.160 15.940 ;
      LAYER met2 ;
        RECT 2156.960 1700.410 2157.240 1702.400 ;
        RECT 2155.720 1700.270 2157.240 1700.410 ;
        RECT 2155.720 1678.230 2155.860 1700.270 ;
        RECT 2156.960 1700.000 2157.240 1700.270 ;
        RECT 2152.900 1677.910 2153.160 1678.230 ;
        RECT 2155.660 1677.910 2155.920 1678.230 ;
        RECT 1959.240 18.030 1959.500 18.350 ;
        RECT 2041.580 18.205 2041.840 18.350 ;
        RECT 2042.960 18.205 2043.220 18.350 ;
        RECT 1959.300 2.400 1959.440 18.030 ;
        RECT 2041.570 17.835 2041.850 18.205 ;
        RECT 2042.950 17.835 2043.230 18.205 ;
        RECT 2152.960 15.970 2153.100 1677.910 ;
        RECT 2152.900 15.650 2153.160 15.970 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
      LAYER via2 ;
        RECT 2041.570 17.880 2041.850 18.160 ;
        RECT 2042.950 17.880 2043.230 18.160 ;
      LAYER met3 ;
        RECT 2041.545 18.170 2041.875 18.185 ;
        RECT 2042.925 18.170 2043.255 18.185 ;
        RECT 2041.545 17.870 2043.255 18.170 ;
        RECT 2041.545 17.855 2041.875 17.870 ;
        RECT 2042.925 17.855 2043.255 17.870 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2152.485 1685.125 2152.655 1685.975 ;
        RECT 2080.725 14.025 2080.895 20.655 ;
        RECT 2095.445 19.805 2095.615 20.655 ;
      LAYER mcon ;
        RECT 2152.485 1685.805 2152.655 1685.975 ;
        RECT 2080.725 20.485 2080.895 20.655 ;
        RECT 2095.445 20.485 2095.615 20.655 ;
      LAYER met1 ;
        RECT 2152.425 1685.960 2152.715 1686.005 ;
        RECT 2166.210 1685.960 2166.530 1686.020 ;
        RECT 2152.425 1685.820 2166.530 1685.960 ;
        RECT 2152.425 1685.775 2152.715 1685.820 ;
        RECT 2166.210 1685.760 2166.530 1685.820 ;
        RECT 2101.350 1685.280 2101.670 1685.340 ;
        RECT 2152.425 1685.280 2152.715 1685.325 ;
        RECT 2101.350 1685.140 2152.715 1685.280 ;
        RECT 2101.350 1685.080 2101.670 1685.140 ;
        RECT 2152.425 1685.095 2152.715 1685.140 ;
        RECT 2080.665 20.640 2080.955 20.685 ;
        RECT 2095.385 20.640 2095.675 20.685 ;
        RECT 2080.665 20.500 2095.675 20.640 ;
        RECT 2080.665 20.455 2080.955 20.500 ;
        RECT 2095.385 20.455 2095.675 20.500 ;
        RECT 2095.385 19.960 2095.675 20.005 ;
        RECT 2101.350 19.960 2101.670 20.020 ;
        RECT 2095.385 19.820 2101.670 19.960 ;
        RECT 2095.385 19.775 2095.675 19.820 ;
        RECT 2101.350 19.760 2101.670 19.820 ;
        RECT 1977.150 14.180 1977.470 14.240 ;
        RECT 2080.665 14.180 2080.955 14.225 ;
        RECT 1977.150 14.040 2080.955 14.180 ;
        RECT 1977.150 13.980 1977.470 14.040 ;
        RECT 2080.665 13.995 2080.955 14.040 ;
      LAYER via ;
        RECT 2166.240 1685.760 2166.500 1686.020 ;
        RECT 2101.380 1685.080 2101.640 1685.340 ;
        RECT 2101.380 19.760 2101.640 20.020 ;
        RECT 1977.180 13.980 1977.440 14.240 ;
      LAYER met2 ;
        RECT 2166.160 1700.000 2166.440 1702.400 ;
        RECT 2166.300 1686.050 2166.440 1700.000 ;
        RECT 2166.240 1685.730 2166.500 1686.050 ;
        RECT 2101.380 1685.050 2101.640 1685.370 ;
        RECT 2101.440 20.050 2101.580 1685.050 ;
        RECT 2101.380 19.730 2101.640 20.050 ;
        RECT 1977.180 13.950 1977.440 14.270 ;
        RECT 1977.240 2.400 1977.380 13.950 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1995.090 18.940 1995.410 19.000 ;
        RECT 2174.030 18.940 2174.350 19.000 ;
        RECT 1995.090 18.800 2174.350 18.940 ;
        RECT 1995.090 18.740 1995.410 18.800 ;
        RECT 2174.030 18.740 2174.350 18.800 ;
      LAYER via ;
        RECT 1995.120 18.740 1995.380 19.000 ;
        RECT 2174.060 18.740 2174.320 19.000 ;
      LAYER met2 ;
        RECT 2175.360 1700.410 2175.640 1702.400 ;
        RECT 2174.120 1700.270 2175.640 1700.410 ;
        RECT 2174.120 19.030 2174.260 1700.270 ;
        RECT 2175.360 1700.000 2175.640 1700.270 ;
        RECT 1995.120 18.710 1995.380 19.030 ;
        RECT 2174.060 18.710 2174.320 19.030 ;
        RECT 1995.180 2.400 1995.320 18.710 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2162.605 1685.125 2164.615 1685.295 ;
        RECT 2162.605 1684.785 2162.775 1685.125 ;
        RECT 2179.165 1683.765 2179.335 1685.295 ;
        RECT 2017.705 18.445 2018.795 18.615 ;
        RECT 2041.165 18.445 2041.335 21.335 ;
        RECT 2017.705 17.085 2017.875 18.445 ;
        RECT 2094.985 17.425 2095.155 19.975 ;
        RECT 2106.485 17.425 2106.655 19.975 ;
      LAYER mcon ;
        RECT 2164.445 1685.125 2164.615 1685.295 ;
        RECT 2179.165 1685.125 2179.335 1685.295 ;
        RECT 2041.165 21.165 2041.335 21.335 ;
        RECT 2018.625 18.445 2018.795 18.615 ;
        RECT 2094.985 19.805 2095.155 19.975 ;
        RECT 2106.485 19.805 2106.655 19.975 ;
      LAYER met1 ;
        RECT 2164.385 1685.280 2164.675 1685.325 ;
        RECT 2179.105 1685.280 2179.395 1685.325 ;
        RECT 2164.385 1685.140 2179.395 1685.280 ;
        RECT 2164.385 1685.095 2164.675 1685.140 ;
        RECT 2179.105 1685.095 2179.395 1685.140 ;
        RECT 2122.050 1684.940 2122.370 1685.000 ;
        RECT 2162.545 1684.940 2162.835 1684.985 ;
        RECT 2122.050 1684.800 2162.835 1684.940 ;
        RECT 2122.050 1684.740 2122.370 1684.800 ;
        RECT 2162.545 1684.755 2162.835 1684.800 ;
        RECT 2179.105 1683.920 2179.395 1683.965 ;
        RECT 2184.610 1683.920 2184.930 1683.980 ;
        RECT 2179.105 1683.780 2184.930 1683.920 ;
        RECT 2179.105 1683.735 2179.395 1683.780 ;
        RECT 2184.610 1683.720 2184.930 1683.780 ;
        RECT 2041.105 21.320 2041.395 21.365 ;
        RECT 2043.390 21.320 2043.710 21.380 ;
        RECT 2041.105 21.180 2043.710 21.320 ;
        RECT 2041.105 21.135 2041.395 21.180 ;
        RECT 2043.390 21.120 2043.710 21.180 ;
        RECT 2043.390 19.960 2043.710 20.020 ;
        RECT 2094.925 19.960 2095.215 20.005 ;
        RECT 2043.390 19.820 2095.215 19.960 ;
        RECT 2043.390 19.760 2043.710 19.820 ;
        RECT 2094.925 19.775 2095.215 19.820 ;
        RECT 2106.425 19.960 2106.715 20.005 ;
        RECT 2122.050 19.960 2122.370 20.020 ;
        RECT 2106.425 19.820 2122.370 19.960 ;
        RECT 2106.425 19.775 2106.715 19.820 ;
        RECT 2122.050 19.760 2122.370 19.820 ;
        RECT 2018.565 18.600 2018.855 18.645 ;
        RECT 2041.105 18.600 2041.395 18.645 ;
        RECT 2018.565 18.460 2041.395 18.600 ;
        RECT 2018.565 18.415 2018.855 18.460 ;
        RECT 2041.105 18.415 2041.395 18.460 ;
        RECT 2094.925 17.580 2095.215 17.625 ;
        RECT 2106.425 17.580 2106.715 17.625 ;
        RECT 2094.925 17.440 2106.715 17.580 ;
        RECT 2094.925 17.395 2095.215 17.440 ;
        RECT 2106.425 17.395 2106.715 17.440 ;
        RECT 2012.570 17.240 2012.890 17.300 ;
        RECT 2017.645 17.240 2017.935 17.285 ;
        RECT 2012.570 17.100 2017.935 17.240 ;
        RECT 2012.570 17.040 2012.890 17.100 ;
        RECT 2017.645 17.055 2017.935 17.100 ;
      LAYER via ;
        RECT 2122.080 1684.740 2122.340 1685.000 ;
        RECT 2184.640 1683.720 2184.900 1683.980 ;
        RECT 2043.420 21.120 2043.680 21.380 ;
        RECT 2043.420 19.760 2043.680 20.020 ;
        RECT 2122.080 19.760 2122.340 20.020 ;
        RECT 2012.600 17.040 2012.860 17.300 ;
      LAYER met2 ;
        RECT 2184.560 1700.000 2184.840 1702.400 ;
        RECT 2122.080 1684.710 2122.340 1685.030 ;
        RECT 2043.420 21.090 2043.680 21.410 ;
        RECT 2043.480 20.050 2043.620 21.090 ;
        RECT 2122.140 20.050 2122.280 1684.710 ;
        RECT 2184.700 1684.010 2184.840 1700.000 ;
        RECT 2184.640 1683.690 2184.900 1684.010 ;
        RECT 2043.420 19.730 2043.680 20.050 ;
        RECT 2122.080 19.730 2122.340 20.050 ;
        RECT 2012.600 17.010 2012.860 17.330 ;
        RECT 2012.660 2.400 2012.800 17.010 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2193.810 1684.940 2194.130 1685.000 ;
        RECT 2163.080 1684.800 2194.130 1684.940 ;
        RECT 2135.390 1684.600 2135.710 1684.660 ;
        RECT 2163.080 1684.600 2163.220 1684.800 ;
        RECT 2193.810 1684.740 2194.130 1684.800 ;
        RECT 2135.390 1684.460 2163.220 1684.600 ;
        RECT 2135.390 1684.400 2135.710 1684.460 ;
        RECT 2135.390 15.200 2135.710 15.260 ;
        RECT 2094.080 15.060 2135.710 15.200 ;
        RECT 2030.510 14.860 2030.830 14.920 ;
        RECT 2045.690 14.860 2046.010 14.920 ;
        RECT 2030.510 14.720 2046.010 14.860 ;
        RECT 2030.510 14.660 2030.830 14.720 ;
        RECT 2045.690 14.660 2046.010 14.720 ;
        RECT 2047.070 14.860 2047.390 14.920 ;
        RECT 2094.080 14.860 2094.220 15.060 ;
        RECT 2135.390 15.000 2135.710 15.060 ;
        RECT 2047.070 14.720 2094.220 14.860 ;
        RECT 2047.070 14.660 2047.390 14.720 ;
      LAYER via ;
        RECT 2135.420 1684.400 2135.680 1684.660 ;
        RECT 2193.840 1684.740 2194.100 1685.000 ;
        RECT 2030.540 14.660 2030.800 14.920 ;
        RECT 2045.720 14.660 2045.980 14.920 ;
        RECT 2047.100 14.660 2047.360 14.920 ;
        RECT 2135.420 15.000 2135.680 15.260 ;
      LAYER met2 ;
        RECT 2193.760 1700.000 2194.040 1702.400 ;
        RECT 2193.900 1685.030 2194.040 1700.000 ;
        RECT 2193.840 1684.710 2194.100 1685.030 ;
        RECT 2135.420 1684.370 2135.680 1684.690 ;
        RECT 2135.480 15.290 2135.620 1684.370 ;
        RECT 2135.420 14.970 2135.680 15.290 ;
        RECT 2030.540 14.630 2030.800 14.950 ;
        RECT 2045.720 14.690 2045.980 14.950 ;
        RECT 2047.100 14.690 2047.360 14.950 ;
        RECT 2045.720 14.630 2047.360 14.690 ;
        RECT 2030.600 2.400 2030.740 14.630 ;
        RECT 2045.780 14.550 2047.300 14.630 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2203.010 1684.600 2203.330 1684.660 ;
        RECT 2163.540 1684.460 2203.330 1684.600 ;
        RECT 2156.090 1684.260 2156.410 1684.320 ;
        RECT 2163.540 1684.260 2163.680 1684.460 ;
        RECT 2203.010 1684.400 2203.330 1684.460 ;
        RECT 2156.090 1684.120 2163.680 1684.260 ;
        RECT 2156.090 1684.060 2156.410 1684.120 ;
        RECT 2048.450 16.560 2048.770 16.620 ;
        RECT 2156.090 16.560 2156.410 16.620 ;
        RECT 2048.450 16.420 2156.410 16.560 ;
        RECT 2048.450 16.360 2048.770 16.420 ;
        RECT 2156.090 16.360 2156.410 16.420 ;
      LAYER via ;
        RECT 2156.120 1684.060 2156.380 1684.320 ;
        RECT 2203.040 1684.400 2203.300 1684.660 ;
        RECT 2048.480 16.360 2048.740 16.620 ;
        RECT 2156.120 16.360 2156.380 16.620 ;
      LAYER met2 ;
        RECT 2202.960 1700.000 2203.240 1702.400 ;
        RECT 2203.100 1684.690 2203.240 1700.000 ;
        RECT 2203.040 1684.370 2203.300 1684.690 ;
        RECT 2156.120 1684.030 2156.380 1684.350 ;
        RECT 2156.180 16.650 2156.320 1684.030 ;
        RECT 2048.480 16.330 2048.740 16.650 ;
        RECT 2156.120 16.330 2156.380 16.650 ;
        RECT 2048.540 2.400 2048.680 16.330 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1539.230 1678.140 1539.550 1678.200 ;
        RECT 1540.150 1678.140 1540.470 1678.200 ;
        RECT 1539.230 1678.000 1540.470 1678.140 ;
        RECT 1539.230 1677.940 1539.550 1678.000 ;
        RECT 1540.150 1677.940 1540.470 1678.000 ;
        RECT 765.510 67.900 765.830 67.960 ;
        RECT 1539.230 67.900 1539.550 67.960 ;
        RECT 765.510 67.760 1539.550 67.900 ;
        RECT 765.510 67.700 765.830 67.760 ;
        RECT 1539.230 67.700 1539.550 67.760 ;
      LAYER via ;
        RECT 1539.260 1677.940 1539.520 1678.200 ;
        RECT 1540.180 1677.940 1540.440 1678.200 ;
        RECT 765.540 67.700 765.800 67.960 ;
        RECT 1539.260 67.700 1539.520 67.960 ;
      LAYER met2 ;
        RECT 1541.480 1700.410 1541.760 1702.400 ;
        RECT 1540.240 1700.270 1541.760 1700.410 ;
        RECT 1540.240 1678.230 1540.380 1700.270 ;
        RECT 1541.480 1700.000 1541.760 1700.270 ;
        RECT 1539.260 1677.910 1539.520 1678.230 ;
        RECT 1540.180 1677.910 1540.440 1678.230 ;
        RECT 1539.320 67.990 1539.460 1677.910 ;
        RECT 765.540 67.670 765.800 67.990 ;
        RECT 1539.260 67.670 1539.520 67.990 ;
        RECT 765.600 16.730 765.740 67.670 ;
        RECT 763.760 16.590 765.740 16.730 ;
        RECT 763.760 2.400 763.900 16.590 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2071.985 2.805 2072.155 16.235 ;
        RECT 2083.945 15.385 2084.115 16.235 ;
        RECT 2091.305 15.385 2091.475 16.915 ;
      LAYER mcon ;
        RECT 2091.305 16.745 2091.475 16.915 ;
        RECT 2071.985 16.065 2072.155 16.235 ;
        RECT 2083.945 16.065 2084.115 16.235 ;
      LAYER met1 ;
        RECT 2176.790 1684.260 2177.110 1684.320 ;
        RECT 2212.210 1684.260 2212.530 1684.320 ;
        RECT 2176.790 1684.120 2212.530 1684.260 ;
        RECT 2176.790 1684.060 2177.110 1684.120 ;
        RECT 2212.210 1684.060 2212.530 1684.120 ;
        RECT 2091.245 16.900 2091.535 16.945 ;
        RECT 2176.790 16.900 2177.110 16.960 ;
        RECT 2091.245 16.760 2177.110 16.900 ;
        RECT 2091.245 16.715 2091.535 16.760 ;
        RECT 2176.790 16.700 2177.110 16.760 ;
        RECT 2071.925 16.220 2072.215 16.265 ;
        RECT 2083.885 16.220 2084.175 16.265 ;
        RECT 2071.925 16.080 2084.175 16.220 ;
        RECT 2071.925 16.035 2072.215 16.080 ;
        RECT 2083.885 16.035 2084.175 16.080 ;
        RECT 2083.885 15.540 2084.175 15.585 ;
        RECT 2091.245 15.540 2091.535 15.585 ;
        RECT 2083.885 15.400 2091.535 15.540 ;
        RECT 2083.885 15.355 2084.175 15.400 ;
        RECT 2091.245 15.355 2091.535 15.400 ;
        RECT 2066.390 2.960 2066.710 3.020 ;
        RECT 2071.925 2.960 2072.215 3.005 ;
        RECT 2066.390 2.820 2072.215 2.960 ;
        RECT 2066.390 2.760 2066.710 2.820 ;
        RECT 2071.925 2.775 2072.215 2.820 ;
      LAYER via ;
        RECT 2176.820 1684.060 2177.080 1684.320 ;
        RECT 2212.240 1684.060 2212.500 1684.320 ;
        RECT 2176.820 16.700 2177.080 16.960 ;
        RECT 2066.420 2.760 2066.680 3.020 ;
      LAYER met2 ;
        RECT 2212.160 1700.000 2212.440 1702.400 ;
        RECT 2212.300 1684.350 2212.440 1700.000 ;
        RECT 2176.820 1684.030 2177.080 1684.350 ;
        RECT 2212.240 1684.030 2212.500 1684.350 ;
        RECT 2176.880 16.990 2177.020 1684.030 ;
        RECT 2176.820 16.670 2177.080 16.990 ;
        RECT 2066.420 2.730 2066.680 3.050 ;
        RECT 2066.480 2.400 2066.620 2.730 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2190.590 1683.920 2190.910 1683.980 ;
        RECT 2221.410 1683.920 2221.730 1683.980 ;
        RECT 2190.590 1683.780 2221.730 1683.920 ;
        RECT 2190.590 1683.720 2190.910 1683.780 ;
        RECT 2221.410 1683.720 2221.730 1683.780 ;
        RECT 2084.330 16.220 2084.650 16.280 ;
        RECT 2190.590 16.220 2190.910 16.280 ;
        RECT 2084.330 16.080 2190.910 16.220 ;
        RECT 2084.330 16.020 2084.650 16.080 ;
        RECT 2190.590 16.020 2190.910 16.080 ;
      LAYER via ;
        RECT 2190.620 1683.720 2190.880 1683.980 ;
        RECT 2221.440 1683.720 2221.700 1683.980 ;
        RECT 2084.360 16.020 2084.620 16.280 ;
        RECT 2190.620 16.020 2190.880 16.280 ;
      LAYER met2 ;
        RECT 2221.360 1700.000 2221.640 1702.400 ;
        RECT 2221.500 1684.010 2221.640 1700.000 ;
        RECT 2190.620 1683.690 2190.880 1684.010 ;
        RECT 2221.440 1683.690 2221.700 1684.010 ;
        RECT 2190.680 16.310 2190.820 1683.690 ;
        RECT 2084.360 15.990 2084.620 16.310 ;
        RECT 2190.620 15.990 2190.880 16.310 ;
        RECT 2084.420 2.400 2084.560 15.990 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2104.110 1688.340 2104.430 1688.400 ;
        RECT 2230.610 1688.340 2230.930 1688.400 ;
        RECT 2104.110 1688.200 2230.930 1688.340 ;
        RECT 2104.110 1688.140 2104.430 1688.200 ;
        RECT 2230.610 1688.140 2230.930 1688.200 ;
        RECT 2101.810 20.640 2102.130 20.700 ;
        RECT 2104.110 20.640 2104.430 20.700 ;
        RECT 2101.810 20.500 2104.430 20.640 ;
        RECT 2101.810 20.440 2102.130 20.500 ;
        RECT 2104.110 20.440 2104.430 20.500 ;
      LAYER via ;
        RECT 2104.140 1688.140 2104.400 1688.400 ;
        RECT 2230.640 1688.140 2230.900 1688.400 ;
        RECT 2101.840 20.440 2102.100 20.700 ;
        RECT 2104.140 20.440 2104.400 20.700 ;
      LAYER met2 ;
        RECT 2230.560 1700.000 2230.840 1702.400 ;
        RECT 2230.700 1688.430 2230.840 1700.000 ;
        RECT 2104.140 1688.110 2104.400 1688.430 ;
        RECT 2230.640 1688.110 2230.900 1688.430 ;
        RECT 2104.200 20.730 2104.340 1688.110 ;
        RECT 2101.840 20.410 2102.100 20.730 ;
        RECT 2104.140 20.410 2104.400 20.730 ;
        RECT 2101.900 2.400 2102.040 20.410 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2124.810 1686.300 2125.130 1686.360 ;
        RECT 2239.810 1686.300 2240.130 1686.360 ;
        RECT 2124.810 1686.160 2240.130 1686.300 ;
        RECT 2124.810 1686.100 2125.130 1686.160 ;
        RECT 2239.810 1686.100 2240.130 1686.160 ;
        RECT 2119.750 20.640 2120.070 20.700 ;
        RECT 2124.810 20.640 2125.130 20.700 ;
        RECT 2119.750 20.500 2125.130 20.640 ;
        RECT 2119.750 20.440 2120.070 20.500 ;
        RECT 2124.810 20.440 2125.130 20.500 ;
      LAYER via ;
        RECT 2124.840 1686.100 2125.100 1686.360 ;
        RECT 2239.840 1686.100 2240.100 1686.360 ;
        RECT 2119.780 20.440 2120.040 20.700 ;
        RECT 2124.840 20.440 2125.100 20.700 ;
      LAYER met2 ;
        RECT 2239.760 1700.000 2240.040 1702.400 ;
        RECT 2239.900 1686.390 2240.040 1700.000 ;
        RECT 2124.840 1686.070 2125.100 1686.390 ;
        RECT 2239.840 1686.070 2240.100 1686.390 ;
        RECT 2124.900 20.730 2125.040 1686.070 ;
        RECT 2119.780 20.410 2120.040 20.730 ;
        RECT 2124.840 20.410 2125.100 20.730 ;
        RECT 2119.840 2.400 2119.980 20.410 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2163.065 19.635 2163.235 19.975 ;
        RECT 2163.065 19.465 2164.155 19.635 ;
      LAYER mcon ;
        RECT 2163.065 19.805 2163.235 19.975 ;
        RECT 2163.985 19.465 2164.155 19.635 ;
      LAYER met1 ;
        RECT 2211.290 1686.640 2211.610 1686.700 ;
        RECT 2249.010 1686.640 2249.330 1686.700 ;
        RECT 2211.290 1686.500 2249.330 1686.640 ;
        RECT 2211.290 1686.440 2211.610 1686.500 ;
        RECT 2249.010 1686.440 2249.330 1686.500 ;
        RECT 2137.690 19.960 2138.010 20.020 ;
        RECT 2163.005 19.960 2163.295 20.005 ;
        RECT 2137.690 19.820 2163.295 19.960 ;
        RECT 2137.690 19.760 2138.010 19.820 ;
        RECT 2163.005 19.775 2163.295 19.820 ;
        RECT 2163.925 19.620 2164.215 19.665 ;
        RECT 2211.290 19.620 2211.610 19.680 ;
        RECT 2163.925 19.480 2211.610 19.620 ;
        RECT 2163.925 19.435 2164.215 19.480 ;
        RECT 2211.290 19.420 2211.610 19.480 ;
      LAYER via ;
        RECT 2211.320 1686.440 2211.580 1686.700 ;
        RECT 2249.040 1686.440 2249.300 1686.700 ;
        RECT 2137.720 19.760 2137.980 20.020 ;
        RECT 2211.320 19.420 2211.580 19.680 ;
      LAYER met2 ;
        RECT 2248.960 1700.000 2249.240 1702.400 ;
        RECT 2249.100 1686.730 2249.240 1700.000 ;
        RECT 2211.320 1686.410 2211.580 1686.730 ;
        RECT 2249.040 1686.410 2249.300 1686.730 ;
        RECT 2137.720 19.730 2137.980 20.050 ;
        RECT 2137.780 2.400 2137.920 19.730 ;
        RECT 2211.380 19.710 2211.520 1686.410 ;
        RECT 2211.320 19.390 2211.580 19.710 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2258.210 1685.620 2258.530 1685.680 ;
        RECT 2164.000 1685.480 2258.530 1685.620 ;
        RECT 2159.310 1685.280 2159.630 1685.340 ;
        RECT 2164.000 1685.280 2164.140 1685.480 ;
        RECT 2258.210 1685.420 2258.530 1685.480 ;
        RECT 2159.310 1685.140 2164.140 1685.280 ;
        RECT 2159.310 1685.080 2159.630 1685.140 ;
        RECT 2155.630 20.640 2155.950 20.700 ;
        RECT 2159.310 20.640 2159.630 20.700 ;
        RECT 2155.630 20.500 2159.630 20.640 ;
        RECT 2155.630 20.440 2155.950 20.500 ;
        RECT 2159.310 20.440 2159.630 20.500 ;
      LAYER via ;
        RECT 2159.340 1685.080 2159.600 1685.340 ;
        RECT 2258.240 1685.420 2258.500 1685.680 ;
        RECT 2155.660 20.440 2155.920 20.700 ;
        RECT 2159.340 20.440 2159.600 20.700 ;
      LAYER met2 ;
        RECT 2258.160 1700.000 2258.440 1702.400 ;
        RECT 2258.300 1685.710 2258.440 1700.000 ;
        RECT 2258.240 1685.390 2258.500 1685.710 ;
        RECT 2159.340 1685.050 2159.600 1685.370 ;
        RECT 2159.400 20.730 2159.540 1685.050 ;
        RECT 2155.660 20.410 2155.920 20.730 ;
        RECT 2159.340 20.410 2159.600 20.730 ;
        RECT 2155.720 2.400 2155.860 20.410 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2267.410 1684.600 2267.730 1684.660 ;
        RECT 2235.760 1684.460 2267.730 1684.600 ;
        RECT 2232.450 1683.920 2232.770 1683.980 ;
        RECT 2235.760 1683.920 2235.900 1684.460 ;
        RECT 2267.410 1684.400 2267.730 1684.460 ;
        RECT 2232.450 1683.780 2235.900 1683.920 ;
        RECT 2232.450 1683.720 2232.770 1683.780 ;
        RECT 2172.650 18.600 2172.970 18.660 ;
        RECT 2232.450 18.600 2232.770 18.660 ;
        RECT 2172.650 18.460 2232.770 18.600 ;
        RECT 2172.650 18.400 2172.970 18.460 ;
        RECT 2232.450 18.400 2232.770 18.460 ;
      LAYER via ;
        RECT 2232.480 1683.720 2232.740 1683.980 ;
        RECT 2267.440 1684.400 2267.700 1684.660 ;
        RECT 2172.680 18.400 2172.940 18.660 ;
        RECT 2232.480 18.400 2232.740 18.660 ;
      LAYER met2 ;
        RECT 2267.360 1700.000 2267.640 1702.400 ;
        RECT 2267.500 1684.690 2267.640 1700.000 ;
        RECT 2267.440 1684.370 2267.700 1684.690 ;
        RECT 2232.480 1683.690 2232.740 1684.010 ;
        RECT 2232.540 18.690 2232.680 1683.690 ;
        RECT 2172.680 18.370 2172.940 18.690 ;
        RECT 2232.480 18.370 2232.740 18.690 ;
        RECT 2172.740 9.250 2172.880 18.370 ;
        RECT 2172.740 9.110 2173.340 9.250 ;
        RECT 2173.200 2.400 2173.340 9.110 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2238.890 1683.920 2239.210 1683.980 ;
        RECT 2276.610 1683.920 2276.930 1683.980 ;
        RECT 2238.890 1683.780 2276.930 1683.920 ;
        RECT 2238.890 1683.720 2239.210 1683.780 ;
        RECT 2276.610 1683.720 2276.930 1683.780 ;
        RECT 2191.050 18.940 2191.370 19.000 ;
        RECT 2238.890 18.940 2239.210 19.000 ;
        RECT 2191.050 18.800 2239.210 18.940 ;
        RECT 2191.050 18.740 2191.370 18.800 ;
        RECT 2238.890 18.740 2239.210 18.800 ;
      LAYER via ;
        RECT 2238.920 1683.720 2239.180 1683.980 ;
        RECT 2276.640 1683.720 2276.900 1683.980 ;
        RECT 2191.080 18.740 2191.340 19.000 ;
        RECT 2238.920 18.740 2239.180 19.000 ;
      LAYER met2 ;
        RECT 2276.560 1700.000 2276.840 1702.400 ;
        RECT 2276.700 1684.010 2276.840 1700.000 ;
        RECT 2238.920 1683.690 2239.180 1684.010 ;
        RECT 2276.640 1683.690 2276.900 1684.010 ;
        RECT 2238.980 19.030 2239.120 1683.690 ;
        RECT 2191.080 18.710 2191.340 19.030 ;
        RECT 2238.920 18.710 2239.180 19.030 ;
        RECT 2191.140 2.400 2191.280 18.710 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2246.250 1688.340 2246.570 1688.400 ;
        RECT 2285.810 1688.340 2286.130 1688.400 ;
        RECT 2246.250 1688.200 2286.130 1688.340 ;
        RECT 2246.250 1688.140 2246.570 1688.200 ;
        RECT 2285.810 1688.140 2286.130 1688.200 ;
        RECT 2208.990 16.560 2209.310 16.620 ;
        RECT 2245.790 16.560 2246.110 16.620 ;
        RECT 2208.990 16.420 2246.110 16.560 ;
        RECT 2208.990 16.360 2209.310 16.420 ;
        RECT 2245.790 16.360 2246.110 16.420 ;
      LAYER via ;
        RECT 2246.280 1688.140 2246.540 1688.400 ;
        RECT 2285.840 1688.140 2286.100 1688.400 ;
        RECT 2209.020 16.360 2209.280 16.620 ;
        RECT 2245.820 16.360 2246.080 16.620 ;
      LAYER met2 ;
        RECT 2285.760 1700.000 2286.040 1702.400 ;
        RECT 2285.900 1688.430 2286.040 1700.000 ;
        RECT 2246.280 1688.110 2246.540 1688.430 ;
        RECT 2285.840 1688.110 2286.100 1688.430 ;
        RECT 2246.340 1672.530 2246.480 1688.110 ;
        RECT 2245.880 1672.390 2246.480 1672.530 ;
        RECT 2245.880 16.650 2246.020 1672.390 ;
        RECT 2209.020 16.330 2209.280 16.650 ;
        RECT 2245.820 16.330 2246.080 16.650 ;
        RECT 2209.080 2.400 2209.220 16.330 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2259.590 1690.040 2259.910 1690.100 ;
        RECT 2295.010 1690.040 2295.330 1690.100 ;
        RECT 2259.590 1689.900 2295.330 1690.040 ;
        RECT 2259.590 1689.840 2259.910 1689.900 ;
        RECT 2295.010 1689.840 2295.330 1689.900 ;
        RECT 2226.930 15.200 2227.250 15.260 ;
        RECT 2259.590 15.200 2259.910 15.260 ;
        RECT 2226.930 15.060 2259.910 15.200 ;
        RECT 2226.930 15.000 2227.250 15.060 ;
        RECT 2259.590 15.000 2259.910 15.060 ;
      LAYER via ;
        RECT 2259.620 1689.840 2259.880 1690.100 ;
        RECT 2295.040 1689.840 2295.300 1690.100 ;
        RECT 2226.960 15.000 2227.220 15.260 ;
        RECT 2259.620 15.000 2259.880 15.260 ;
      LAYER met2 ;
        RECT 2294.960 1700.000 2295.240 1702.400 ;
        RECT 2295.100 1690.130 2295.240 1700.000 ;
        RECT 2259.620 1689.810 2259.880 1690.130 ;
        RECT 2295.040 1689.810 2295.300 1690.130 ;
        RECT 2259.680 15.290 2259.820 1689.810 ;
        RECT 2226.960 14.970 2227.220 15.290 ;
        RECT 2259.620 14.970 2259.880 15.290 ;
        RECT 2227.020 2.400 2227.160 14.970 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1547.125 1642.285 1547.295 1656.395 ;
        RECT 1546.665 1497.445 1546.835 1545.555 ;
        RECT 1546.665 1400.885 1546.835 1448.655 ;
        RECT 1546.665 1304.325 1546.835 1352.095 ;
        RECT 1546.665 1256.045 1546.835 1303.815 ;
        RECT 1546.665 1062.585 1546.835 1076.695 ;
        RECT 1547.125 1014.305 1547.295 1028.415 ;
        RECT 1546.665 966.025 1546.835 980.135 ;
        RECT 1546.665 820.845 1546.835 862.495 ;
        RECT 1546.665 614.125 1546.835 662.235 ;
        RECT 1546.665 386.325 1546.835 434.775 ;
        RECT 1547.125 241.825 1547.295 330.395 ;
        RECT 1546.665 144.925 1546.835 210.375 ;
      LAYER mcon ;
        RECT 1547.125 1656.225 1547.295 1656.395 ;
        RECT 1546.665 1545.385 1546.835 1545.555 ;
        RECT 1546.665 1448.485 1546.835 1448.655 ;
        RECT 1546.665 1351.925 1546.835 1352.095 ;
        RECT 1546.665 1303.645 1546.835 1303.815 ;
        RECT 1546.665 1076.525 1546.835 1076.695 ;
        RECT 1547.125 1028.245 1547.295 1028.415 ;
        RECT 1546.665 979.965 1546.835 980.135 ;
        RECT 1546.665 862.325 1546.835 862.495 ;
        RECT 1546.665 662.065 1546.835 662.235 ;
        RECT 1546.665 434.605 1546.835 434.775 ;
        RECT 1547.125 330.225 1547.295 330.395 ;
        RECT 1546.665 210.205 1546.835 210.375 ;
      LAYER met1 ;
        RECT 1547.065 1656.380 1547.355 1656.425 ;
        RECT 1548.430 1656.380 1548.750 1656.440 ;
        RECT 1547.065 1656.240 1548.750 1656.380 ;
        RECT 1547.065 1656.195 1547.355 1656.240 ;
        RECT 1548.430 1656.180 1548.750 1656.240 ;
        RECT 1547.050 1642.440 1547.370 1642.500 ;
        RECT 1546.855 1642.300 1547.370 1642.440 ;
        RECT 1547.050 1642.240 1547.370 1642.300 ;
        RECT 1546.590 1545.540 1546.910 1545.600 ;
        RECT 1546.395 1545.400 1546.910 1545.540 ;
        RECT 1546.590 1545.340 1546.910 1545.400 ;
        RECT 1546.605 1497.600 1546.895 1497.645 ;
        RECT 1547.050 1497.600 1547.370 1497.660 ;
        RECT 1546.605 1497.460 1547.370 1497.600 ;
        RECT 1546.605 1497.415 1546.895 1497.460 ;
        RECT 1547.050 1497.400 1547.370 1497.460 ;
        RECT 1546.590 1449.320 1546.910 1449.380 ;
        RECT 1547.970 1449.320 1548.290 1449.380 ;
        RECT 1546.590 1449.180 1548.290 1449.320 ;
        RECT 1546.590 1449.120 1546.910 1449.180 ;
        RECT 1547.970 1449.120 1548.290 1449.180 ;
        RECT 1546.590 1448.640 1546.910 1448.700 ;
        RECT 1546.395 1448.500 1546.910 1448.640 ;
        RECT 1546.590 1448.440 1546.910 1448.500 ;
        RECT 1546.605 1401.040 1546.895 1401.085 ;
        RECT 1547.050 1401.040 1547.370 1401.100 ;
        RECT 1546.605 1400.900 1547.370 1401.040 ;
        RECT 1546.605 1400.855 1546.895 1400.900 ;
        RECT 1547.050 1400.840 1547.370 1400.900 ;
        RECT 1546.590 1352.760 1546.910 1352.820 ;
        RECT 1547.970 1352.760 1548.290 1352.820 ;
        RECT 1546.590 1352.620 1548.290 1352.760 ;
        RECT 1546.590 1352.560 1546.910 1352.620 ;
        RECT 1547.970 1352.560 1548.290 1352.620 ;
        RECT 1546.590 1352.080 1546.910 1352.140 ;
        RECT 1546.395 1351.940 1546.910 1352.080 ;
        RECT 1546.590 1351.880 1546.910 1351.940 ;
        RECT 1546.605 1304.480 1546.895 1304.525 ;
        RECT 1547.050 1304.480 1547.370 1304.540 ;
        RECT 1546.605 1304.340 1547.370 1304.480 ;
        RECT 1546.605 1304.295 1546.895 1304.340 ;
        RECT 1547.050 1304.280 1547.370 1304.340 ;
        RECT 1546.605 1303.800 1546.895 1303.845 ;
        RECT 1547.050 1303.800 1547.370 1303.860 ;
        RECT 1546.605 1303.660 1547.370 1303.800 ;
        RECT 1546.605 1303.615 1546.895 1303.660 ;
        RECT 1547.050 1303.600 1547.370 1303.660 ;
        RECT 1546.590 1256.200 1546.910 1256.260 ;
        RECT 1546.395 1256.060 1546.910 1256.200 ;
        RECT 1546.590 1256.000 1546.910 1256.060 ;
        RECT 1547.510 1207.580 1547.830 1207.640 ;
        RECT 1547.970 1207.580 1548.290 1207.640 ;
        RECT 1547.510 1207.440 1548.290 1207.580 ;
        RECT 1547.510 1207.380 1547.830 1207.440 ;
        RECT 1547.970 1207.380 1548.290 1207.440 ;
        RECT 1546.590 1124.760 1546.910 1125.020 ;
        RECT 1546.680 1124.280 1546.820 1124.760 ;
        RECT 1547.050 1124.280 1547.370 1124.340 ;
        RECT 1546.680 1124.140 1547.370 1124.280 ;
        RECT 1547.050 1124.080 1547.370 1124.140 ;
        RECT 1546.590 1076.680 1546.910 1076.740 ;
        RECT 1546.395 1076.540 1546.910 1076.680 ;
        RECT 1546.590 1076.480 1546.910 1076.540 ;
        RECT 1546.605 1062.740 1546.895 1062.785 ;
        RECT 1547.050 1062.740 1547.370 1062.800 ;
        RECT 1546.605 1062.600 1547.370 1062.740 ;
        RECT 1546.605 1062.555 1546.895 1062.600 ;
        RECT 1547.050 1062.540 1547.370 1062.600 ;
        RECT 1547.050 1028.400 1547.370 1028.460 ;
        RECT 1546.855 1028.260 1547.370 1028.400 ;
        RECT 1547.050 1028.200 1547.370 1028.260 ;
        RECT 1547.050 1014.460 1547.370 1014.520 ;
        RECT 1546.855 1014.320 1547.370 1014.460 ;
        RECT 1547.050 1014.260 1547.370 1014.320 ;
        RECT 1546.590 980.120 1546.910 980.180 ;
        RECT 1546.395 979.980 1546.910 980.120 ;
        RECT 1546.590 979.920 1546.910 979.980 ;
        RECT 1546.605 966.180 1546.895 966.225 ;
        RECT 1547.050 966.180 1547.370 966.240 ;
        RECT 1546.605 966.040 1547.370 966.180 ;
        RECT 1546.605 965.995 1546.895 966.040 ;
        RECT 1547.050 965.980 1547.370 966.040 ;
        RECT 1547.050 883.900 1547.370 883.960 ;
        RECT 1546.680 883.760 1547.370 883.900 ;
        RECT 1546.680 883.280 1546.820 883.760 ;
        RECT 1547.050 883.700 1547.370 883.760 ;
        RECT 1546.590 883.020 1546.910 883.280 ;
        RECT 1546.590 862.480 1546.910 862.540 ;
        RECT 1546.395 862.340 1546.910 862.480 ;
        RECT 1546.590 862.280 1546.910 862.340 ;
        RECT 1546.590 821.000 1546.910 821.060 ;
        RECT 1546.395 820.860 1546.910 821.000 ;
        RECT 1546.590 820.800 1546.910 820.860 ;
        RECT 1546.590 765.920 1546.910 765.980 ;
        RECT 1547.510 765.920 1547.830 765.980 ;
        RECT 1546.590 765.780 1547.830 765.920 ;
        RECT 1546.590 765.720 1546.910 765.780 ;
        RECT 1547.510 765.720 1547.830 765.780 ;
        RECT 1546.590 676.500 1546.910 676.560 ;
        RECT 1547.970 676.500 1548.290 676.560 ;
        RECT 1546.590 676.360 1548.290 676.500 ;
        RECT 1546.590 676.300 1546.910 676.360 ;
        RECT 1547.970 676.300 1548.290 676.360 ;
        RECT 1546.590 662.220 1546.910 662.280 ;
        RECT 1546.395 662.080 1546.910 662.220 ;
        RECT 1546.590 662.020 1546.910 662.080 ;
        RECT 1546.605 614.280 1546.895 614.325 ;
        RECT 1547.510 614.280 1547.830 614.340 ;
        RECT 1546.605 614.140 1547.830 614.280 ;
        RECT 1546.605 614.095 1546.895 614.140 ;
        RECT 1547.510 614.080 1547.830 614.140 ;
        RECT 1546.590 566.000 1546.910 566.060 ;
        RECT 1547.510 566.000 1547.830 566.060 ;
        RECT 1546.590 565.860 1547.830 566.000 ;
        RECT 1546.590 565.800 1546.910 565.860 ;
        RECT 1547.510 565.800 1547.830 565.860 ;
        RECT 1546.590 434.760 1546.910 434.820 ;
        RECT 1546.395 434.620 1546.910 434.760 ;
        RECT 1546.590 434.560 1546.910 434.620 ;
        RECT 1546.590 386.480 1546.910 386.540 ;
        RECT 1546.395 386.340 1546.910 386.480 ;
        RECT 1546.590 386.280 1546.910 386.340 ;
        RECT 1547.050 330.860 1547.370 331.120 ;
        RECT 1547.140 330.425 1547.280 330.860 ;
        RECT 1547.065 330.195 1547.355 330.425 ;
        RECT 1547.050 241.980 1547.370 242.040 ;
        RECT 1546.855 241.840 1547.370 241.980 ;
        RECT 1547.050 241.780 1547.370 241.840 ;
        RECT 1546.605 210.360 1546.895 210.405 ;
        RECT 1547.050 210.360 1547.370 210.420 ;
        RECT 1546.605 210.220 1547.370 210.360 ;
        RECT 1546.605 210.175 1546.895 210.220 ;
        RECT 1547.050 210.160 1547.370 210.220 ;
        RECT 1546.590 145.080 1546.910 145.140 ;
        RECT 1546.395 144.940 1546.910 145.080 ;
        RECT 1546.590 144.880 1546.910 144.940 ;
        RECT 786.210 71.640 786.530 71.700 ;
        RECT 1547.050 71.640 1547.370 71.700 ;
        RECT 786.210 71.500 1547.370 71.640 ;
        RECT 786.210 71.440 786.530 71.500 ;
        RECT 1547.050 71.440 1547.370 71.500 ;
      LAYER via ;
        RECT 1548.460 1656.180 1548.720 1656.440 ;
        RECT 1547.080 1642.240 1547.340 1642.500 ;
        RECT 1546.620 1545.340 1546.880 1545.600 ;
        RECT 1547.080 1497.400 1547.340 1497.660 ;
        RECT 1546.620 1449.120 1546.880 1449.380 ;
        RECT 1548.000 1449.120 1548.260 1449.380 ;
        RECT 1546.620 1448.440 1546.880 1448.700 ;
        RECT 1547.080 1400.840 1547.340 1401.100 ;
        RECT 1546.620 1352.560 1546.880 1352.820 ;
        RECT 1548.000 1352.560 1548.260 1352.820 ;
        RECT 1546.620 1351.880 1546.880 1352.140 ;
        RECT 1547.080 1304.280 1547.340 1304.540 ;
        RECT 1547.080 1303.600 1547.340 1303.860 ;
        RECT 1546.620 1256.000 1546.880 1256.260 ;
        RECT 1547.540 1207.380 1547.800 1207.640 ;
        RECT 1548.000 1207.380 1548.260 1207.640 ;
        RECT 1546.620 1124.760 1546.880 1125.020 ;
        RECT 1547.080 1124.080 1547.340 1124.340 ;
        RECT 1546.620 1076.480 1546.880 1076.740 ;
        RECT 1547.080 1062.540 1547.340 1062.800 ;
        RECT 1547.080 1028.200 1547.340 1028.460 ;
        RECT 1547.080 1014.260 1547.340 1014.520 ;
        RECT 1546.620 979.920 1546.880 980.180 ;
        RECT 1547.080 965.980 1547.340 966.240 ;
        RECT 1547.080 883.700 1547.340 883.960 ;
        RECT 1546.620 883.020 1546.880 883.280 ;
        RECT 1546.620 862.280 1546.880 862.540 ;
        RECT 1546.620 820.800 1546.880 821.060 ;
        RECT 1546.620 765.720 1546.880 765.980 ;
        RECT 1547.540 765.720 1547.800 765.980 ;
        RECT 1546.620 676.300 1546.880 676.560 ;
        RECT 1548.000 676.300 1548.260 676.560 ;
        RECT 1546.620 662.020 1546.880 662.280 ;
        RECT 1547.540 614.080 1547.800 614.340 ;
        RECT 1546.620 565.800 1546.880 566.060 ;
        RECT 1547.540 565.800 1547.800 566.060 ;
        RECT 1546.620 434.560 1546.880 434.820 ;
        RECT 1546.620 386.280 1546.880 386.540 ;
        RECT 1547.080 330.860 1547.340 331.120 ;
        RECT 1547.080 241.780 1547.340 242.040 ;
        RECT 1547.080 210.160 1547.340 210.420 ;
        RECT 1546.620 144.880 1546.880 145.140 ;
        RECT 786.240 71.440 786.500 71.700 ;
        RECT 1547.080 71.440 1547.340 71.700 ;
      LAYER met2 ;
        RECT 1550.680 1700.410 1550.960 1702.400 ;
        RECT 1548.520 1700.270 1550.960 1700.410 ;
        RECT 1548.520 1656.470 1548.660 1700.270 ;
        RECT 1550.680 1700.000 1550.960 1700.270 ;
        RECT 1548.460 1656.150 1548.720 1656.470 ;
        RECT 1547.080 1642.210 1547.340 1642.530 ;
        RECT 1547.140 1559.650 1547.280 1642.210 ;
        RECT 1546.680 1559.510 1547.280 1559.650 ;
        RECT 1546.680 1545.630 1546.820 1559.510 ;
        RECT 1546.620 1545.310 1546.880 1545.630 ;
        RECT 1547.080 1497.370 1547.340 1497.690 ;
        RECT 1547.140 1497.205 1547.280 1497.370 ;
        RECT 1547.070 1496.835 1547.350 1497.205 ;
        RECT 1547.990 1496.835 1548.270 1497.205 ;
        RECT 1548.060 1449.410 1548.200 1496.835 ;
        RECT 1546.620 1449.090 1546.880 1449.410 ;
        RECT 1548.000 1449.090 1548.260 1449.410 ;
        RECT 1546.680 1448.730 1546.820 1449.090 ;
        RECT 1546.620 1448.410 1546.880 1448.730 ;
        RECT 1547.080 1400.810 1547.340 1401.130 ;
        RECT 1547.140 1400.645 1547.280 1400.810 ;
        RECT 1547.070 1400.275 1547.350 1400.645 ;
        RECT 1547.990 1400.275 1548.270 1400.645 ;
        RECT 1548.060 1352.850 1548.200 1400.275 ;
        RECT 1546.620 1352.530 1546.880 1352.850 ;
        RECT 1548.000 1352.530 1548.260 1352.850 ;
        RECT 1546.680 1352.170 1546.820 1352.530 ;
        RECT 1546.620 1351.850 1546.880 1352.170 ;
        RECT 1547.080 1304.250 1547.340 1304.570 ;
        RECT 1547.140 1303.890 1547.280 1304.250 ;
        RECT 1547.080 1303.570 1547.340 1303.890 ;
        RECT 1546.620 1255.970 1546.880 1256.290 ;
        RECT 1546.680 1255.805 1546.820 1255.970 ;
        RECT 1546.610 1255.435 1546.890 1255.805 ;
        RECT 1547.530 1255.435 1547.810 1255.805 ;
        RECT 1547.600 1207.670 1547.740 1255.435 ;
        RECT 1547.540 1207.350 1547.800 1207.670 ;
        RECT 1548.000 1207.350 1548.260 1207.670 ;
        RECT 1548.060 1159.810 1548.200 1207.350 ;
        RECT 1546.680 1159.670 1548.200 1159.810 ;
        RECT 1546.680 1125.050 1546.820 1159.670 ;
        RECT 1546.620 1124.730 1546.880 1125.050 ;
        RECT 1547.080 1124.050 1547.340 1124.370 ;
        RECT 1547.140 1110.850 1547.280 1124.050 ;
        RECT 1546.680 1110.710 1547.280 1110.850 ;
        RECT 1546.680 1076.770 1546.820 1110.710 ;
        RECT 1546.620 1076.450 1546.880 1076.770 ;
        RECT 1547.080 1062.510 1547.340 1062.830 ;
        RECT 1547.140 1028.490 1547.280 1062.510 ;
        RECT 1547.080 1028.170 1547.340 1028.490 ;
        RECT 1547.140 1014.550 1547.280 1014.705 ;
        RECT 1547.080 1014.290 1547.340 1014.550 ;
        RECT 1546.680 1014.230 1547.340 1014.290 ;
        RECT 1546.680 1014.150 1547.280 1014.230 ;
        RECT 1546.680 980.210 1546.820 1014.150 ;
        RECT 1546.620 979.890 1546.880 980.210 ;
        RECT 1547.080 965.950 1547.340 966.270 ;
        RECT 1547.140 932.010 1547.280 965.950 ;
        RECT 1546.220 931.870 1547.280 932.010 ;
        RECT 1546.220 919.205 1546.360 931.870 ;
        RECT 1546.150 918.835 1546.430 919.205 ;
        RECT 1547.070 918.155 1547.350 918.525 ;
        RECT 1547.140 883.990 1547.280 918.155 ;
        RECT 1547.080 883.670 1547.340 883.990 ;
        RECT 1546.620 882.990 1546.880 883.310 ;
        RECT 1546.680 862.570 1546.820 882.990 ;
        RECT 1546.620 862.250 1546.880 862.570 ;
        RECT 1546.620 820.770 1546.880 821.090 ;
        RECT 1546.680 814.370 1546.820 820.770 ;
        RECT 1546.680 814.230 1547.280 814.370 ;
        RECT 1547.140 766.090 1547.280 814.230 ;
        RECT 1546.680 766.010 1547.280 766.090 ;
        RECT 1546.620 765.950 1547.280 766.010 ;
        RECT 1546.620 765.690 1546.880 765.950 ;
        RECT 1547.540 765.690 1547.800 766.010 ;
        RECT 1546.680 765.535 1546.820 765.690 ;
        RECT 1547.600 717.810 1547.740 765.690 ;
        RECT 1547.600 717.670 1548.200 717.810 ;
        RECT 1548.060 676.590 1548.200 717.670 ;
        RECT 1546.620 676.270 1546.880 676.590 ;
        RECT 1548.000 676.270 1548.260 676.590 ;
        RECT 1546.680 662.310 1546.820 676.270 ;
        RECT 1546.620 661.990 1546.880 662.310 ;
        RECT 1547.540 614.050 1547.800 614.370 ;
        RECT 1547.600 566.090 1547.740 614.050 ;
        RECT 1546.620 565.770 1546.880 566.090 ;
        RECT 1547.540 565.770 1547.800 566.090 ;
        RECT 1546.680 507.010 1546.820 565.770 ;
        RECT 1546.220 506.870 1546.820 507.010 ;
        RECT 1546.220 496.810 1546.360 506.870 ;
        RECT 1546.220 496.670 1546.820 496.810 ;
        RECT 1546.680 434.850 1546.820 496.670 ;
        RECT 1546.620 434.530 1546.880 434.850 ;
        RECT 1546.620 386.250 1546.880 386.570 ;
        RECT 1546.680 338.370 1546.820 386.250 ;
        RECT 1546.680 338.230 1547.280 338.370 ;
        RECT 1547.140 331.150 1547.280 338.230 ;
        RECT 1547.080 330.830 1547.340 331.150 ;
        RECT 1547.080 241.750 1547.340 242.070 ;
        RECT 1547.140 210.450 1547.280 241.750 ;
        RECT 1547.080 210.130 1547.340 210.450 ;
        RECT 1546.620 144.850 1546.880 145.170 ;
        RECT 1546.680 96.290 1546.820 144.850 ;
        RECT 1546.680 96.150 1547.280 96.290 ;
        RECT 1547.140 71.730 1547.280 96.150 ;
        RECT 786.240 71.410 786.500 71.730 ;
        RECT 1547.080 71.410 1547.340 71.730 ;
        RECT 786.300 16.730 786.440 71.410 ;
        RECT 781.700 16.590 786.440 16.730 ;
        RECT 781.700 2.400 781.840 16.590 ;
        RECT 781.490 -4.800 782.050 2.400 ;
      LAYER via2 ;
        RECT 1547.070 1496.880 1547.350 1497.160 ;
        RECT 1547.990 1496.880 1548.270 1497.160 ;
        RECT 1547.070 1400.320 1547.350 1400.600 ;
        RECT 1547.990 1400.320 1548.270 1400.600 ;
        RECT 1546.610 1255.480 1546.890 1255.760 ;
        RECT 1547.530 1255.480 1547.810 1255.760 ;
        RECT 1546.150 918.880 1546.430 919.160 ;
        RECT 1547.070 918.200 1547.350 918.480 ;
      LAYER met3 ;
        RECT 1547.045 1497.170 1547.375 1497.185 ;
        RECT 1547.965 1497.170 1548.295 1497.185 ;
        RECT 1547.045 1496.870 1548.295 1497.170 ;
        RECT 1547.045 1496.855 1547.375 1496.870 ;
        RECT 1547.965 1496.855 1548.295 1496.870 ;
        RECT 1547.045 1400.610 1547.375 1400.625 ;
        RECT 1547.965 1400.610 1548.295 1400.625 ;
        RECT 1547.045 1400.310 1548.295 1400.610 ;
        RECT 1547.045 1400.295 1547.375 1400.310 ;
        RECT 1547.965 1400.295 1548.295 1400.310 ;
        RECT 1546.585 1255.770 1546.915 1255.785 ;
        RECT 1547.505 1255.770 1547.835 1255.785 ;
        RECT 1546.585 1255.470 1547.835 1255.770 ;
        RECT 1546.585 1255.455 1546.915 1255.470 ;
        RECT 1547.505 1255.455 1547.835 1255.470 ;
        RECT 1546.125 919.170 1546.455 919.185 ;
        RECT 1546.125 918.870 1548.050 919.170 ;
        RECT 1546.125 918.855 1546.455 918.870 ;
        RECT 1547.045 918.490 1547.375 918.505 ;
        RECT 1547.750 918.490 1548.050 918.870 ;
        RECT 1547.045 918.190 1548.050 918.490 ;
        RECT 1547.045 918.175 1547.375 918.190 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2266.950 1685.960 2267.270 1686.020 ;
        RECT 2303.750 1685.960 2304.070 1686.020 ;
        RECT 2266.950 1685.820 2304.070 1685.960 ;
        RECT 2266.950 1685.760 2267.270 1685.820 ;
        RECT 2303.750 1685.760 2304.070 1685.820 ;
        RECT 2244.870 19.280 2245.190 19.340 ;
        RECT 2266.950 19.280 2267.270 19.340 ;
        RECT 2244.870 19.140 2267.270 19.280 ;
        RECT 2244.870 19.080 2245.190 19.140 ;
        RECT 2266.950 19.080 2267.270 19.140 ;
      LAYER via ;
        RECT 2266.980 1685.760 2267.240 1686.020 ;
        RECT 2303.780 1685.760 2304.040 1686.020 ;
        RECT 2244.900 19.080 2245.160 19.340 ;
        RECT 2266.980 19.080 2267.240 19.340 ;
      LAYER met2 ;
        RECT 2303.700 1700.000 2303.980 1702.400 ;
        RECT 2303.840 1686.050 2303.980 1700.000 ;
        RECT 2266.980 1685.730 2267.240 1686.050 ;
        RECT 2303.780 1685.730 2304.040 1686.050 ;
        RECT 2267.040 19.370 2267.180 1685.730 ;
        RECT 2244.900 19.050 2245.160 19.370 ;
        RECT 2266.980 19.050 2267.240 19.370 ;
        RECT 2244.960 2.400 2245.100 19.050 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2287.190 1683.920 2287.510 1683.980 ;
        RECT 2312.950 1683.920 2313.270 1683.980 ;
        RECT 2287.190 1683.780 2313.270 1683.920 ;
        RECT 2287.190 1683.720 2287.510 1683.780 ;
        RECT 2312.950 1683.720 2313.270 1683.780 ;
        RECT 2262.350 17.240 2262.670 17.300 ;
        RECT 2287.190 17.240 2287.510 17.300 ;
        RECT 2262.350 17.100 2287.510 17.240 ;
        RECT 2262.350 17.040 2262.670 17.100 ;
        RECT 2287.190 17.040 2287.510 17.100 ;
      LAYER via ;
        RECT 2287.220 1683.720 2287.480 1683.980 ;
        RECT 2312.980 1683.720 2313.240 1683.980 ;
        RECT 2262.380 17.040 2262.640 17.300 ;
        RECT 2287.220 17.040 2287.480 17.300 ;
      LAYER met2 ;
        RECT 2312.900 1700.000 2313.180 1702.400 ;
        RECT 2313.040 1684.010 2313.180 1700.000 ;
        RECT 2287.220 1683.690 2287.480 1684.010 ;
        RECT 2312.980 1683.690 2313.240 1684.010 ;
        RECT 2287.280 17.330 2287.420 1683.690 ;
        RECT 2262.380 17.010 2262.640 17.330 ;
        RECT 2287.220 17.010 2287.480 17.330 ;
        RECT 2262.440 2.400 2262.580 17.010 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2300.990 1684.600 2301.310 1684.660 ;
        RECT 2322.150 1684.600 2322.470 1684.660 ;
        RECT 2300.990 1684.460 2322.470 1684.600 ;
        RECT 2300.990 1684.400 2301.310 1684.460 ;
        RECT 2322.150 1684.400 2322.470 1684.460 ;
        RECT 2300.990 14.180 2301.310 14.240 ;
        RECT 2280.380 14.040 2301.310 14.180 ;
        RECT 2280.380 13.900 2280.520 14.040 ;
        RECT 2300.990 13.980 2301.310 14.040 ;
        RECT 2280.290 13.640 2280.610 13.900 ;
      LAYER via ;
        RECT 2301.020 1684.400 2301.280 1684.660 ;
        RECT 2322.180 1684.400 2322.440 1684.660 ;
        RECT 2301.020 13.980 2301.280 14.240 ;
        RECT 2280.320 13.640 2280.580 13.900 ;
      LAYER met2 ;
        RECT 2322.100 1700.000 2322.380 1702.400 ;
        RECT 2322.240 1684.690 2322.380 1700.000 ;
        RECT 2301.020 1684.370 2301.280 1684.690 ;
        RECT 2322.180 1684.370 2322.440 1684.690 ;
        RECT 2301.080 14.270 2301.220 1684.370 ;
        RECT 2301.020 13.950 2301.280 14.270 ;
        RECT 2280.320 13.610 2280.580 13.930 ;
        RECT 2280.380 2.400 2280.520 13.610 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2321.690 1684.260 2322.010 1684.320 ;
        RECT 2331.350 1684.260 2331.670 1684.320 ;
        RECT 2321.690 1684.120 2331.670 1684.260 ;
        RECT 2321.690 1684.060 2322.010 1684.120 ;
        RECT 2331.350 1684.060 2331.670 1684.120 ;
        RECT 2298.230 16.900 2298.550 16.960 ;
        RECT 2321.690 16.900 2322.010 16.960 ;
        RECT 2298.230 16.760 2322.010 16.900 ;
        RECT 2298.230 16.700 2298.550 16.760 ;
        RECT 2321.690 16.700 2322.010 16.760 ;
      LAYER via ;
        RECT 2321.720 1684.060 2321.980 1684.320 ;
        RECT 2331.380 1684.060 2331.640 1684.320 ;
        RECT 2298.260 16.700 2298.520 16.960 ;
        RECT 2321.720 16.700 2321.980 16.960 ;
      LAYER met2 ;
        RECT 2331.300 1700.000 2331.580 1702.400 ;
        RECT 2331.440 1684.350 2331.580 1700.000 ;
        RECT 2321.720 1684.030 2321.980 1684.350 ;
        RECT 2331.380 1684.030 2331.640 1684.350 ;
        RECT 2321.780 16.990 2321.920 1684.030 ;
        RECT 2298.260 16.670 2298.520 16.990 ;
        RECT 2321.720 16.670 2321.980 16.990 ;
        RECT 2298.320 2.400 2298.460 16.670 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2318.010 1689.360 2318.330 1689.420 ;
        RECT 2340.550 1689.360 2340.870 1689.420 ;
        RECT 2318.010 1689.220 2340.870 1689.360 ;
        RECT 2318.010 1689.160 2318.330 1689.220 ;
        RECT 2340.550 1689.160 2340.870 1689.220 ;
        RECT 2316.170 14.180 2316.490 14.240 ;
        RECT 2318.010 14.180 2318.330 14.240 ;
        RECT 2316.170 14.040 2318.330 14.180 ;
        RECT 2316.170 13.980 2316.490 14.040 ;
        RECT 2318.010 13.980 2318.330 14.040 ;
      LAYER via ;
        RECT 2318.040 1689.160 2318.300 1689.420 ;
        RECT 2340.580 1689.160 2340.840 1689.420 ;
        RECT 2316.200 13.980 2316.460 14.240 ;
        RECT 2318.040 13.980 2318.300 14.240 ;
      LAYER met2 ;
        RECT 2340.500 1700.000 2340.780 1702.400 ;
        RECT 2340.640 1689.450 2340.780 1700.000 ;
        RECT 2318.040 1689.130 2318.300 1689.450 ;
        RECT 2340.580 1689.130 2340.840 1689.450 ;
        RECT 2318.100 14.270 2318.240 1689.130 ;
        RECT 2316.200 13.950 2316.460 14.270 ;
        RECT 2318.040 13.950 2318.300 14.270 ;
        RECT 2316.260 2.400 2316.400 13.950 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2338.710 1684.260 2339.030 1684.320 ;
        RECT 2349.750 1684.260 2350.070 1684.320 ;
        RECT 2338.710 1684.120 2350.070 1684.260 ;
        RECT 2338.710 1684.060 2339.030 1684.120 ;
        RECT 2349.750 1684.060 2350.070 1684.120 ;
        RECT 2334.110 18.600 2334.430 18.660 ;
        RECT 2338.710 18.600 2339.030 18.660 ;
        RECT 2334.110 18.460 2339.030 18.600 ;
        RECT 2334.110 18.400 2334.430 18.460 ;
        RECT 2338.710 18.400 2339.030 18.460 ;
      LAYER via ;
        RECT 2338.740 1684.060 2339.000 1684.320 ;
        RECT 2349.780 1684.060 2350.040 1684.320 ;
        RECT 2334.140 18.400 2334.400 18.660 ;
        RECT 2338.740 18.400 2339.000 18.660 ;
      LAYER met2 ;
        RECT 2349.700 1700.000 2349.980 1702.400 ;
        RECT 2349.840 1684.350 2349.980 1700.000 ;
        RECT 2338.740 1684.030 2339.000 1684.350 ;
        RECT 2349.780 1684.030 2350.040 1684.350 ;
        RECT 2338.800 18.690 2338.940 1684.030 ;
        RECT 2334.140 18.370 2334.400 18.690 ;
        RECT 2338.740 18.370 2339.000 18.690 ;
        RECT 2334.200 2.400 2334.340 18.370 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2353.430 1678.140 2353.750 1678.200 ;
        RECT 2357.110 1678.140 2357.430 1678.200 ;
        RECT 2353.430 1678.000 2357.430 1678.140 ;
        RECT 2353.430 1677.940 2353.750 1678.000 ;
        RECT 2357.110 1677.940 2357.430 1678.000 ;
        RECT 2351.590 15.540 2351.910 15.600 ;
        RECT 2353.430 15.540 2353.750 15.600 ;
        RECT 2351.590 15.400 2353.750 15.540 ;
        RECT 2351.590 15.340 2351.910 15.400 ;
        RECT 2353.430 15.340 2353.750 15.400 ;
      LAYER via ;
        RECT 2353.460 1677.940 2353.720 1678.200 ;
        RECT 2357.140 1677.940 2357.400 1678.200 ;
        RECT 2351.620 15.340 2351.880 15.600 ;
        RECT 2353.460 15.340 2353.720 15.600 ;
      LAYER met2 ;
        RECT 2358.900 1700.410 2359.180 1702.400 ;
        RECT 2357.200 1700.270 2359.180 1700.410 ;
        RECT 2357.200 1678.230 2357.340 1700.270 ;
        RECT 2358.900 1700.000 2359.180 1700.270 ;
        RECT 2353.460 1677.910 2353.720 1678.230 ;
        RECT 2357.140 1677.910 2357.400 1678.230 ;
        RECT 2353.520 15.630 2353.660 1677.910 ;
        RECT 2351.620 15.310 2351.880 15.630 ;
        RECT 2353.460 15.310 2353.720 15.630 ;
        RECT 2351.680 2.400 2351.820 15.310 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2366.770 20.640 2367.090 20.700 ;
        RECT 2369.530 20.640 2369.850 20.700 ;
        RECT 2366.770 20.500 2369.850 20.640 ;
        RECT 2366.770 20.440 2367.090 20.500 ;
        RECT 2369.530 20.440 2369.850 20.500 ;
      LAYER via ;
        RECT 2366.800 20.440 2367.060 20.700 ;
        RECT 2369.560 20.440 2369.820 20.700 ;
      LAYER met2 ;
        RECT 2368.100 1700.410 2368.380 1702.400 ;
        RECT 2366.860 1700.270 2368.380 1700.410 ;
        RECT 2366.860 20.730 2367.000 1700.270 ;
        RECT 2368.100 1700.000 2368.380 1700.270 ;
        RECT 2366.800 20.410 2367.060 20.730 ;
        RECT 2369.560 20.410 2369.820 20.730 ;
        RECT 2369.620 2.400 2369.760 20.410 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2377.350 1688.340 2377.670 1688.400 ;
        RECT 2387.930 1688.340 2388.250 1688.400 ;
        RECT 2377.350 1688.200 2388.250 1688.340 ;
        RECT 2377.350 1688.140 2377.670 1688.200 ;
        RECT 2387.930 1688.140 2388.250 1688.200 ;
      LAYER via ;
        RECT 2377.380 1688.140 2377.640 1688.400 ;
        RECT 2387.960 1688.140 2388.220 1688.400 ;
      LAYER met2 ;
        RECT 2377.300 1700.000 2377.580 1702.400 ;
        RECT 2377.440 1688.430 2377.580 1700.000 ;
        RECT 2377.380 1688.110 2377.640 1688.430 ;
        RECT 2387.960 1688.110 2388.220 1688.430 ;
        RECT 2388.020 17.410 2388.160 1688.110 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.400 2387.700 17.270 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2386.550 1690.040 2386.870 1690.100 ;
        RECT 2401.270 1690.040 2401.590 1690.100 ;
        RECT 2386.550 1689.900 2401.590 1690.040 ;
        RECT 2386.550 1689.840 2386.870 1689.900 ;
        RECT 2401.270 1689.840 2401.590 1689.900 ;
        RECT 2401.730 2.960 2402.050 3.020 ;
        RECT 2405.410 2.960 2405.730 3.020 ;
        RECT 2401.730 2.820 2405.730 2.960 ;
        RECT 2401.730 2.760 2402.050 2.820 ;
        RECT 2405.410 2.760 2405.730 2.820 ;
      LAYER via ;
        RECT 2386.580 1689.840 2386.840 1690.100 ;
        RECT 2401.300 1689.840 2401.560 1690.100 ;
        RECT 2401.760 2.760 2402.020 3.020 ;
        RECT 2405.440 2.760 2405.700 3.020 ;
      LAYER met2 ;
        RECT 2386.500 1700.000 2386.780 1702.400 ;
        RECT 2386.640 1690.130 2386.780 1700.000 ;
        RECT 2386.580 1689.810 2386.840 1690.130 ;
        RECT 2401.300 1689.810 2401.560 1690.130 ;
        RECT 2401.360 1688.170 2401.500 1689.810 ;
        RECT 2401.360 1688.030 2401.960 1688.170 ;
        RECT 2401.820 3.050 2401.960 1688.030 ;
        RECT 2401.760 2.730 2402.020 3.050 ;
        RECT 2405.440 2.730 2405.700 3.050 ;
        RECT 2405.500 2.400 2405.640 2.730 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 800.010 71.980 800.330 72.040 ;
        RECT 1559.930 71.980 1560.250 72.040 ;
        RECT 800.010 71.840 1560.250 71.980 ;
        RECT 800.010 71.780 800.330 71.840 ;
        RECT 1559.930 71.780 1560.250 71.840 ;
      LAYER via ;
        RECT 800.040 71.780 800.300 72.040 ;
        RECT 1559.960 71.780 1560.220 72.040 ;
      LAYER met2 ;
        RECT 1559.880 1700.000 1560.160 1702.400 ;
        RECT 1560.020 72.070 1560.160 1700.000 ;
        RECT 800.040 71.750 800.300 72.070 ;
        RECT 1559.960 71.750 1560.220 72.070 ;
        RECT 800.100 17.410 800.240 71.750 ;
        RECT 799.640 17.270 800.240 17.410 ;
        RECT 799.640 2.400 799.780 17.270 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1478.125 1642.285 1478.295 1690.395 ;
        RECT 1478.585 1466.165 1478.755 1490.475 ;
        RECT 1477.205 1345.465 1477.375 1393.575 ;
        RECT 1477.205 1200.285 1477.375 1297.015 ;
        RECT 1477.665 1138.745 1477.835 1186.855 ;
        RECT 1477.205 1055.445 1477.375 1077.035 ;
        RECT 1478.125 917.745 1478.295 942.395 ;
        RECT 1477.665 807.245 1477.835 855.355 ;
        RECT 1478.125 703.885 1478.295 751.995 ;
        RECT 1477.665 607.325 1477.835 655.435 ;
        RECT 1478.125 510.765 1478.295 558.875 ;
      LAYER mcon ;
        RECT 1478.125 1690.225 1478.295 1690.395 ;
        RECT 1478.585 1490.305 1478.755 1490.475 ;
        RECT 1477.205 1393.405 1477.375 1393.575 ;
        RECT 1477.205 1296.845 1477.375 1297.015 ;
        RECT 1477.665 1186.685 1477.835 1186.855 ;
        RECT 1477.205 1076.865 1477.375 1077.035 ;
        RECT 1478.125 942.225 1478.295 942.395 ;
        RECT 1477.665 855.185 1477.835 855.355 ;
        RECT 1478.125 751.825 1478.295 751.995 ;
        RECT 1477.665 655.265 1477.835 655.435 ;
        RECT 1478.125 558.705 1478.295 558.875 ;
      LAYER met1 ;
        RECT 1478.065 1690.380 1478.355 1690.425 ;
        RECT 1478.970 1690.380 1479.290 1690.440 ;
        RECT 1478.065 1690.240 1479.290 1690.380 ;
        RECT 1478.065 1690.195 1478.355 1690.240 ;
        RECT 1478.970 1690.180 1479.290 1690.240 ;
        RECT 1478.050 1642.440 1478.370 1642.500 ;
        RECT 1477.855 1642.300 1478.370 1642.440 ;
        RECT 1478.050 1642.240 1478.370 1642.300 ;
        RECT 1478.510 1490.460 1478.830 1490.520 ;
        RECT 1478.315 1490.320 1478.830 1490.460 ;
        RECT 1478.510 1490.260 1478.830 1490.320 ;
        RECT 1478.510 1466.320 1478.830 1466.380 ;
        RECT 1478.315 1466.180 1478.830 1466.320 ;
        RECT 1478.510 1466.120 1478.830 1466.180 ;
        RECT 1477.130 1400.700 1477.450 1400.760 ;
        RECT 1478.510 1400.700 1478.830 1400.760 ;
        RECT 1477.130 1400.560 1478.830 1400.700 ;
        RECT 1477.130 1400.500 1477.450 1400.560 ;
        RECT 1478.510 1400.500 1478.830 1400.560 ;
        RECT 1477.130 1393.560 1477.450 1393.620 ;
        RECT 1476.935 1393.420 1477.450 1393.560 ;
        RECT 1477.130 1393.360 1477.450 1393.420 ;
        RECT 1477.145 1345.620 1477.435 1345.665 ;
        RECT 1478.050 1345.620 1478.370 1345.680 ;
        RECT 1477.145 1345.480 1478.370 1345.620 ;
        RECT 1477.145 1345.435 1477.435 1345.480 ;
        RECT 1478.050 1345.420 1478.370 1345.480 ;
        RECT 1477.130 1304.140 1477.450 1304.200 ;
        RECT 1478.050 1304.140 1478.370 1304.200 ;
        RECT 1477.130 1304.000 1478.370 1304.140 ;
        RECT 1477.130 1303.940 1477.450 1304.000 ;
        RECT 1478.050 1303.940 1478.370 1304.000 ;
        RECT 1477.130 1297.000 1477.450 1297.060 ;
        RECT 1476.935 1296.860 1477.450 1297.000 ;
        RECT 1477.130 1296.800 1477.450 1296.860 ;
        RECT 1477.145 1200.440 1477.435 1200.485 ;
        RECT 1477.590 1200.440 1477.910 1200.500 ;
        RECT 1477.145 1200.300 1477.910 1200.440 ;
        RECT 1477.145 1200.255 1477.435 1200.300 ;
        RECT 1477.590 1200.240 1477.910 1200.300 ;
        RECT 1477.590 1186.840 1477.910 1186.900 ;
        RECT 1477.395 1186.700 1477.910 1186.840 ;
        RECT 1477.590 1186.640 1477.910 1186.700 ;
        RECT 1477.590 1138.900 1477.910 1138.960 ;
        RECT 1477.395 1138.760 1477.910 1138.900 ;
        RECT 1477.590 1138.700 1477.910 1138.760 ;
        RECT 1477.590 1124.760 1477.910 1125.020 ;
        RECT 1477.680 1124.280 1477.820 1124.760 ;
        RECT 1478.050 1124.280 1478.370 1124.340 ;
        RECT 1477.680 1124.140 1478.370 1124.280 ;
        RECT 1478.050 1124.080 1478.370 1124.140 ;
        RECT 1477.145 1077.020 1477.435 1077.065 ;
        RECT 1478.050 1077.020 1478.370 1077.080 ;
        RECT 1477.145 1076.880 1478.370 1077.020 ;
        RECT 1477.145 1076.835 1477.435 1076.880 ;
        RECT 1478.050 1076.820 1478.370 1076.880 ;
        RECT 1477.130 1055.600 1477.450 1055.660 ;
        RECT 1476.935 1055.460 1477.450 1055.600 ;
        RECT 1477.130 1055.400 1477.450 1055.460 ;
        RECT 1477.130 1031.460 1477.450 1031.520 ;
        RECT 1478.510 1031.460 1478.830 1031.520 ;
        RECT 1477.130 1031.320 1478.830 1031.460 ;
        RECT 1477.130 1031.260 1477.450 1031.320 ;
        RECT 1478.510 1031.260 1478.830 1031.320 ;
        RECT 1477.130 1000.520 1477.450 1000.580 ;
        RECT 1478.510 1000.520 1478.830 1000.580 ;
        RECT 1477.130 1000.380 1478.830 1000.520 ;
        RECT 1477.130 1000.320 1477.450 1000.380 ;
        RECT 1478.510 1000.320 1478.830 1000.380 ;
        RECT 1478.050 942.380 1478.370 942.440 ;
        RECT 1477.855 942.240 1478.370 942.380 ;
        RECT 1478.050 942.180 1478.370 942.240 ;
        RECT 1478.050 917.900 1478.370 917.960 ;
        RECT 1477.855 917.760 1478.370 917.900 ;
        RECT 1478.050 917.700 1478.370 917.760 ;
        RECT 1477.590 855.340 1477.910 855.400 ;
        RECT 1477.395 855.200 1477.910 855.340 ;
        RECT 1477.590 855.140 1477.910 855.200 ;
        RECT 1477.590 807.400 1477.910 807.460 ;
        RECT 1477.395 807.260 1477.910 807.400 ;
        RECT 1477.590 807.200 1477.910 807.260 ;
        RECT 1478.050 759.120 1478.370 759.180 ;
        RECT 1478.050 758.980 1478.740 759.120 ;
        RECT 1478.050 758.920 1478.370 758.980 ;
        RECT 1478.600 758.500 1478.740 758.980 ;
        RECT 1478.510 758.240 1478.830 758.500 ;
        RECT 1478.065 751.980 1478.355 752.025 ;
        RECT 1478.510 751.980 1478.830 752.040 ;
        RECT 1478.065 751.840 1478.830 751.980 ;
        RECT 1478.065 751.795 1478.355 751.840 ;
        RECT 1478.510 751.780 1478.830 751.840 ;
        RECT 1478.050 704.040 1478.370 704.100 ;
        RECT 1477.855 703.900 1478.370 704.040 ;
        RECT 1478.050 703.840 1478.370 703.900 ;
        RECT 1477.590 655.420 1477.910 655.480 ;
        RECT 1477.395 655.280 1477.910 655.420 ;
        RECT 1477.590 655.220 1477.910 655.280 ;
        RECT 1477.605 607.480 1477.895 607.525 ;
        RECT 1478.050 607.480 1478.370 607.540 ;
        RECT 1477.605 607.340 1478.370 607.480 ;
        RECT 1477.605 607.295 1477.895 607.340 ;
        RECT 1478.050 607.280 1478.370 607.340 ;
        RECT 1478.050 593.680 1478.370 593.940 ;
        RECT 1478.140 593.260 1478.280 593.680 ;
        RECT 1478.050 593.000 1478.370 593.260 ;
        RECT 1478.050 558.860 1478.370 558.920 ;
        RECT 1477.855 558.720 1478.370 558.860 ;
        RECT 1478.050 558.660 1478.370 558.720 ;
        RECT 1478.065 510.920 1478.355 510.965 ;
        RECT 1478.510 510.920 1478.830 510.980 ;
        RECT 1478.065 510.780 1478.830 510.920 ;
        RECT 1478.065 510.735 1478.355 510.780 ;
        RECT 1478.510 510.720 1478.830 510.780 ;
        RECT 1477.590 400.760 1477.910 400.820 ;
        RECT 1478.510 400.760 1478.830 400.820 ;
        RECT 1477.590 400.620 1478.830 400.760 ;
        RECT 1477.590 400.560 1477.910 400.620 ;
        RECT 1478.510 400.560 1478.830 400.620 ;
        RECT 1477.590 289.720 1477.910 289.980 ;
        RECT 1477.680 289.240 1477.820 289.720 ;
        RECT 1478.050 289.240 1478.370 289.300 ;
        RECT 1477.680 289.100 1478.370 289.240 ;
        RECT 1478.050 289.040 1478.370 289.100 ;
        RECT 1478.050 241.300 1478.370 241.360 ;
        RECT 1478.510 241.300 1478.830 241.360 ;
        RECT 1478.050 241.160 1478.830 241.300 ;
        RECT 1478.050 241.100 1478.370 241.160 ;
        RECT 1478.510 241.100 1478.830 241.160 ;
        RECT 1478.510 191.460 1478.830 191.720 ;
        RECT 1478.600 191.040 1478.740 191.460 ;
        RECT 1478.510 190.780 1478.830 191.040 ;
        RECT 1477.590 144.740 1477.910 144.800 ;
        RECT 1478.050 144.740 1478.370 144.800 ;
        RECT 1477.590 144.600 1478.370 144.740 ;
        RECT 1477.590 144.540 1477.910 144.600 ;
        RECT 1478.050 144.540 1478.370 144.600 ;
        RECT 648.210 75.720 648.530 75.780 ;
        RECT 1477.590 75.720 1477.910 75.780 ;
        RECT 648.210 75.580 1477.910 75.720 ;
        RECT 648.210 75.520 648.530 75.580 ;
        RECT 1477.590 75.520 1477.910 75.580 ;
      LAYER via ;
        RECT 1479.000 1690.180 1479.260 1690.440 ;
        RECT 1478.080 1642.240 1478.340 1642.500 ;
        RECT 1478.540 1490.260 1478.800 1490.520 ;
        RECT 1478.540 1466.120 1478.800 1466.380 ;
        RECT 1477.160 1400.500 1477.420 1400.760 ;
        RECT 1478.540 1400.500 1478.800 1400.760 ;
        RECT 1477.160 1393.360 1477.420 1393.620 ;
        RECT 1478.080 1345.420 1478.340 1345.680 ;
        RECT 1477.160 1303.940 1477.420 1304.200 ;
        RECT 1478.080 1303.940 1478.340 1304.200 ;
        RECT 1477.160 1296.800 1477.420 1297.060 ;
        RECT 1477.620 1200.240 1477.880 1200.500 ;
        RECT 1477.620 1186.640 1477.880 1186.900 ;
        RECT 1477.620 1138.700 1477.880 1138.960 ;
        RECT 1477.620 1124.760 1477.880 1125.020 ;
        RECT 1478.080 1124.080 1478.340 1124.340 ;
        RECT 1478.080 1076.820 1478.340 1077.080 ;
        RECT 1477.160 1055.400 1477.420 1055.660 ;
        RECT 1477.160 1031.260 1477.420 1031.520 ;
        RECT 1478.540 1031.260 1478.800 1031.520 ;
        RECT 1477.160 1000.320 1477.420 1000.580 ;
        RECT 1478.540 1000.320 1478.800 1000.580 ;
        RECT 1478.080 942.180 1478.340 942.440 ;
        RECT 1478.080 917.700 1478.340 917.960 ;
        RECT 1477.620 855.140 1477.880 855.400 ;
        RECT 1477.620 807.200 1477.880 807.460 ;
        RECT 1478.080 758.920 1478.340 759.180 ;
        RECT 1478.540 758.240 1478.800 758.500 ;
        RECT 1478.540 751.780 1478.800 752.040 ;
        RECT 1478.080 703.840 1478.340 704.100 ;
        RECT 1477.620 655.220 1477.880 655.480 ;
        RECT 1478.080 607.280 1478.340 607.540 ;
        RECT 1478.080 593.680 1478.340 593.940 ;
        RECT 1478.080 593.000 1478.340 593.260 ;
        RECT 1478.080 558.660 1478.340 558.920 ;
        RECT 1478.540 510.720 1478.800 510.980 ;
        RECT 1477.620 400.560 1477.880 400.820 ;
        RECT 1478.540 400.560 1478.800 400.820 ;
        RECT 1477.620 289.720 1477.880 289.980 ;
        RECT 1478.080 289.040 1478.340 289.300 ;
        RECT 1478.080 241.100 1478.340 241.360 ;
        RECT 1478.540 241.100 1478.800 241.360 ;
        RECT 1478.540 191.460 1478.800 191.720 ;
        RECT 1478.540 190.780 1478.800 191.040 ;
        RECT 1477.620 144.540 1477.880 144.800 ;
        RECT 1478.080 144.540 1478.340 144.800 ;
        RECT 648.240 75.520 648.500 75.780 ;
        RECT 1477.620 75.520 1477.880 75.780 ;
      LAYER met2 ;
        RECT 1480.300 1700.410 1480.580 1702.400 ;
        RECT 1479.060 1700.270 1480.580 1700.410 ;
        RECT 1479.060 1690.470 1479.200 1700.270 ;
        RECT 1480.300 1700.000 1480.580 1700.270 ;
        RECT 1479.000 1690.150 1479.260 1690.470 ;
        RECT 1478.080 1642.210 1478.340 1642.530 ;
        RECT 1478.140 1559.650 1478.280 1642.210 ;
        RECT 1477.680 1559.510 1478.280 1559.650 ;
        RECT 1477.680 1515.450 1477.820 1559.510 ;
        RECT 1477.680 1515.310 1478.740 1515.450 ;
        RECT 1478.600 1490.550 1478.740 1515.310 ;
        RECT 1478.540 1490.230 1478.800 1490.550 ;
        RECT 1478.540 1466.090 1478.800 1466.410 ;
        RECT 1478.600 1400.790 1478.740 1466.090 ;
        RECT 1477.160 1400.470 1477.420 1400.790 ;
        RECT 1478.540 1400.470 1478.800 1400.790 ;
        RECT 1477.220 1393.650 1477.360 1400.470 ;
        RECT 1477.160 1393.330 1477.420 1393.650 ;
        RECT 1478.080 1345.390 1478.340 1345.710 ;
        RECT 1478.140 1304.230 1478.280 1345.390 ;
        RECT 1477.160 1303.910 1477.420 1304.230 ;
        RECT 1478.080 1303.910 1478.340 1304.230 ;
        RECT 1477.220 1297.090 1477.360 1303.910 ;
        RECT 1477.160 1296.770 1477.420 1297.090 ;
        RECT 1477.620 1200.210 1477.880 1200.530 ;
        RECT 1477.680 1186.930 1477.820 1200.210 ;
        RECT 1477.620 1186.610 1477.880 1186.930 ;
        RECT 1477.620 1138.670 1477.880 1138.990 ;
        RECT 1477.680 1125.050 1477.820 1138.670 ;
        RECT 1477.620 1124.730 1477.880 1125.050 ;
        RECT 1478.080 1124.050 1478.340 1124.370 ;
        RECT 1478.140 1077.110 1478.280 1124.050 ;
        RECT 1478.080 1076.790 1478.340 1077.110 ;
        RECT 1477.160 1055.370 1477.420 1055.690 ;
        RECT 1477.220 1031.550 1477.360 1055.370 ;
        RECT 1477.160 1031.230 1477.420 1031.550 ;
        RECT 1478.540 1031.230 1478.800 1031.550 ;
        RECT 1478.600 1000.610 1478.740 1031.230 ;
        RECT 1477.160 1000.290 1477.420 1000.610 ;
        RECT 1478.540 1000.290 1478.800 1000.610 ;
        RECT 1477.220 952.525 1477.360 1000.290 ;
        RECT 1477.150 952.155 1477.430 952.525 ;
        RECT 1478.070 952.155 1478.350 952.525 ;
        RECT 1478.140 942.470 1478.280 952.155 ;
        RECT 1478.080 942.150 1478.340 942.470 ;
        RECT 1478.080 917.670 1478.340 917.990 ;
        RECT 1478.140 879.650 1478.280 917.670 ;
        RECT 1477.680 879.510 1478.280 879.650 ;
        RECT 1477.680 855.430 1477.820 879.510 ;
        RECT 1477.620 855.110 1477.880 855.430 ;
        RECT 1477.620 807.170 1477.880 807.490 ;
        RECT 1477.680 776.970 1477.820 807.170 ;
        RECT 1477.680 776.830 1478.280 776.970 ;
        RECT 1478.140 759.210 1478.280 776.830 ;
        RECT 1478.080 758.890 1478.340 759.210 ;
        RECT 1478.540 758.210 1478.800 758.530 ;
        RECT 1478.600 752.070 1478.740 758.210 ;
        RECT 1478.540 751.750 1478.800 752.070 ;
        RECT 1478.080 703.810 1478.340 704.130 ;
        RECT 1478.140 703.530 1478.280 703.810 ;
        RECT 1478.140 703.390 1478.740 703.530 ;
        RECT 1478.600 656.725 1478.740 703.390 ;
        RECT 1478.530 656.355 1478.810 656.725 ;
        RECT 1477.610 655.675 1477.890 656.045 ;
        RECT 1477.680 655.510 1477.820 655.675 ;
        RECT 1477.620 655.190 1477.880 655.510 ;
        RECT 1478.080 607.250 1478.340 607.570 ;
        RECT 1478.140 593.970 1478.280 607.250 ;
        RECT 1478.080 593.650 1478.340 593.970 ;
        RECT 1478.080 592.970 1478.340 593.290 ;
        RECT 1478.140 558.950 1478.280 592.970 ;
        RECT 1478.080 558.630 1478.340 558.950 ;
        RECT 1478.540 510.690 1478.800 511.010 ;
        RECT 1478.600 400.850 1478.740 510.690 ;
        RECT 1477.620 400.530 1477.880 400.850 ;
        RECT 1478.540 400.530 1478.800 400.850 ;
        RECT 1477.680 332.930 1477.820 400.530 ;
        RECT 1477.680 332.790 1478.280 332.930 ;
        RECT 1478.140 331.570 1478.280 332.790 ;
        RECT 1477.680 331.430 1478.280 331.570 ;
        RECT 1477.680 290.010 1477.820 331.430 ;
        RECT 1477.620 289.690 1477.880 290.010 ;
        RECT 1478.080 289.010 1478.340 289.330 ;
        RECT 1478.140 241.390 1478.280 289.010 ;
        RECT 1478.080 241.070 1478.340 241.390 ;
        RECT 1478.540 241.070 1478.800 241.390 ;
        RECT 1478.600 191.750 1478.740 241.070 ;
        RECT 1478.540 191.430 1478.800 191.750 ;
        RECT 1478.540 190.750 1478.800 191.070 ;
        RECT 1478.600 145.250 1478.740 190.750 ;
        RECT 1478.140 145.110 1478.740 145.250 ;
        RECT 1478.140 144.830 1478.280 145.110 ;
        RECT 1477.620 144.510 1477.880 144.830 ;
        RECT 1478.080 144.510 1478.340 144.830 ;
        RECT 1477.680 75.810 1477.820 144.510 ;
        RECT 648.240 75.490 648.500 75.810 ;
        RECT 1477.620 75.490 1477.880 75.810 ;
        RECT 648.300 17.410 648.440 75.490 ;
        RECT 645.080 17.270 648.440 17.410 ;
        RECT 645.080 2.400 645.220 17.270 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 1477.150 952.200 1477.430 952.480 ;
        RECT 1478.070 952.200 1478.350 952.480 ;
        RECT 1478.530 656.400 1478.810 656.680 ;
        RECT 1477.610 655.720 1477.890 656.000 ;
      LAYER met3 ;
        RECT 1477.125 952.490 1477.455 952.505 ;
        RECT 1478.045 952.490 1478.375 952.505 ;
        RECT 1477.125 952.190 1478.375 952.490 ;
        RECT 1477.125 952.175 1477.455 952.190 ;
        RECT 1478.045 952.175 1478.375 952.190 ;
        RECT 1478.505 656.690 1478.835 656.705 ;
        RECT 1476.910 656.390 1478.835 656.690 ;
        RECT 1476.910 656.010 1477.210 656.390 ;
        RECT 1478.505 656.375 1478.835 656.390 ;
        RECT 1477.585 656.010 1477.915 656.025 ;
        RECT 1476.910 655.710 1477.915 656.010 ;
        RECT 1477.585 655.695 1477.915 655.710 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2398.970 1687.660 2399.290 1687.720 ;
        RECT 2398.970 1687.520 2404.720 1687.660 ;
        RECT 2398.970 1687.460 2399.290 1687.520 ;
        RECT 2404.580 1686.640 2404.720 1687.520 ;
        RECT 2429.790 1686.640 2430.110 1686.700 ;
        RECT 2404.580 1686.500 2430.110 1686.640 ;
        RECT 2429.790 1686.440 2430.110 1686.500 ;
      LAYER via ;
        RECT 2399.000 1687.460 2399.260 1687.720 ;
        RECT 2429.820 1686.440 2430.080 1686.700 ;
      LAYER met2 ;
        RECT 2398.920 1700.000 2399.200 1702.400 ;
        RECT 2399.060 1687.750 2399.200 1700.000 ;
        RECT 2399.000 1687.430 2399.260 1687.750 ;
        RECT 2429.820 1686.410 2430.080 1686.730 ;
        RECT 2429.880 3.130 2430.020 1686.410 ;
        RECT 2428.960 2.990 2430.020 3.130 ;
        RECT 2428.960 2.400 2429.100 2.990 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2408.170 1687.660 2408.490 1687.720 ;
        RECT 2414.150 1687.660 2414.470 1687.720 ;
        RECT 2408.170 1687.520 2414.470 1687.660 ;
        RECT 2408.170 1687.460 2408.490 1687.520 ;
        RECT 2414.150 1687.460 2414.470 1687.520 ;
        RECT 2414.150 16.900 2414.470 16.960 ;
        RECT 2446.810 16.900 2447.130 16.960 ;
        RECT 2414.150 16.760 2447.130 16.900 ;
        RECT 2414.150 16.700 2414.470 16.760 ;
        RECT 2446.810 16.700 2447.130 16.760 ;
      LAYER via ;
        RECT 2408.200 1687.460 2408.460 1687.720 ;
        RECT 2414.180 1687.460 2414.440 1687.720 ;
        RECT 2414.180 16.700 2414.440 16.960 ;
        RECT 2446.840 16.700 2447.100 16.960 ;
      LAYER met2 ;
        RECT 2408.120 1700.000 2408.400 1702.400 ;
        RECT 2408.260 1687.750 2408.400 1700.000 ;
        RECT 2408.200 1687.430 2408.460 1687.750 ;
        RECT 2414.180 1687.430 2414.440 1687.750 ;
        RECT 2414.240 16.990 2414.380 1687.430 ;
        RECT 2414.180 16.670 2414.440 16.990 ;
        RECT 2446.840 16.670 2447.100 16.990 ;
        RECT 2446.900 2.400 2447.040 16.670 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2417.370 1688.340 2417.690 1688.400 ;
        RECT 2421.050 1688.340 2421.370 1688.400 ;
        RECT 2417.370 1688.200 2421.370 1688.340 ;
        RECT 2417.370 1688.140 2417.690 1688.200 ;
        RECT 2421.050 1688.140 2421.370 1688.200 ;
        RECT 2421.050 18.260 2421.370 18.320 ;
        RECT 2464.750 18.260 2465.070 18.320 ;
        RECT 2421.050 18.120 2465.070 18.260 ;
        RECT 2421.050 18.060 2421.370 18.120 ;
        RECT 2464.750 18.060 2465.070 18.120 ;
      LAYER via ;
        RECT 2417.400 1688.140 2417.660 1688.400 ;
        RECT 2421.080 1688.140 2421.340 1688.400 ;
        RECT 2421.080 18.060 2421.340 18.320 ;
        RECT 2464.780 18.060 2465.040 18.320 ;
      LAYER met2 ;
        RECT 2417.320 1700.000 2417.600 1702.400 ;
        RECT 2417.460 1688.430 2417.600 1700.000 ;
        RECT 2417.400 1688.110 2417.660 1688.430 ;
        RECT 2421.080 1688.110 2421.340 1688.430 ;
        RECT 2421.140 18.350 2421.280 1688.110 ;
        RECT 2421.080 18.030 2421.340 18.350 ;
        RECT 2464.780 18.030 2465.040 18.350 ;
        RECT 2464.840 2.400 2464.980 18.030 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2426.570 1687.320 2426.890 1687.380 ;
        RECT 2466.590 1687.320 2466.910 1687.380 ;
        RECT 2426.570 1687.180 2466.910 1687.320 ;
        RECT 2426.570 1687.120 2426.890 1687.180 ;
        RECT 2466.590 1687.120 2466.910 1687.180 ;
        RECT 2466.590 15.880 2466.910 15.940 ;
        RECT 2482.690 15.880 2483.010 15.940 ;
        RECT 2466.590 15.740 2483.010 15.880 ;
        RECT 2466.590 15.680 2466.910 15.740 ;
        RECT 2482.690 15.680 2483.010 15.740 ;
      LAYER via ;
        RECT 2426.600 1687.120 2426.860 1687.380 ;
        RECT 2466.620 1687.120 2466.880 1687.380 ;
        RECT 2466.620 15.680 2466.880 15.940 ;
        RECT 2482.720 15.680 2482.980 15.940 ;
      LAYER met2 ;
        RECT 2426.520 1700.000 2426.800 1702.400 ;
        RECT 2426.660 1687.410 2426.800 1700.000 ;
        RECT 2426.600 1687.090 2426.860 1687.410 ;
        RECT 2466.620 1687.090 2466.880 1687.410 ;
        RECT 2466.680 15.970 2466.820 1687.090 ;
        RECT 2466.620 15.650 2466.880 15.970 ;
        RECT 2482.720 15.650 2482.980 15.970 ;
        RECT 2482.780 2.400 2482.920 15.650 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2435.770 1689.360 2436.090 1689.420 ;
        RECT 2498.790 1689.360 2499.110 1689.420 ;
        RECT 2435.770 1689.220 2499.110 1689.360 ;
        RECT 2435.770 1689.160 2436.090 1689.220 ;
        RECT 2498.790 1689.160 2499.110 1689.220 ;
        RECT 2498.790 2.960 2499.110 3.020 ;
        RECT 2500.630 2.960 2500.950 3.020 ;
        RECT 2498.790 2.820 2500.950 2.960 ;
        RECT 2498.790 2.760 2499.110 2.820 ;
        RECT 2500.630 2.760 2500.950 2.820 ;
      LAYER via ;
        RECT 2435.800 1689.160 2436.060 1689.420 ;
        RECT 2498.820 1689.160 2499.080 1689.420 ;
        RECT 2498.820 2.760 2499.080 3.020 ;
        RECT 2500.660 2.760 2500.920 3.020 ;
      LAYER met2 ;
        RECT 2435.720 1700.000 2436.000 1702.400 ;
        RECT 2435.860 1689.450 2436.000 1700.000 ;
        RECT 2435.800 1689.130 2436.060 1689.450 ;
        RECT 2498.820 1689.130 2499.080 1689.450 ;
        RECT 2498.880 3.050 2499.020 1689.130 ;
        RECT 2498.820 2.730 2499.080 3.050 ;
        RECT 2500.660 2.730 2500.920 3.050 ;
        RECT 2500.720 2.400 2500.860 2.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2444.970 1688.680 2445.290 1688.740 ;
        RECT 2513.050 1688.680 2513.370 1688.740 ;
        RECT 2444.970 1688.540 2499.480 1688.680 ;
        RECT 2444.970 1688.480 2445.290 1688.540 ;
        RECT 2499.340 1688.340 2499.480 1688.540 ;
        RECT 2504.400 1688.540 2513.370 1688.680 ;
        RECT 2504.400 1688.340 2504.540 1688.540 ;
        RECT 2513.050 1688.480 2513.370 1688.540 ;
        RECT 2499.340 1688.200 2504.540 1688.340 ;
      LAYER via ;
        RECT 2445.000 1688.480 2445.260 1688.740 ;
        RECT 2513.080 1688.480 2513.340 1688.740 ;
      LAYER met2 ;
        RECT 2444.920 1700.000 2445.200 1702.400 ;
        RECT 2445.060 1688.770 2445.200 1700.000 ;
        RECT 2445.000 1688.450 2445.260 1688.770 ;
        RECT 2513.080 1688.450 2513.340 1688.770 ;
        RECT 2513.140 16.050 2513.280 1688.450 ;
        RECT 2513.140 15.910 2518.340 16.050 ;
        RECT 2518.200 2.400 2518.340 15.910 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2494.725 1688.185 2494.895 1690.395 ;
        RECT 2498.865 1686.485 2499.035 1688.355 ;
      LAYER mcon ;
        RECT 2494.725 1690.225 2494.895 1690.395 ;
        RECT 2498.865 1688.185 2499.035 1688.355 ;
      LAYER met1 ;
        RECT 2454.170 1690.380 2454.490 1690.440 ;
        RECT 2494.665 1690.380 2494.955 1690.425 ;
        RECT 2454.170 1690.240 2494.955 1690.380 ;
        RECT 2454.170 1690.180 2454.490 1690.240 ;
        RECT 2494.665 1690.195 2494.955 1690.240 ;
        RECT 2494.665 1688.340 2494.955 1688.385 ;
        RECT 2498.805 1688.340 2499.095 1688.385 ;
        RECT 2494.665 1688.200 2499.095 1688.340 ;
        RECT 2494.665 1688.155 2494.955 1688.200 ;
        RECT 2498.805 1688.155 2499.095 1688.200 ;
        RECT 2498.805 1686.640 2499.095 1686.685 ;
        RECT 2533.290 1686.640 2533.610 1686.700 ;
        RECT 2498.805 1686.500 2533.610 1686.640 ;
        RECT 2498.805 1686.455 2499.095 1686.500 ;
        RECT 2533.290 1686.440 2533.610 1686.500 ;
        RECT 2533.290 2.960 2533.610 3.020 ;
        RECT 2536.050 2.960 2536.370 3.020 ;
        RECT 2533.290 2.820 2536.370 2.960 ;
        RECT 2533.290 2.760 2533.610 2.820 ;
        RECT 2536.050 2.760 2536.370 2.820 ;
      LAYER via ;
        RECT 2454.200 1690.180 2454.460 1690.440 ;
        RECT 2533.320 1686.440 2533.580 1686.700 ;
        RECT 2533.320 2.760 2533.580 3.020 ;
        RECT 2536.080 2.760 2536.340 3.020 ;
      LAYER met2 ;
        RECT 2454.120 1700.000 2454.400 1702.400 ;
        RECT 2454.260 1690.470 2454.400 1700.000 ;
        RECT 2454.200 1690.150 2454.460 1690.470 ;
        RECT 2533.320 1686.410 2533.580 1686.730 ;
        RECT 2533.380 3.050 2533.520 1686.410 ;
        RECT 2533.320 2.730 2533.580 3.050 ;
        RECT 2536.080 2.730 2536.340 3.050 ;
        RECT 2536.140 2.400 2536.280 2.730 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2478.180 1688.200 2484.300 1688.340 ;
        RECT 2463.370 1688.000 2463.690 1688.060 ;
        RECT 2478.180 1688.000 2478.320 1688.200 ;
        RECT 2463.370 1687.860 2478.320 1688.000 ;
        RECT 2484.160 1688.000 2484.300 1688.200 ;
        RECT 2553.990 1688.000 2554.310 1688.060 ;
        RECT 2484.160 1687.860 2554.310 1688.000 ;
        RECT 2463.370 1687.800 2463.690 1687.860 ;
        RECT 2553.990 1687.800 2554.310 1687.860 ;
      LAYER via ;
        RECT 2463.400 1687.800 2463.660 1688.060 ;
        RECT 2554.020 1687.800 2554.280 1688.060 ;
      LAYER met2 ;
        RECT 2463.320 1700.000 2463.600 1702.400 ;
        RECT 2463.460 1688.090 2463.600 1700.000 ;
        RECT 2463.400 1687.770 2463.660 1688.090 ;
        RECT 2554.020 1687.770 2554.280 1688.090 ;
        RECT 2554.080 2.400 2554.220 1687.770 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2472.570 1687.660 2472.890 1687.720 ;
        RECT 2567.790 1687.660 2568.110 1687.720 ;
        RECT 2472.570 1687.520 2568.110 1687.660 ;
        RECT 2472.570 1687.460 2472.890 1687.520 ;
        RECT 2567.790 1687.460 2568.110 1687.520 ;
        RECT 2567.790 2.960 2568.110 3.020 ;
        RECT 2571.930 2.960 2572.250 3.020 ;
        RECT 2567.790 2.820 2572.250 2.960 ;
        RECT 2567.790 2.760 2568.110 2.820 ;
        RECT 2571.930 2.760 2572.250 2.820 ;
      LAYER via ;
        RECT 2472.600 1687.460 2472.860 1687.720 ;
        RECT 2567.820 1687.460 2568.080 1687.720 ;
        RECT 2567.820 2.760 2568.080 3.020 ;
        RECT 2571.960 2.760 2572.220 3.020 ;
      LAYER met2 ;
        RECT 2472.520 1700.000 2472.800 1702.400 ;
        RECT 2472.660 1687.750 2472.800 1700.000 ;
        RECT 2472.600 1687.430 2472.860 1687.750 ;
        RECT 2567.820 1687.430 2568.080 1687.750 ;
        RECT 2567.880 3.050 2568.020 1687.430 ;
        RECT 2567.820 2.730 2568.080 3.050 ;
        RECT 2571.960 2.730 2572.220 3.050 ;
        RECT 2572.020 2.400 2572.160 2.730 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2481.310 1687.320 2481.630 1687.380 ;
        RECT 2588.030 1687.320 2588.350 1687.380 ;
        RECT 2481.310 1687.180 2588.350 1687.320 ;
        RECT 2481.310 1687.120 2481.630 1687.180 ;
        RECT 2588.030 1687.120 2588.350 1687.180 ;
      LAYER via ;
        RECT 2481.340 1687.120 2481.600 1687.380 ;
        RECT 2588.060 1687.120 2588.320 1687.380 ;
      LAYER met2 ;
        RECT 2481.260 1700.000 2481.540 1702.400 ;
        RECT 2481.400 1687.410 2481.540 1700.000 ;
        RECT 2481.340 1687.090 2481.600 1687.410 ;
        RECT 2588.060 1687.090 2588.320 1687.410 ;
        RECT 2588.120 3.130 2588.260 1687.090 ;
        RECT 2588.120 2.990 2589.640 3.130 ;
        RECT 2589.500 2.400 2589.640 2.990 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1567.290 1689.360 1567.610 1689.420 ;
        RECT 1570.510 1689.360 1570.830 1689.420 ;
        RECT 1567.290 1689.220 1570.830 1689.360 ;
        RECT 1567.290 1689.160 1567.610 1689.220 ;
        RECT 1570.510 1689.160 1570.830 1689.220 ;
        RECT 827.610 71.300 827.930 71.360 ;
        RECT 1567.290 71.300 1567.610 71.360 ;
        RECT 827.610 71.160 1567.610 71.300 ;
        RECT 827.610 71.100 827.930 71.160 ;
        RECT 1567.290 71.100 1567.610 71.160 ;
      LAYER via ;
        RECT 1567.320 1689.160 1567.580 1689.420 ;
        RECT 1570.540 1689.160 1570.800 1689.420 ;
        RECT 827.640 71.100 827.900 71.360 ;
        RECT 1567.320 71.100 1567.580 71.360 ;
      LAYER met2 ;
        RECT 1572.300 1700.410 1572.580 1702.400 ;
        RECT 1570.600 1700.270 1572.580 1700.410 ;
        RECT 1570.600 1689.450 1570.740 1700.270 ;
        RECT 1572.300 1700.000 1572.580 1700.270 ;
        RECT 1567.320 1689.130 1567.580 1689.450 ;
        RECT 1570.540 1689.130 1570.800 1689.450 ;
        RECT 1567.380 71.390 1567.520 1689.130 ;
        RECT 827.640 71.070 827.900 71.390 ;
        RECT 1567.320 71.070 1567.580 71.390 ;
        RECT 827.700 16.730 827.840 71.070 ;
        RECT 823.560 16.590 827.840 16.730 ;
        RECT 823.560 2.400 823.700 16.590 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2490.510 1686.980 2490.830 1687.040 ;
        RECT 2601.830 1686.980 2602.150 1687.040 ;
        RECT 2490.510 1686.840 2602.150 1686.980 ;
        RECT 2490.510 1686.780 2490.830 1686.840 ;
        RECT 2601.830 1686.780 2602.150 1686.840 ;
        RECT 2601.830 2.960 2602.150 3.020 ;
        RECT 2607.350 2.960 2607.670 3.020 ;
        RECT 2601.830 2.820 2607.670 2.960 ;
        RECT 2601.830 2.760 2602.150 2.820 ;
        RECT 2607.350 2.760 2607.670 2.820 ;
      LAYER via ;
        RECT 2490.540 1686.780 2490.800 1687.040 ;
        RECT 2601.860 1686.780 2602.120 1687.040 ;
        RECT 2601.860 2.760 2602.120 3.020 ;
        RECT 2607.380 2.760 2607.640 3.020 ;
      LAYER met2 ;
        RECT 2490.460 1700.000 2490.740 1702.400 ;
        RECT 2490.600 1687.070 2490.740 1700.000 ;
        RECT 2490.540 1686.750 2490.800 1687.070 ;
        RECT 2601.860 1686.750 2602.120 1687.070 ;
        RECT 2601.920 3.050 2602.060 1686.750 ;
        RECT 2601.860 2.730 2602.120 3.050 ;
        RECT 2607.380 2.730 2607.640 3.050 ;
        RECT 2607.440 2.400 2607.580 2.730 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2615.245 18.105 2615.415 19.295 ;
      LAYER mcon ;
        RECT 2615.245 19.125 2615.415 19.295 ;
      LAYER met1 ;
        RECT 2499.710 1688.680 2500.030 1688.740 ;
        RECT 2503.850 1688.680 2504.170 1688.740 ;
        RECT 2499.710 1688.540 2504.170 1688.680 ;
        RECT 2499.710 1688.480 2500.030 1688.540 ;
        RECT 2503.850 1688.480 2504.170 1688.540 ;
        RECT 2615.185 19.280 2615.475 19.325 ;
        RECT 2625.290 19.280 2625.610 19.340 ;
        RECT 2615.185 19.140 2625.610 19.280 ;
        RECT 2615.185 19.095 2615.475 19.140 ;
        RECT 2625.290 19.080 2625.610 19.140 ;
        RECT 2503.850 18.260 2504.170 18.320 ;
        RECT 2615.185 18.260 2615.475 18.305 ;
        RECT 2503.850 18.120 2615.475 18.260 ;
        RECT 2503.850 18.060 2504.170 18.120 ;
        RECT 2615.185 18.075 2615.475 18.120 ;
      LAYER via ;
        RECT 2499.740 1688.480 2500.000 1688.740 ;
        RECT 2503.880 1688.480 2504.140 1688.740 ;
        RECT 2625.320 19.080 2625.580 19.340 ;
        RECT 2503.880 18.060 2504.140 18.320 ;
      LAYER met2 ;
        RECT 2499.660 1700.000 2499.940 1702.400 ;
        RECT 2499.800 1688.770 2499.940 1700.000 ;
        RECT 2499.740 1688.450 2500.000 1688.770 ;
        RECT 2503.880 1688.450 2504.140 1688.770 ;
        RECT 2503.940 18.350 2504.080 1688.450 ;
        RECT 2625.320 19.050 2625.580 19.370 ;
        RECT 2503.880 18.030 2504.140 18.350 ;
        RECT 2625.380 2.400 2625.520 19.050 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2511.210 17.240 2511.530 17.300 ;
        RECT 2643.230 17.240 2643.550 17.300 ;
        RECT 2511.210 17.100 2643.550 17.240 ;
        RECT 2511.210 17.040 2511.530 17.100 ;
        RECT 2643.230 17.040 2643.550 17.100 ;
      LAYER via ;
        RECT 2511.240 17.040 2511.500 17.300 ;
        RECT 2643.260 17.040 2643.520 17.300 ;
      LAYER met2 ;
        RECT 2508.860 1700.410 2509.140 1702.400 ;
        RECT 2508.860 1700.270 2511.440 1700.410 ;
        RECT 2508.860 1700.000 2509.140 1700.270 ;
        RECT 2511.300 17.330 2511.440 1700.270 ;
        RECT 2511.240 17.010 2511.500 17.330 ;
        RECT 2643.260 17.010 2643.520 17.330 ;
        RECT 2643.320 2.400 2643.460 17.010 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2570.165 1683.765 2570.335 1684.955 ;
      LAYER mcon ;
        RECT 2570.165 1684.785 2570.335 1684.955 ;
      LAYER met1 ;
        RECT 2517.190 1689.700 2517.510 1689.760 ;
        RECT 2518.110 1689.700 2518.430 1689.760 ;
        RECT 2517.190 1689.560 2518.430 1689.700 ;
        RECT 2517.190 1689.500 2517.510 1689.560 ;
        RECT 2518.110 1689.500 2518.430 1689.560 ;
        RECT 2517.190 1684.940 2517.510 1685.000 ;
        RECT 2570.105 1684.940 2570.395 1684.985 ;
        RECT 2517.190 1684.800 2570.395 1684.940 ;
        RECT 2517.190 1684.740 2517.510 1684.800 ;
        RECT 2570.105 1684.755 2570.395 1684.800 ;
        RECT 2570.105 1683.920 2570.395 1683.965 ;
        RECT 2656.570 1683.920 2656.890 1683.980 ;
        RECT 2570.105 1683.780 2622.300 1683.920 ;
        RECT 2570.105 1683.735 2570.395 1683.780 ;
        RECT 2622.160 1683.580 2622.300 1683.780 ;
        RECT 2628.600 1683.780 2637.480 1683.920 ;
        RECT 2628.600 1683.580 2628.740 1683.780 ;
        RECT 2622.160 1683.440 2628.740 1683.580 ;
        RECT 2637.340 1683.580 2637.480 1683.780 ;
        RECT 2642.860 1683.780 2646.680 1683.920 ;
        RECT 2642.860 1683.580 2643.000 1683.780 ;
        RECT 2637.340 1683.440 2643.000 1683.580 ;
        RECT 2646.540 1683.580 2646.680 1683.780 ;
        RECT 2649.760 1683.780 2656.890 1683.920 ;
        RECT 2649.760 1683.580 2649.900 1683.780 ;
        RECT 2656.570 1683.720 2656.890 1683.780 ;
        RECT 2646.540 1683.440 2649.900 1683.580 ;
      LAYER via ;
        RECT 2517.220 1689.500 2517.480 1689.760 ;
        RECT 2518.140 1689.500 2518.400 1689.760 ;
        RECT 2517.220 1684.740 2517.480 1685.000 ;
        RECT 2656.600 1683.720 2656.860 1683.980 ;
      LAYER met2 ;
        RECT 2518.060 1700.000 2518.340 1702.400 ;
        RECT 2518.200 1689.790 2518.340 1700.000 ;
        RECT 2517.220 1689.470 2517.480 1689.790 ;
        RECT 2518.140 1689.470 2518.400 1689.790 ;
        RECT 2517.280 1685.030 2517.420 1689.470 ;
        RECT 2517.220 1684.710 2517.480 1685.030 ;
        RECT 2656.600 1683.690 2656.860 1684.010 ;
        RECT 2656.660 16.730 2656.800 1683.690 ;
        RECT 2656.660 16.590 2661.400 16.730 ;
        RECT 2661.260 2.400 2661.400 16.590 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2527.310 1688.680 2527.630 1688.740 ;
        RECT 2531.910 1688.680 2532.230 1688.740 ;
        RECT 2527.310 1688.540 2532.230 1688.680 ;
        RECT 2527.310 1688.480 2527.630 1688.540 ;
        RECT 2531.910 1688.480 2532.230 1688.540 ;
        RECT 2531.910 14.860 2532.230 14.920 ;
        RECT 2678.650 14.860 2678.970 14.920 ;
        RECT 2531.910 14.720 2678.970 14.860 ;
        RECT 2531.910 14.660 2532.230 14.720 ;
        RECT 2678.650 14.660 2678.970 14.720 ;
      LAYER via ;
        RECT 2527.340 1688.480 2527.600 1688.740 ;
        RECT 2531.940 1688.480 2532.200 1688.740 ;
        RECT 2531.940 14.660 2532.200 14.920 ;
        RECT 2678.680 14.660 2678.940 14.920 ;
      LAYER met2 ;
        RECT 2527.260 1700.000 2527.540 1702.400 ;
        RECT 2527.400 1688.770 2527.540 1700.000 ;
        RECT 2527.340 1688.450 2527.600 1688.770 ;
        RECT 2531.940 1688.450 2532.200 1688.770 ;
        RECT 2532.000 14.950 2532.140 1688.450 ;
        RECT 2531.940 14.630 2532.200 14.950 ;
        RECT 2678.680 14.630 2678.940 14.950 ;
        RECT 2678.740 2.400 2678.880 14.630 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2536.510 1685.620 2536.830 1685.680 ;
        RECT 2691.070 1685.620 2691.390 1685.680 ;
        RECT 2536.510 1685.480 2691.390 1685.620 ;
        RECT 2536.510 1685.420 2536.830 1685.480 ;
        RECT 2691.070 1685.420 2691.390 1685.480 ;
      LAYER via ;
        RECT 2536.540 1685.420 2536.800 1685.680 ;
        RECT 2691.100 1685.420 2691.360 1685.680 ;
      LAYER met2 ;
        RECT 2536.460 1700.000 2536.740 1702.400 ;
        RECT 2536.600 1685.710 2536.740 1700.000 ;
        RECT 2536.540 1685.390 2536.800 1685.710 ;
        RECT 2691.100 1685.390 2691.360 1685.710 ;
        RECT 2691.160 16.730 2691.300 1685.390 ;
        RECT 2691.160 16.590 2696.820 16.730 ;
        RECT 2696.680 2.400 2696.820 16.590 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2545.710 1690.380 2546.030 1690.440 ;
        RECT 2711.770 1690.380 2712.090 1690.440 ;
        RECT 2545.710 1690.240 2712.090 1690.380 ;
        RECT 2545.710 1690.180 2546.030 1690.240 ;
        RECT 2711.770 1690.180 2712.090 1690.240 ;
      LAYER via ;
        RECT 2545.740 1690.180 2546.000 1690.440 ;
        RECT 2711.800 1690.180 2712.060 1690.440 ;
      LAYER met2 ;
        RECT 2545.660 1700.000 2545.940 1702.400 ;
        RECT 2545.800 1690.470 2545.940 1700.000 ;
        RECT 2545.740 1690.150 2546.000 1690.470 ;
        RECT 2711.800 1690.150 2712.060 1690.470 ;
        RECT 2711.860 16.730 2712.000 1690.150 ;
        RECT 2711.860 16.590 2714.760 16.730 ;
        RECT 2714.620 2.400 2714.760 16.590 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2554.910 1688.680 2555.230 1688.740 ;
        RECT 2559.510 1688.680 2559.830 1688.740 ;
        RECT 2554.910 1688.540 2559.830 1688.680 ;
        RECT 2554.910 1688.480 2555.230 1688.540 ;
        RECT 2559.510 1688.480 2559.830 1688.540 ;
        RECT 2559.510 15.540 2559.830 15.600 ;
        RECT 2559.510 15.400 2695.440 15.540 ;
        RECT 2559.510 15.340 2559.830 15.400 ;
        RECT 2695.300 15.200 2695.440 15.400 ;
        RECT 2732.470 15.200 2732.790 15.260 ;
        RECT 2695.300 15.060 2732.790 15.200 ;
        RECT 2732.470 15.000 2732.790 15.060 ;
      LAYER via ;
        RECT 2554.940 1688.480 2555.200 1688.740 ;
        RECT 2559.540 1688.480 2559.800 1688.740 ;
        RECT 2559.540 15.340 2559.800 15.600 ;
        RECT 2732.500 15.000 2732.760 15.260 ;
      LAYER met2 ;
        RECT 2554.860 1700.000 2555.140 1702.400 ;
        RECT 2555.000 1688.770 2555.140 1700.000 ;
        RECT 2554.940 1688.450 2555.200 1688.770 ;
        RECT 2559.540 1688.450 2559.800 1688.770 ;
        RECT 2559.600 15.630 2559.740 1688.450 ;
        RECT 2559.540 15.310 2559.800 15.630 ;
        RECT 2732.500 14.970 2732.760 15.290 ;
        RECT 2732.560 2.400 2732.700 14.970 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2564.110 1690.040 2564.430 1690.100 ;
        RECT 2735.690 1690.040 2736.010 1690.100 ;
        RECT 2564.110 1689.900 2736.010 1690.040 ;
        RECT 2564.110 1689.840 2564.430 1689.900 ;
        RECT 2735.690 1689.840 2736.010 1689.900 ;
        RECT 2735.690 16.220 2736.010 16.280 ;
        RECT 2750.410 16.220 2750.730 16.280 ;
        RECT 2735.690 16.080 2750.730 16.220 ;
        RECT 2735.690 16.020 2736.010 16.080 ;
        RECT 2750.410 16.020 2750.730 16.080 ;
      LAYER via ;
        RECT 2564.140 1689.840 2564.400 1690.100 ;
        RECT 2735.720 1689.840 2735.980 1690.100 ;
        RECT 2735.720 16.020 2735.980 16.280 ;
        RECT 2750.440 16.020 2750.700 16.280 ;
      LAYER met2 ;
        RECT 2564.060 1700.000 2564.340 1702.400 ;
        RECT 2564.200 1690.130 2564.340 1700.000 ;
        RECT 2564.140 1689.810 2564.400 1690.130 ;
        RECT 2735.720 1689.810 2735.980 1690.130 ;
        RECT 2735.780 16.310 2735.920 1689.810 ;
        RECT 2735.720 15.990 2735.980 16.310 ;
        RECT 2750.440 15.990 2750.700 16.310 ;
        RECT 2750.500 2.400 2750.640 15.990 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2573.310 1689.360 2573.630 1689.420 ;
        RECT 2573.310 1689.220 2593.780 1689.360 ;
        RECT 2573.310 1689.160 2573.630 1689.220 ;
        RECT 2593.640 1689.020 2593.780 1689.220 ;
        RECT 2766.970 1689.020 2767.290 1689.080 ;
        RECT 2593.640 1688.880 2767.290 1689.020 ;
        RECT 2766.970 1688.820 2767.290 1688.880 ;
      LAYER via ;
        RECT 2573.340 1689.160 2573.600 1689.420 ;
        RECT 2767.000 1688.820 2767.260 1689.080 ;
      LAYER met2 ;
        RECT 2573.260 1700.000 2573.540 1702.400 ;
        RECT 2573.400 1689.450 2573.540 1700.000 ;
        RECT 2573.340 1689.130 2573.600 1689.450 ;
        RECT 2767.000 1688.790 2767.260 1689.110 ;
        RECT 2767.060 16.730 2767.200 1688.790 ;
        RECT 2767.060 16.590 2768.120 16.730 ;
        RECT 2767.980 2.400 2768.120 16.590 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 841.410 70.960 841.730 71.020 ;
        RECT 1580.630 70.960 1580.950 71.020 ;
        RECT 841.410 70.820 1580.950 70.960 ;
        RECT 841.410 70.760 841.730 70.820 ;
        RECT 1580.630 70.760 1580.950 70.820 ;
      LAYER via ;
        RECT 841.440 70.760 841.700 71.020 ;
        RECT 1580.660 70.760 1580.920 71.020 ;
      LAYER met2 ;
        RECT 1581.500 1700.410 1581.780 1702.400 ;
        RECT 1580.720 1700.270 1581.780 1700.410 ;
        RECT 1580.720 71.050 1580.860 1700.270 ;
        RECT 1581.500 1700.000 1581.780 1700.270 ;
        RECT 841.440 70.730 841.700 71.050 ;
        RECT 1580.660 70.730 1580.920 71.050 ;
        RECT 841.500 17.410 841.640 70.730 ;
        RECT 841.040 17.270 841.640 17.410 ;
        RECT 841.040 2.400 841.180 17.270 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2582.510 1688.680 2582.830 1688.740 ;
        RECT 2587.110 1688.680 2587.430 1688.740 ;
        RECT 2582.510 1688.540 2587.430 1688.680 ;
        RECT 2582.510 1688.480 2582.830 1688.540 ;
        RECT 2587.110 1688.480 2587.430 1688.540 ;
        RECT 2587.110 16.900 2587.430 16.960 ;
        RECT 2785.830 16.900 2786.150 16.960 ;
        RECT 2587.110 16.760 2786.150 16.900 ;
        RECT 2587.110 16.700 2587.430 16.760 ;
        RECT 2785.830 16.700 2786.150 16.760 ;
      LAYER via ;
        RECT 2582.540 1688.480 2582.800 1688.740 ;
        RECT 2587.140 1688.480 2587.400 1688.740 ;
        RECT 2587.140 16.700 2587.400 16.960 ;
        RECT 2785.860 16.700 2786.120 16.960 ;
      LAYER met2 ;
        RECT 2582.460 1700.000 2582.740 1702.400 ;
        RECT 2582.600 1688.770 2582.740 1700.000 ;
        RECT 2582.540 1688.450 2582.800 1688.770 ;
        RECT 2587.140 1688.450 2587.400 1688.770 ;
        RECT 2587.200 16.990 2587.340 1688.450 ;
        RECT 2587.140 16.670 2587.400 16.990 ;
        RECT 2785.860 16.670 2786.120 16.990 ;
        RECT 2785.920 2.400 2786.060 16.670 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2591.710 1688.340 2592.030 1688.400 ;
        RECT 2801.470 1688.340 2801.790 1688.400 ;
        RECT 2591.710 1688.200 2801.790 1688.340 ;
        RECT 2591.710 1688.140 2592.030 1688.200 ;
        RECT 2801.470 1688.140 2801.790 1688.200 ;
      LAYER via ;
        RECT 2591.740 1688.140 2592.000 1688.400 ;
        RECT 2801.500 1688.140 2801.760 1688.400 ;
      LAYER met2 ;
        RECT 2591.660 1700.000 2591.940 1702.400 ;
        RECT 2591.800 1688.430 2591.940 1700.000 ;
        RECT 2591.740 1688.110 2592.000 1688.430 ;
        RECT 2801.500 1688.110 2801.760 1688.430 ;
        RECT 2801.560 17.410 2801.700 1688.110 ;
        RECT 2801.560 17.270 2804.000 17.410 ;
        RECT 2803.860 2.400 2804.000 17.270 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2600.910 19.960 2601.230 20.020 ;
        RECT 2821.710 19.960 2822.030 20.020 ;
        RECT 2600.910 19.820 2822.030 19.960 ;
        RECT 2600.910 19.760 2601.230 19.820 ;
        RECT 2821.710 19.760 2822.030 19.820 ;
      LAYER via ;
        RECT 2600.940 19.760 2601.200 20.020 ;
        RECT 2821.740 19.760 2822.000 20.020 ;
      LAYER met2 ;
        RECT 2600.860 1700.000 2601.140 1702.400 ;
        RECT 2601.000 20.050 2601.140 1700.000 ;
        RECT 2600.940 19.730 2601.200 20.050 ;
        RECT 2821.740 19.730 2822.000 20.050 ;
        RECT 2821.800 2.400 2821.940 19.730 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2610.110 1688.000 2610.430 1688.060 ;
        RECT 2610.110 1687.860 2633.340 1688.000 ;
        RECT 2610.110 1687.800 2610.430 1687.860 ;
        RECT 2633.200 1687.660 2633.340 1687.860 ;
        RECT 2835.970 1687.660 2836.290 1687.720 ;
        RECT 2633.200 1687.520 2836.290 1687.660 ;
        RECT 2835.970 1687.460 2836.290 1687.520 ;
      LAYER via ;
        RECT 2610.140 1687.800 2610.400 1688.060 ;
        RECT 2836.000 1687.460 2836.260 1687.720 ;
      LAYER met2 ;
        RECT 2610.060 1700.000 2610.340 1702.400 ;
        RECT 2610.200 1688.090 2610.340 1700.000 ;
        RECT 2610.140 1687.770 2610.400 1688.090 ;
        RECT 2836.000 1687.430 2836.260 1687.750 ;
        RECT 2836.060 17.410 2836.200 1687.430 ;
        RECT 2836.060 17.270 2839.420 17.410 ;
        RECT 2839.280 2.400 2839.420 17.270 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2621.610 18.600 2621.930 18.660 ;
        RECT 2857.130 18.600 2857.450 18.660 ;
        RECT 2621.610 18.460 2857.450 18.600 ;
        RECT 2621.610 18.400 2621.930 18.460 ;
        RECT 2857.130 18.400 2857.450 18.460 ;
      LAYER via ;
        RECT 2621.640 18.400 2621.900 18.660 ;
        RECT 2857.160 18.400 2857.420 18.660 ;
      LAYER met2 ;
        RECT 2619.260 1700.410 2619.540 1702.400 ;
        RECT 2619.260 1700.270 2621.840 1700.410 ;
        RECT 2619.260 1700.000 2619.540 1700.270 ;
        RECT 2621.700 18.690 2621.840 1700.270 ;
        RECT 2621.640 18.370 2621.900 18.690 ;
        RECT 2857.160 18.370 2857.420 18.690 ;
        RECT 2857.220 2.400 2857.360 18.370 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2628.460 1700.000 2628.740 1702.400 ;
        RECT 2628.600 16.845 2628.740 1700.000 ;
        RECT 2628.530 16.475 2628.810 16.845 ;
        RECT 2875.090 16.475 2875.370 16.845 ;
        RECT 2875.160 2.400 2875.300 16.475 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 2628.530 16.520 2628.810 16.800 ;
        RECT 2875.090 16.520 2875.370 16.800 ;
      LAYER met3 ;
        RECT 2628.505 16.810 2628.835 16.825 ;
        RECT 2875.065 16.810 2875.395 16.825 ;
        RECT 2628.505 16.510 2875.395 16.810 ;
        RECT 2628.505 16.495 2628.835 16.510 ;
        RECT 2875.065 16.495 2875.395 16.510 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2637.710 1683.920 2638.030 1683.980 ;
        RECT 2642.310 1683.920 2642.630 1683.980 ;
        RECT 2637.710 1683.780 2642.630 1683.920 ;
        RECT 2637.710 1683.720 2638.030 1683.780 ;
        RECT 2642.310 1683.720 2642.630 1683.780 ;
        RECT 2642.310 17.580 2642.630 17.640 ;
        RECT 2893.010 17.580 2893.330 17.640 ;
        RECT 2642.310 17.440 2893.330 17.580 ;
        RECT 2642.310 17.380 2642.630 17.440 ;
        RECT 2893.010 17.380 2893.330 17.440 ;
      LAYER via ;
        RECT 2637.740 1683.720 2638.000 1683.980 ;
        RECT 2642.340 1683.720 2642.600 1683.980 ;
        RECT 2642.340 17.380 2642.600 17.640 ;
        RECT 2893.040 17.380 2893.300 17.640 ;
      LAYER met2 ;
        RECT 2637.660 1700.000 2637.940 1702.400 ;
        RECT 2637.800 1684.010 2637.940 1700.000 ;
        RECT 2637.740 1683.690 2638.000 1684.010 ;
        RECT 2642.340 1683.690 2642.600 1684.010 ;
        RECT 2642.400 17.670 2642.540 1683.690 ;
        RECT 2642.340 17.350 2642.600 17.670 ;
        RECT 2893.040 17.350 2893.300 17.670 ;
        RECT 2893.100 2.400 2893.240 17.350 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2646.910 1683.920 2647.230 1683.980 ;
        RECT 2649.210 1683.920 2649.530 1683.980 ;
        RECT 2646.910 1683.780 2649.530 1683.920 ;
        RECT 2646.910 1683.720 2647.230 1683.780 ;
        RECT 2649.210 1683.720 2649.530 1683.780 ;
        RECT 2649.210 17.920 2649.530 17.980 ;
        RECT 2910.950 17.920 2911.270 17.980 ;
        RECT 2649.210 17.780 2911.270 17.920 ;
        RECT 2649.210 17.720 2649.530 17.780 ;
        RECT 2910.950 17.720 2911.270 17.780 ;
      LAYER via ;
        RECT 2646.940 1683.720 2647.200 1683.980 ;
        RECT 2649.240 1683.720 2649.500 1683.980 ;
        RECT 2649.240 17.720 2649.500 17.980 ;
        RECT 2910.980 17.720 2911.240 17.980 ;
      LAYER met2 ;
        RECT 2646.860 1700.000 2647.140 1702.400 ;
        RECT 2647.000 1684.010 2647.140 1700.000 ;
        RECT 2646.940 1683.690 2647.200 1684.010 ;
        RECT 2649.240 1683.690 2649.500 1684.010 ;
        RECT 2649.300 18.010 2649.440 1683.690 ;
        RECT 2649.240 17.690 2649.500 18.010 ;
        RECT 2910.980 17.690 2911.240 18.010 ;
        RECT 2911.040 2.400 2911.180 17.690 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 858.890 45.120 859.210 45.180 ;
        RECT 1588.450 45.120 1588.770 45.180 ;
        RECT 858.890 44.980 1588.770 45.120 ;
        RECT 858.890 44.920 859.210 44.980 ;
        RECT 1588.450 44.920 1588.770 44.980 ;
      LAYER via ;
        RECT 858.920 44.920 859.180 45.180 ;
        RECT 1588.480 44.920 1588.740 45.180 ;
      LAYER met2 ;
        RECT 1590.700 1700.410 1590.980 1702.400 ;
        RECT 1588.540 1700.270 1590.980 1700.410 ;
        RECT 1588.540 45.210 1588.680 1700.270 ;
        RECT 1590.700 1700.000 1590.980 1700.270 ;
        RECT 858.920 44.890 859.180 45.210 ;
        RECT 1588.480 44.890 1588.740 45.210 ;
        RECT 858.980 2.400 859.120 44.890 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1594.965 1587.205 1595.135 1630.895 ;
        RECT 1594.965 524.365 1595.135 593.895 ;
        RECT 1595.425 331.245 1595.595 338.215 ;
        RECT 1594.965 234.685 1595.135 300.135 ;
      LAYER mcon ;
        RECT 1594.965 1630.725 1595.135 1630.895 ;
        RECT 1594.965 593.725 1595.135 593.895 ;
        RECT 1595.425 338.045 1595.595 338.215 ;
        RECT 1594.965 299.965 1595.135 300.135 ;
      LAYER met1 ;
        RECT 1594.890 1630.880 1595.210 1630.940 ;
        RECT 1594.695 1630.740 1595.210 1630.880 ;
        RECT 1594.890 1630.680 1595.210 1630.740 ;
        RECT 1594.905 1587.360 1595.195 1587.405 ;
        RECT 1595.810 1587.360 1596.130 1587.420 ;
        RECT 1594.905 1587.220 1596.130 1587.360 ;
        RECT 1594.905 1587.175 1595.195 1587.220 ;
        RECT 1595.810 1587.160 1596.130 1587.220 ;
        RECT 1595.810 1546.220 1596.130 1546.280 ;
        RECT 1594.980 1546.080 1596.130 1546.220 ;
        RECT 1594.980 1545.600 1595.120 1546.080 ;
        RECT 1595.810 1546.020 1596.130 1546.080 ;
        RECT 1594.890 1545.340 1595.210 1545.600 ;
        RECT 1594.890 1400.700 1595.210 1400.760 ;
        RECT 1595.350 1400.700 1595.670 1400.760 ;
        RECT 1594.890 1400.560 1595.670 1400.700 ;
        RECT 1594.890 1400.500 1595.210 1400.560 ;
        RECT 1595.350 1400.500 1595.670 1400.560 ;
        RECT 1594.890 1304.140 1595.210 1304.200 ;
        RECT 1595.350 1304.140 1595.670 1304.200 ;
        RECT 1594.890 1304.000 1595.670 1304.140 ;
        RECT 1594.890 1303.940 1595.210 1304.000 ;
        RECT 1595.350 1303.940 1595.670 1304.000 ;
        RECT 1594.890 1159.300 1595.210 1159.360 ;
        RECT 1595.350 1159.300 1595.670 1159.360 ;
        RECT 1594.890 1159.160 1595.670 1159.300 ;
        RECT 1594.890 1159.100 1595.210 1159.160 ;
        RECT 1595.350 1159.100 1595.670 1159.160 ;
        RECT 1594.890 1062.740 1595.210 1062.800 ;
        RECT 1595.350 1062.740 1595.670 1062.800 ;
        RECT 1594.890 1062.600 1595.670 1062.740 ;
        RECT 1594.890 1062.540 1595.210 1062.600 ;
        RECT 1595.350 1062.540 1595.670 1062.600 ;
        RECT 1594.430 979.780 1594.750 979.840 ;
        RECT 1595.350 979.780 1595.670 979.840 ;
        RECT 1594.430 979.640 1595.670 979.780 ;
        RECT 1594.430 979.580 1594.750 979.640 ;
        RECT 1595.350 979.580 1595.670 979.640 ;
        RECT 1594.890 917.900 1595.210 917.960 ;
        RECT 1595.350 917.900 1595.670 917.960 ;
        RECT 1594.890 917.760 1595.670 917.900 ;
        RECT 1594.890 917.700 1595.210 917.760 ;
        RECT 1595.350 917.700 1595.670 917.760 ;
        RECT 1594.890 910.760 1595.210 910.820 ;
        RECT 1595.350 910.760 1595.670 910.820 ;
        RECT 1594.890 910.620 1595.670 910.760 ;
        RECT 1594.890 910.560 1595.210 910.620 ;
        RECT 1595.350 910.560 1595.670 910.620 ;
        RECT 1594.430 786.660 1594.750 786.720 ;
        RECT 1595.350 786.660 1595.670 786.720 ;
        RECT 1594.430 786.520 1595.670 786.660 ;
        RECT 1594.430 786.460 1594.750 786.520 ;
        RECT 1595.350 786.460 1595.670 786.520 ;
        RECT 1594.890 765.920 1595.210 765.980 ;
        RECT 1595.350 765.920 1595.670 765.980 ;
        RECT 1594.890 765.780 1595.670 765.920 ;
        RECT 1594.890 765.720 1595.210 765.780 ;
        RECT 1595.350 765.720 1595.670 765.780 ;
        RECT 1594.890 689.900 1595.210 690.160 ;
        RECT 1594.980 689.760 1595.120 689.900 ;
        RECT 1595.350 689.760 1595.670 689.820 ;
        RECT 1594.980 689.620 1595.670 689.760 ;
        RECT 1595.350 689.560 1595.670 689.620 ;
        RECT 1594.890 593.880 1595.210 593.940 ;
        RECT 1594.695 593.740 1595.210 593.880 ;
        RECT 1594.890 593.680 1595.210 593.740 ;
        RECT 1594.890 524.520 1595.210 524.580 ;
        RECT 1594.695 524.380 1595.210 524.520 ;
        RECT 1594.890 524.320 1595.210 524.380 ;
        RECT 1594.890 496.780 1595.210 497.040 ;
        RECT 1594.980 496.640 1595.120 496.780 ;
        RECT 1595.350 496.640 1595.670 496.700 ;
        RECT 1594.980 496.500 1595.670 496.640 ;
        RECT 1595.350 496.440 1595.670 496.500 ;
        RECT 1594.890 434.560 1595.210 434.820 ;
        RECT 1594.980 434.420 1595.120 434.560 ;
        RECT 1595.350 434.420 1595.670 434.480 ;
        RECT 1594.980 434.280 1595.670 434.420 ;
        RECT 1595.350 434.220 1595.670 434.280 ;
        RECT 1595.350 338.200 1595.670 338.260 ;
        RECT 1595.155 338.060 1595.670 338.200 ;
        RECT 1595.350 338.000 1595.670 338.060 ;
        RECT 1595.350 331.400 1595.670 331.460 ;
        RECT 1595.155 331.260 1595.670 331.400 ;
        RECT 1595.350 331.200 1595.670 331.260 ;
        RECT 1594.890 300.120 1595.210 300.180 ;
        RECT 1594.695 299.980 1595.210 300.120 ;
        RECT 1594.890 299.920 1595.210 299.980 ;
        RECT 1594.890 234.840 1595.210 234.900 ;
        RECT 1594.695 234.700 1595.210 234.840 ;
        RECT 1594.890 234.640 1595.210 234.700 ;
        RECT 1595.350 158.820 1595.670 159.080 ;
        RECT 1595.440 158.400 1595.580 158.820 ;
        RECT 1595.350 158.140 1595.670 158.400 ;
        RECT 876.830 45.460 877.150 45.520 ;
        RECT 1594.430 45.460 1594.750 45.520 ;
        RECT 876.830 45.320 1594.750 45.460 ;
        RECT 876.830 45.260 877.150 45.320 ;
        RECT 1594.430 45.260 1594.750 45.320 ;
      LAYER via ;
        RECT 1594.920 1630.680 1595.180 1630.940 ;
        RECT 1595.840 1587.160 1596.100 1587.420 ;
        RECT 1595.840 1546.020 1596.100 1546.280 ;
        RECT 1594.920 1545.340 1595.180 1545.600 ;
        RECT 1594.920 1400.500 1595.180 1400.760 ;
        RECT 1595.380 1400.500 1595.640 1400.760 ;
        RECT 1594.920 1303.940 1595.180 1304.200 ;
        RECT 1595.380 1303.940 1595.640 1304.200 ;
        RECT 1594.920 1159.100 1595.180 1159.360 ;
        RECT 1595.380 1159.100 1595.640 1159.360 ;
        RECT 1594.920 1062.540 1595.180 1062.800 ;
        RECT 1595.380 1062.540 1595.640 1062.800 ;
        RECT 1594.460 979.580 1594.720 979.840 ;
        RECT 1595.380 979.580 1595.640 979.840 ;
        RECT 1594.920 917.700 1595.180 917.960 ;
        RECT 1595.380 917.700 1595.640 917.960 ;
        RECT 1594.920 910.560 1595.180 910.820 ;
        RECT 1595.380 910.560 1595.640 910.820 ;
        RECT 1594.460 786.460 1594.720 786.720 ;
        RECT 1595.380 786.460 1595.640 786.720 ;
        RECT 1594.920 765.720 1595.180 765.980 ;
        RECT 1595.380 765.720 1595.640 765.980 ;
        RECT 1594.920 689.900 1595.180 690.160 ;
        RECT 1595.380 689.560 1595.640 689.820 ;
        RECT 1594.920 593.680 1595.180 593.940 ;
        RECT 1594.920 524.320 1595.180 524.580 ;
        RECT 1594.920 496.780 1595.180 497.040 ;
        RECT 1595.380 496.440 1595.640 496.700 ;
        RECT 1594.920 434.560 1595.180 434.820 ;
        RECT 1595.380 434.220 1595.640 434.480 ;
        RECT 1595.380 338.000 1595.640 338.260 ;
        RECT 1595.380 331.200 1595.640 331.460 ;
        RECT 1594.920 299.920 1595.180 300.180 ;
        RECT 1594.920 234.640 1595.180 234.900 ;
        RECT 1595.380 158.820 1595.640 159.080 ;
        RECT 1595.380 158.140 1595.640 158.400 ;
        RECT 876.860 45.260 877.120 45.520 ;
        RECT 1594.460 45.260 1594.720 45.520 ;
      LAYER met2 ;
        RECT 1599.900 1700.410 1600.180 1702.400 ;
        RECT 1597.740 1700.270 1600.180 1700.410 ;
        RECT 1597.740 1688.850 1597.880 1700.270 ;
        RECT 1599.900 1700.000 1600.180 1700.270 ;
        RECT 1594.980 1688.710 1597.880 1688.850 ;
        RECT 1594.980 1630.970 1595.120 1688.710 ;
        RECT 1594.920 1630.650 1595.180 1630.970 ;
        RECT 1595.840 1587.130 1596.100 1587.450 ;
        RECT 1595.900 1546.310 1596.040 1587.130 ;
        RECT 1595.840 1545.990 1596.100 1546.310 ;
        RECT 1594.920 1545.310 1595.180 1545.630 ;
        RECT 1594.980 1497.090 1595.120 1545.310 ;
        RECT 1594.520 1496.950 1595.120 1497.090 ;
        RECT 1594.520 1472.610 1594.660 1496.950 ;
        RECT 1594.520 1472.470 1595.580 1472.610 ;
        RECT 1595.440 1414.130 1595.580 1472.470 ;
        RECT 1594.980 1413.990 1595.580 1414.130 ;
        RECT 1594.980 1400.790 1595.120 1413.990 ;
        RECT 1594.920 1400.470 1595.180 1400.790 ;
        RECT 1595.380 1400.470 1595.640 1400.790 ;
        RECT 1595.440 1317.570 1595.580 1400.470 ;
        RECT 1594.980 1317.430 1595.580 1317.570 ;
        RECT 1594.980 1304.230 1595.120 1317.430 ;
        RECT 1594.920 1303.910 1595.180 1304.230 ;
        RECT 1595.380 1303.910 1595.640 1304.230 ;
        RECT 1595.440 1221.010 1595.580 1303.910 ;
        RECT 1594.980 1220.870 1595.580 1221.010 ;
        RECT 1594.980 1159.390 1595.120 1220.870 ;
        RECT 1594.920 1159.070 1595.180 1159.390 ;
        RECT 1595.380 1159.070 1595.640 1159.390 ;
        RECT 1595.440 1124.450 1595.580 1159.070 ;
        RECT 1594.980 1124.310 1595.580 1124.450 ;
        RECT 1594.980 1062.830 1595.120 1124.310 ;
        RECT 1594.920 1062.510 1595.180 1062.830 ;
        RECT 1595.380 1062.510 1595.640 1062.830 ;
        RECT 1595.440 1027.890 1595.580 1062.510 ;
        RECT 1594.980 1027.750 1595.580 1027.890 ;
        RECT 1594.980 980.290 1595.120 1027.750 ;
        RECT 1594.520 980.150 1595.120 980.290 ;
        RECT 1594.520 979.870 1594.660 980.150 ;
        RECT 1594.460 979.550 1594.720 979.870 ;
        RECT 1595.380 979.550 1595.640 979.870 ;
        RECT 1595.440 917.990 1595.580 979.550 ;
        RECT 1594.920 917.670 1595.180 917.990 ;
        RECT 1595.380 917.670 1595.640 917.990 ;
        RECT 1594.980 910.850 1595.120 917.670 ;
        RECT 1594.920 910.530 1595.180 910.850 ;
        RECT 1595.380 910.530 1595.640 910.850 ;
        RECT 1595.440 834.770 1595.580 910.530 ;
        RECT 1594.980 834.630 1595.580 834.770 ;
        RECT 1594.980 787.170 1595.120 834.630 ;
        RECT 1594.520 787.030 1595.120 787.170 ;
        RECT 1594.520 786.750 1594.660 787.030 ;
        RECT 1594.460 786.430 1594.720 786.750 ;
        RECT 1595.380 786.430 1595.640 786.750 ;
        RECT 1595.440 766.010 1595.580 786.430 ;
        RECT 1594.920 765.690 1595.180 766.010 ;
        RECT 1595.380 765.690 1595.640 766.010 ;
        RECT 1594.980 690.190 1595.120 765.690 ;
        RECT 1594.920 689.870 1595.180 690.190 ;
        RECT 1595.380 689.530 1595.640 689.850 ;
        RECT 1595.440 641.650 1595.580 689.530 ;
        RECT 1594.980 641.510 1595.580 641.650 ;
        RECT 1594.980 593.970 1595.120 641.510 ;
        RECT 1594.920 593.650 1595.180 593.970 ;
        RECT 1594.920 524.290 1595.180 524.610 ;
        RECT 1594.980 497.070 1595.120 524.290 ;
        RECT 1594.920 496.750 1595.180 497.070 ;
        RECT 1595.380 496.410 1595.640 496.730 ;
        RECT 1595.440 448.530 1595.580 496.410 ;
        RECT 1594.980 448.390 1595.580 448.530 ;
        RECT 1594.980 434.850 1595.120 448.390 ;
        RECT 1594.920 434.530 1595.180 434.850 ;
        RECT 1595.380 434.190 1595.640 434.510 ;
        RECT 1595.440 338.290 1595.580 434.190 ;
        RECT 1595.380 337.970 1595.640 338.290 ;
        RECT 1595.380 331.400 1595.640 331.490 ;
        RECT 1594.980 331.260 1595.640 331.400 ;
        RECT 1594.980 300.210 1595.120 331.260 ;
        RECT 1595.380 331.170 1595.640 331.260 ;
        RECT 1594.920 299.890 1595.180 300.210 ;
        RECT 1594.920 234.610 1595.180 234.930 ;
        RECT 1594.980 234.330 1595.120 234.610 ;
        RECT 1594.980 234.190 1595.580 234.330 ;
        RECT 1595.440 159.110 1595.580 234.190 ;
        RECT 1595.380 158.790 1595.640 159.110 ;
        RECT 1595.380 158.110 1595.640 158.430 ;
        RECT 1595.440 130.290 1595.580 158.110 ;
        RECT 1594.980 130.150 1595.580 130.290 ;
        RECT 1594.980 72.490 1595.120 130.150 ;
        RECT 1594.520 72.350 1595.120 72.490 ;
        RECT 1594.520 45.550 1594.660 72.350 ;
        RECT 876.860 45.230 877.120 45.550 ;
        RECT 1594.460 45.230 1594.720 45.550 ;
        RECT 876.920 2.400 877.060 45.230 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 894.770 45.800 895.090 45.860 ;
        RECT 1607.770 45.800 1608.090 45.860 ;
        RECT 894.770 45.660 1608.090 45.800 ;
        RECT 894.770 45.600 895.090 45.660 ;
        RECT 1607.770 45.600 1608.090 45.660 ;
      LAYER via ;
        RECT 894.800 45.600 895.060 45.860 ;
        RECT 1607.800 45.600 1608.060 45.860 ;
      LAYER met2 ;
        RECT 1609.100 1700.410 1609.380 1702.400 ;
        RECT 1607.860 1700.270 1609.380 1700.410 ;
        RECT 1607.860 45.890 1608.000 1700.270 ;
        RECT 1609.100 1700.000 1609.380 1700.270 ;
        RECT 894.800 45.570 895.060 45.890 ;
        RECT 1607.800 45.570 1608.060 45.890 ;
        RECT 894.860 2.400 895.000 45.570 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 912.710 46.140 913.030 46.200 ;
        RECT 1616.050 46.140 1616.370 46.200 ;
        RECT 912.710 46.000 1616.370 46.140 ;
        RECT 912.710 45.940 913.030 46.000 ;
        RECT 1616.050 45.940 1616.370 46.000 ;
      LAYER via ;
        RECT 912.740 45.940 913.000 46.200 ;
        RECT 1616.080 45.940 1616.340 46.200 ;
      LAYER met2 ;
        RECT 1618.300 1700.410 1618.580 1702.400 ;
        RECT 1616.140 1700.270 1618.580 1700.410 ;
        RECT 1616.140 46.230 1616.280 1700.270 ;
        RECT 1618.300 1700.000 1618.580 1700.270 ;
        RECT 912.740 45.910 913.000 46.230 ;
        RECT 1616.080 45.910 1616.340 46.230 ;
        RECT 912.800 2.400 912.940 45.910 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1622.565 1449.165 1622.735 1496.935 ;
        RECT 1622.105 1304.325 1622.275 1318.095 ;
        RECT 1622.105 1111.205 1622.275 1124.975 ;
        RECT 1622.105 1097.605 1622.275 1110.695 ;
        RECT 1622.105 1014.305 1622.275 1028.415 ;
        RECT 1622.105 959.225 1622.275 980.475 ;
        RECT 1622.565 807.245 1622.735 855.355 ;
        RECT 1623.025 710.685 1623.195 758.795 ;
        RECT 1622.105 614.125 1622.275 662.235 ;
        RECT 1622.565 427.805 1622.735 475.915 ;
        RECT 1622.105 276.505 1622.275 289.595 ;
        RECT 1622.565 227.885 1622.735 275.995 ;
      LAYER mcon ;
        RECT 1622.565 1496.765 1622.735 1496.935 ;
        RECT 1622.105 1317.925 1622.275 1318.095 ;
        RECT 1622.105 1124.805 1622.275 1124.975 ;
        RECT 1622.105 1110.525 1622.275 1110.695 ;
        RECT 1622.105 1028.245 1622.275 1028.415 ;
        RECT 1622.105 980.305 1622.275 980.475 ;
        RECT 1622.565 855.185 1622.735 855.355 ;
        RECT 1623.025 758.625 1623.195 758.795 ;
        RECT 1622.105 662.065 1622.275 662.235 ;
        RECT 1622.565 475.745 1622.735 475.915 ;
        RECT 1622.105 289.425 1622.275 289.595 ;
        RECT 1622.565 275.825 1622.735 275.995 ;
      LAYER met1 ;
        RECT 1622.030 1666.580 1622.350 1666.640 ;
        RECT 1625.250 1666.580 1625.570 1666.640 ;
        RECT 1622.030 1666.440 1625.570 1666.580 ;
        RECT 1622.030 1666.380 1622.350 1666.440 ;
        RECT 1625.250 1666.380 1625.570 1666.440 ;
        RECT 1622.490 1608.100 1622.810 1608.160 ;
        RECT 1622.120 1607.960 1622.810 1608.100 ;
        RECT 1622.120 1607.820 1622.260 1607.960 ;
        RECT 1622.490 1607.900 1622.810 1607.960 ;
        RECT 1622.030 1607.560 1622.350 1607.820 ;
        RECT 1621.110 1545.880 1621.430 1545.940 ;
        RECT 1622.490 1545.880 1622.810 1545.940 ;
        RECT 1621.110 1545.740 1622.810 1545.880 ;
        RECT 1621.110 1545.680 1621.430 1545.740 ;
        RECT 1622.490 1545.680 1622.810 1545.740 ;
        RECT 1622.490 1496.920 1622.810 1496.980 ;
        RECT 1622.295 1496.780 1622.810 1496.920 ;
        RECT 1622.490 1496.720 1622.810 1496.780 ;
        RECT 1622.490 1449.320 1622.810 1449.380 ;
        RECT 1622.295 1449.180 1622.810 1449.320 ;
        RECT 1622.490 1449.120 1622.810 1449.180 ;
        RECT 1622.030 1401.040 1622.350 1401.100 ;
        RECT 1623.410 1401.040 1623.730 1401.100 ;
        RECT 1622.030 1400.900 1623.730 1401.040 ;
        RECT 1622.030 1400.840 1622.350 1400.900 ;
        RECT 1623.410 1400.840 1623.730 1400.900 ;
        RECT 1622.030 1318.080 1622.350 1318.140 ;
        RECT 1621.835 1317.940 1622.350 1318.080 ;
        RECT 1622.030 1317.880 1622.350 1317.940 ;
        RECT 1622.030 1304.480 1622.350 1304.540 ;
        RECT 1621.835 1304.340 1622.350 1304.480 ;
        RECT 1622.030 1304.280 1622.350 1304.340 ;
        RECT 1621.110 1227.300 1621.430 1227.360 ;
        RECT 1622.030 1227.300 1622.350 1227.360 ;
        RECT 1621.110 1227.160 1622.350 1227.300 ;
        RECT 1621.110 1227.100 1621.430 1227.160 ;
        RECT 1622.030 1227.100 1622.350 1227.160 ;
        RECT 1621.110 1183.440 1621.430 1183.500 ;
        RECT 1622.030 1183.440 1622.350 1183.500 ;
        RECT 1621.110 1183.300 1622.350 1183.440 ;
        RECT 1621.110 1183.240 1621.430 1183.300 ;
        RECT 1622.030 1183.240 1622.350 1183.300 ;
        RECT 1622.030 1124.960 1622.350 1125.020 ;
        RECT 1621.835 1124.820 1622.350 1124.960 ;
        RECT 1622.030 1124.760 1622.350 1124.820 ;
        RECT 1622.030 1111.360 1622.350 1111.420 ;
        RECT 1621.835 1111.220 1622.350 1111.360 ;
        RECT 1622.030 1111.160 1622.350 1111.220 ;
        RECT 1622.030 1110.680 1622.350 1110.740 ;
        RECT 1621.835 1110.540 1622.350 1110.680 ;
        RECT 1622.030 1110.480 1622.350 1110.540 ;
        RECT 1622.030 1097.760 1622.350 1097.820 ;
        RECT 1621.835 1097.620 1622.350 1097.760 ;
        RECT 1622.030 1097.560 1622.350 1097.620 ;
        RECT 1622.030 1028.400 1622.350 1028.460 ;
        RECT 1621.835 1028.260 1622.350 1028.400 ;
        RECT 1622.030 1028.200 1622.350 1028.260 ;
        RECT 1622.030 1014.460 1622.350 1014.520 ;
        RECT 1621.835 1014.320 1622.350 1014.460 ;
        RECT 1622.030 1014.260 1622.350 1014.320 ;
        RECT 1622.030 980.460 1622.350 980.520 ;
        RECT 1621.835 980.320 1622.350 980.460 ;
        RECT 1622.030 980.260 1622.350 980.320 ;
        RECT 1622.030 959.380 1622.350 959.440 ;
        RECT 1621.835 959.240 1622.350 959.380 ;
        RECT 1622.030 959.180 1622.350 959.240 ;
        RECT 1621.110 958.700 1621.430 958.760 ;
        RECT 1622.030 958.700 1622.350 958.760 ;
        RECT 1621.110 958.560 1622.350 958.700 ;
        RECT 1621.110 958.500 1621.430 958.560 ;
        RECT 1622.030 958.500 1622.350 958.560 ;
        RECT 1621.110 877.100 1621.430 877.160 ;
        RECT 1622.490 877.100 1622.810 877.160 ;
        RECT 1621.110 876.960 1622.810 877.100 ;
        RECT 1621.110 876.900 1621.430 876.960 ;
        RECT 1622.490 876.900 1622.810 876.960 ;
        RECT 1622.490 855.340 1622.810 855.400 ;
        RECT 1622.295 855.200 1622.810 855.340 ;
        RECT 1622.490 855.140 1622.810 855.200 ;
        RECT 1622.490 807.400 1622.810 807.460 ;
        RECT 1622.295 807.260 1622.810 807.400 ;
        RECT 1622.490 807.200 1622.810 807.260 ;
        RECT 1622.950 758.780 1623.270 758.840 ;
        RECT 1622.755 758.640 1623.270 758.780 ;
        RECT 1622.950 758.580 1623.270 758.640 ;
        RECT 1622.950 710.840 1623.270 710.900 ;
        RECT 1622.755 710.700 1623.270 710.840 ;
        RECT 1622.950 710.640 1623.270 710.700 ;
        RECT 1622.045 662.220 1622.335 662.265 ;
        RECT 1622.490 662.220 1622.810 662.280 ;
        RECT 1622.045 662.080 1622.810 662.220 ;
        RECT 1622.045 662.035 1622.335 662.080 ;
        RECT 1622.490 662.020 1622.810 662.080 ;
        RECT 1622.030 614.280 1622.350 614.340 ;
        RECT 1621.835 614.140 1622.350 614.280 ;
        RECT 1622.030 614.080 1622.350 614.140 ;
        RECT 1621.110 590.140 1621.430 590.200 ;
        RECT 1622.030 590.140 1622.350 590.200 ;
        RECT 1621.110 590.000 1622.350 590.140 ;
        RECT 1621.110 589.940 1621.430 590.000 ;
        RECT 1622.030 589.940 1622.350 590.000 ;
        RECT 1622.030 524.180 1622.350 524.240 ;
        RECT 1623.410 524.180 1623.730 524.240 ;
        RECT 1622.030 524.040 1623.730 524.180 ;
        RECT 1622.030 523.980 1622.350 524.040 ;
        RECT 1623.410 523.980 1623.730 524.040 ;
        RECT 1622.490 475.900 1622.810 475.960 ;
        RECT 1622.295 475.760 1622.810 475.900 ;
        RECT 1622.490 475.700 1622.810 475.760 ;
        RECT 1622.490 427.960 1622.810 428.020 ;
        RECT 1622.295 427.820 1622.810 427.960 ;
        RECT 1622.490 427.760 1622.810 427.820 ;
        RECT 1622.030 338.200 1622.350 338.260 ;
        RECT 1622.490 338.200 1622.810 338.260 ;
        RECT 1622.030 338.060 1622.810 338.200 ;
        RECT 1622.030 338.000 1622.350 338.060 ;
        RECT 1622.490 338.000 1622.810 338.060 ;
        RECT 1622.030 289.580 1622.350 289.640 ;
        RECT 1621.835 289.440 1622.350 289.580 ;
        RECT 1622.030 289.380 1622.350 289.440 ;
        RECT 1622.045 276.475 1622.335 276.705 ;
        RECT 1622.120 275.980 1622.260 276.475 ;
        RECT 1622.505 275.980 1622.795 276.025 ;
        RECT 1622.120 275.840 1622.795 275.980 ;
        RECT 1622.505 275.795 1622.795 275.840 ;
        RECT 1622.490 228.040 1622.810 228.100 ;
        RECT 1622.295 227.900 1622.810 228.040 ;
        RECT 1622.490 227.840 1622.810 227.900 ;
        RECT 1622.490 131.820 1622.810 131.880 ;
        RECT 1622.120 131.680 1622.810 131.820 ;
        RECT 1622.120 131.540 1622.260 131.680 ;
        RECT 1622.490 131.620 1622.810 131.680 ;
        RECT 1622.030 131.280 1622.350 131.540 ;
        RECT 1622.030 96.800 1622.350 96.860 ;
        RECT 1622.490 96.800 1622.810 96.860 ;
        RECT 1622.030 96.660 1622.810 96.800 ;
        RECT 1622.030 96.600 1622.350 96.660 ;
        RECT 1622.490 96.600 1622.810 96.660 ;
        RECT 930.190 46.480 930.510 46.540 ;
        RECT 1622.030 46.480 1622.350 46.540 ;
        RECT 930.190 46.340 1622.350 46.480 ;
        RECT 930.190 46.280 930.510 46.340 ;
        RECT 1622.030 46.280 1622.350 46.340 ;
      LAYER via ;
        RECT 1622.060 1666.380 1622.320 1666.640 ;
        RECT 1625.280 1666.380 1625.540 1666.640 ;
        RECT 1622.520 1607.900 1622.780 1608.160 ;
        RECT 1622.060 1607.560 1622.320 1607.820 ;
        RECT 1621.140 1545.680 1621.400 1545.940 ;
        RECT 1622.520 1545.680 1622.780 1545.940 ;
        RECT 1622.520 1496.720 1622.780 1496.980 ;
        RECT 1622.520 1449.120 1622.780 1449.380 ;
        RECT 1622.060 1400.840 1622.320 1401.100 ;
        RECT 1623.440 1400.840 1623.700 1401.100 ;
        RECT 1622.060 1317.880 1622.320 1318.140 ;
        RECT 1622.060 1304.280 1622.320 1304.540 ;
        RECT 1621.140 1227.100 1621.400 1227.360 ;
        RECT 1622.060 1227.100 1622.320 1227.360 ;
        RECT 1621.140 1183.240 1621.400 1183.500 ;
        RECT 1622.060 1183.240 1622.320 1183.500 ;
        RECT 1622.060 1124.760 1622.320 1125.020 ;
        RECT 1622.060 1111.160 1622.320 1111.420 ;
        RECT 1622.060 1110.480 1622.320 1110.740 ;
        RECT 1622.060 1097.560 1622.320 1097.820 ;
        RECT 1622.060 1028.200 1622.320 1028.460 ;
        RECT 1622.060 1014.260 1622.320 1014.520 ;
        RECT 1622.060 980.260 1622.320 980.520 ;
        RECT 1622.060 959.180 1622.320 959.440 ;
        RECT 1621.140 958.500 1621.400 958.760 ;
        RECT 1622.060 958.500 1622.320 958.760 ;
        RECT 1621.140 876.900 1621.400 877.160 ;
        RECT 1622.520 876.900 1622.780 877.160 ;
        RECT 1622.520 855.140 1622.780 855.400 ;
        RECT 1622.520 807.200 1622.780 807.460 ;
        RECT 1622.980 758.580 1623.240 758.840 ;
        RECT 1622.980 710.640 1623.240 710.900 ;
        RECT 1622.520 662.020 1622.780 662.280 ;
        RECT 1622.060 614.080 1622.320 614.340 ;
        RECT 1621.140 589.940 1621.400 590.200 ;
        RECT 1622.060 589.940 1622.320 590.200 ;
        RECT 1622.060 523.980 1622.320 524.240 ;
        RECT 1623.440 523.980 1623.700 524.240 ;
        RECT 1622.520 475.700 1622.780 475.960 ;
        RECT 1622.520 427.760 1622.780 428.020 ;
        RECT 1622.060 338.000 1622.320 338.260 ;
        RECT 1622.520 338.000 1622.780 338.260 ;
        RECT 1622.060 289.380 1622.320 289.640 ;
        RECT 1622.520 227.840 1622.780 228.100 ;
        RECT 1622.520 131.620 1622.780 131.880 ;
        RECT 1622.060 131.280 1622.320 131.540 ;
        RECT 1622.060 96.600 1622.320 96.860 ;
        RECT 1622.520 96.600 1622.780 96.860 ;
        RECT 930.220 46.280 930.480 46.540 ;
        RECT 1622.060 46.280 1622.320 46.540 ;
      LAYER met2 ;
        RECT 1627.500 1700.410 1627.780 1702.400 ;
        RECT 1625.340 1700.270 1627.780 1700.410 ;
        RECT 1625.340 1666.670 1625.480 1700.270 ;
        RECT 1627.500 1700.000 1627.780 1700.270 ;
        RECT 1622.060 1666.350 1622.320 1666.670 ;
        RECT 1625.280 1666.350 1625.540 1666.670 ;
        RECT 1622.120 1642.610 1622.260 1666.350 ;
        RECT 1622.120 1642.470 1622.720 1642.610 ;
        RECT 1622.580 1608.190 1622.720 1642.470 ;
        RECT 1622.520 1607.870 1622.780 1608.190 ;
        RECT 1622.060 1607.530 1622.320 1607.850 ;
        RECT 1622.120 1593.765 1622.260 1607.530 ;
        RECT 1621.130 1593.395 1621.410 1593.765 ;
        RECT 1622.050 1593.395 1622.330 1593.765 ;
        RECT 1621.200 1545.970 1621.340 1593.395 ;
        RECT 1621.140 1545.650 1621.400 1545.970 ;
        RECT 1622.520 1545.650 1622.780 1545.970 ;
        RECT 1622.580 1512.050 1622.720 1545.650 ;
        RECT 1622.580 1511.910 1623.180 1512.050 ;
        RECT 1623.040 1510.690 1623.180 1511.910 ;
        RECT 1622.580 1510.550 1623.180 1510.690 ;
        RECT 1622.580 1497.010 1622.720 1510.550 ;
        RECT 1622.520 1496.690 1622.780 1497.010 ;
        RECT 1622.520 1449.090 1622.780 1449.410 ;
        RECT 1622.580 1448.925 1622.720 1449.090 ;
        RECT 1622.510 1448.555 1622.790 1448.925 ;
        RECT 1623.430 1448.555 1623.710 1448.925 ;
        RECT 1623.500 1401.130 1623.640 1448.555 ;
        RECT 1622.060 1400.810 1622.320 1401.130 ;
        RECT 1623.440 1400.810 1623.700 1401.130 ;
        RECT 1622.120 1400.530 1622.260 1400.810 ;
        RECT 1622.120 1400.390 1622.720 1400.530 ;
        RECT 1622.580 1383.530 1622.720 1400.390 ;
        RECT 1622.120 1383.390 1622.720 1383.530 ;
        RECT 1622.120 1318.170 1622.260 1383.390 ;
        RECT 1622.060 1317.850 1622.320 1318.170 ;
        RECT 1622.060 1304.250 1622.320 1304.570 ;
        RECT 1622.120 1303.970 1622.260 1304.250 ;
        RECT 1622.120 1303.830 1622.720 1303.970 ;
        RECT 1622.580 1279.490 1622.720 1303.830 ;
        RECT 1622.120 1279.350 1622.720 1279.490 ;
        RECT 1622.120 1227.390 1622.260 1279.350 ;
        RECT 1621.140 1227.070 1621.400 1227.390 ;
        RECT 1622.060 1227.070 1622.320 1227.390 ;
        RECT 1621.200 1183.530 1621.340 1227.070 ;
        RECT 1621.140 1183.210 1621.400 1183.530 ;
        RECT 1622.060 1183.210 1622.320 1183.530 ;
        RECT 1622.120 1125.050 1622.260 1183.210 ;
        RECT 1622.060 1124.730 1622.320 1125.050 ;
        RECT 1622.060 1111.130 1622.320 1111.450 ;
        RECT 1622.120 1110.770 1622.260 1111.130 ;
        RECT 1622.060 1110.450 1622.320 1110.770 ;
        RECT 1622.060 1097.530 1622.320 1097.850 ;
        RECT 1622.120 1028.490 1622.260 1097.530 ;
        RECT 1622.060 1028.170 1622.320 1028.490 ;
        RECT 1622.060 1014.230 1622.320 1014.550 ;
        RECT 1622.120 980.550 1622.260 1014.230 ;
        RECT 1622.060 980.230 1622.320 980.550 ;
        RECT 1622.060 959.150 1622.320 959.470 ;
        RECT 1622.120 958.790 1622.260 959.150 ;
        RECT 1621.140 958.470 1621.400 958.790 ;
        RECT 1622.060 958.470 1622.320 958.790 ;
        RECT 1621.200 911.045 1621.340 958.470 ;
        RECT 1621.130 910.675 1621.410 911.045 ;
        RECT 1622.510 910.675 1622.790 911.045 ;
        RECT 1622.580 877.190 1622.720 910.675 ;
        RECT 1621.140 876.870 1621.400 877.190 ;
        RECT 1622.520 876.870 1622.780 877.190 ;
        RECT 1621.200 855.965 1621.340 876.870 ;
        RECT 1621.130 855.595 1621.410 855.965 ;
        RECT 1622.050 855.850 1622.330 855.965 ;
        RECT 1622.050 855.710 1622.720 855.850 ;
        RECT 1622.050 855.595 1622.330 855.710 ;
        RECT 1622.580 855.430 1622.720 855.710 ;
        RECT 1622.520 855.110 1622.780 855.430 ;
        RECT 1622.520 807.170 1622.780 807.490 ;
        RECT 1622.580 806.890 1622.720 807.170 ;
        RECT 1622.580 806.750 1623.640 806.890 ;
        RECT 1623.500 759.290 1623.640 806.750 ;
        RECT 1623.040 759.150 1623.640 759.290 ;
        RECT 1623.040 758.870 1623.180 759.150 ;
        RECT 1622.980 758.550 1623.240 758.870 ;
        RECT 1622.980 710.610 1623.240 710.930 ;
        RECT 1623.040 668.850 1623.180 710.610 ;
        RECT 1622.580 668.710 1623.180 668.850 ;
        RECT 1622.580 662.310 1622.720 668.710 ;
        RECT 1622.520 661.990 1622.780 662.310 ;
        RECT 1622.060 614.050 1622.320 614.370 ;
        RECT 1622.120 613.885 1622.260 614.050 ;
        RECT 1621.130 613.515 1621.410 613.885 ;
        RECT 1622.050 613.515 1622.330 613.885 ;
        RECT 1621.200 590.230 1621.340 613.515 ;
        RECT 1621.140 589.910 1621.400 590.230 ;
        RECT 1622.060 589.910 1622.320 590.230 ;
        RECT 1622.120 524.270 1622.260 589.910 ;
        RECT 1622.060 523.950 1622.320 524.270 ;
        RECT 1623.440 523.950 1623.700 524.270 ;
        RECT 1623.500 476.525 1623.640 523.950 ;
        RECT 1622.510 476.155 1622.790 476.525 ;
        RECT 1623.430 476.155 1623.710 476.525 ;
        RECT 1622.580 475.990 1622.720 476.155 ;
        RECT 1622.520 475.670 1622.780 475.990 ;
        RECT 1622.520 427.730 1622.780 428.050 ;
        RECT 1622.580 338.290 1622.720 427.730 ;
        RECT 1622.060 337.970 1622.320 338.290 ;
        RECT 1622.520 337.970 1622.780 338.290 ;
        RECT 1622.120 289.670 1622.260 337.970 ;
        RECT 1622.060 289.350 1622.320 289.670 ;
        RECT 1622.520 227.810 1622.780 228.130 ;
        RECT 1622.580 131.910 1622.720 227.810 ;
        RECT 1622.520 131.590 1622.780 131.910 ;
        RECT 1622.060 131.250 1622.320 131.570 ;
        RECT 1622.120 96.890 1622.260 131.250 ;
        RECT 1622.060 96.570 1622.320 96.890 ;
        RECT 1622.520 96.570 1622.780 96.890 ;
        RECT 1622.580 72.490 1622.720 96.570 ;
        RECT 1622.120 72.350 1622.720 72.490 ;
        RECT 1622.120 46.570 1622.260 72.350 ;
        RECT 930.220 46.250 930.480 46.570 ;
        RECT 1622.060 46.250 1622.320 46.570 ;
        RECT 930.280 2.400 930.420 46.250 ;
        RECT 930.070 -4.800 930.630 2.400 ;
      LAYER via2 ;
        RECT 1621.130 1593.440 1621.410 1593.720 ;
        RECT 1622.050 1593.440 1622.330 1593.720 ;
        RECT 1622.510 1448.600 1622.790 1448.880 ;
        RECT 1623.430 1448.600 1623.710 1448.880 ;
        RECT 1621.130 910.720 1621.410 911.000 ;
        RECT 1622.510 910.720 1622.790 911.000 ;
        RECT 1621.130 855.640 1621.410 855.920 ;
        RECT 1622.050 855.640 1622.330 855.920 ;
        RECT 1621.130 613.560 1621.410 613.840 ;
        RECT 1622.050 613.560 1622.330 613.840 ;
        RECT 1622.510 476.200 1622.790 476.480 ;
        RECT 1623.430 476.200 1623.710 476.480 ;
      LAYER met3 ;
        RECT 1621.105 1593.730 1621.435 1593.745 ;
        RECT 1622.025 1593.730 1622.355 1593.745 ;
        RECT 1621.105 1593.430 1622.355 1593.730 ;
        RECT 1621.105 1593.415 1621.435 1593.430 ;
        RECT 1622.025 1593.415 1622.355 1593.430 ;
        RECT 1622.485 1448.890 1622.815 1448.905 ;
        RECT 1623.405 1448.890 1623.735 1448.905 ;
        RECT 1622.485 1448.590 1623.735 1448.890 ;
        RECT 1622.485 1448.575 1622.815 1448.590 ;
        RECT 1623.405 1448.575 1623.735 1448.590 ;
        RECT 1621.105 911.010 1621.435 911.025 ;
        RECT 1622.485 911.010 1622.815 911.025 ;
        RECT 1621.105 910.710 1622.815 911.010 ;
        RECT 1621.105 910.695 1621.435 910.710 ;
        RECT 1622.485 910.695 1622.815 910.710 ;
        RECT 1621.105 855.930 1621.435 855.945 ;
        RECT 1622.025 855.930 1622.355 855.945 ;
        RECT 1621.105 855.630 1622.355 855.930 ;
        RECT 1621.105 855.615 1621.435 855.630 ;
        RECT 1622.025 855.615 1622.355 855.630 ;
        RECT 1621.105 613.850 1621.435 613.865 ;
        RECT 1622.025 613.850 1622.355 613.865 ;
        RECT 1621.105 613.550 1622.355 613.850 ;
        RECT 1621.105 613.535 1621.435 613.550 ;
        RECT 1622.025 613.535 1622.355 613.550 ;
        RECT 1622.485 476.490 1622.815 476.505 ;
        RECT 1623.405 476.490 1623.735 476.505 ;
        RECT 1622.485 476.190 1623.735 476.490 ;
        RECT 1622.485 476.175 1622.815 476.190 ;
        RECT 1623.405 476.175 1623.735 476.190 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 948.130 46.820 948.450 46.880 ;
        RECT 1635.370 46.820 1635.690 46.880 ;
        RECT 948.130 46.680 1635.690 46.820 ;
        RECT 948.130 46.620 948.450 46.680 ;
        RECT 1635.370 46.620 1635.690 46.680 ;
      LAYER via ;
        RECT 948.160 46.620 948.420 46.880 ;
        RECT 1635.400 46.620 1635.660 46.880 ;
      LAYER met2 ;
        RECT 1636.700 1700.410 1636.980 1702.400 ;
        RECT 1635.460 1700.270 1636.980 1700.410 ;
        RECT 1635.460 46.910 1635.600 1700.270 ;
        RECT 1636.700 1700.000 1636.980 1700.270 ;
        RECT 948.160 46.590 948.420 46.910 ;
        RECT 1635.400 46.590 1635.660 46.910 ;
        RECT 948.220 2.400 948.360 46.590 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 966.070 47.160 966.390 47.220 ;
        RECT 1643.650 47.160 1643.970 47.220 ;
        RECT 966.070 47.020 1643.970 47.160 ;
        RECT 966.070 46.960 966.390 47.020 ;
        RECT 1643.650 46.960 1643.970 47.020 ;
      LAYER via ;
        RECT 966.100 46.960 966.360 47.220 ;
        RECT 1643.680 46.960 1643.940 47.220 ;
      LAYER met2 ;
        RECT 1645.900 1700.410 1646.180 1702.400 ;
        RECT 1643.740 1700.270 1646.180 1700.410 ;
        RECT 1643.740 47.250 1643.880 1700.270 ;
        RECT 1645.900 1700.000 1646.180 1700.270 ;
        RECT 966.100 46.930 966.360 47.250 ;
        RECT 1643.680 46.930 1643.940 47.250 ;
        RECT 966.160 2.400 966.300 46.930 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1650.165 324.785 1650.335 331.415 ;
        RECT 1649.705 269.025 1649.875 317.475 ;
      LAYER mcon ;
        RECT 1650.165 331.245 1650.335 331.415 ;
        RECT 1649.705 317.305 1649.875 317.475 ;
      LAYER met1 ;
        RECT 1650.090 1642.440 1650.410 1642.500 ;
        RECT 1652.850 1642.440 1653.170 1642.500 ;
        RECT 1650.090 1642.300 1653.170 1642.440 ;
        RECT 1650.090 1642.240 1650.410 1642.300 ;
        RECT 1652.850 1642.240 1653.170 1642.300 ;
        RECT 1650.090 1463.060 1650.410 1463.320 ;
        RECT 1650.180 1462.640 1650.320 1463.060 ;
        RECT 1650.090 1462.380 1650.410 1462.640 ;
        RECT 1650.090 1366.500 1650.410 1366.760 ;
        RECT 1650.180 1366.080 1650.320 1366.500 ;
        RECT 1650.090 1365.820 1650.410 1366.080 ;
        RECT 1650.090 1269.940 1650.410 1270.200 ;
        RECT 1650.180 1269.520 1650.320 1269.940 ;
        RECT 1650.090 1269.260 1650.410 1269.520 ;
        RECT 1650.550 1173.240 1650.870 1173.300 ;
        RECT 1650.180 1173.100 1650.870 1173.240 ;
        RECT 1650.180 1172.960 1650.320 1173.100 ;
        RECT 1650.550 1173.040 1650.870 1173.100 ;
        RECT 1650.090 1172.700 1650.410 1172.960 ;
        RECT 1650.550 1076.680 1650.870 1076.740 ;
        RECT 1650.180 1076.540 1650.870 1076.680 ;
        RECT 1650.180 1076.400 1650.320 1076.540 ;
        RECT 1650.550 1076.480 1650.870 1076.540 ;
        RECT 1650.090 1076.140 1650.410 1076.400 ;
        RECT 1650.550 980.120 1650.870 980.180 ;
        RECT 1650.180 979.980 1650.870 980.120 ;
        RECT 1650.180 979.840 1650.320 979.980 ;
        RECT 1650.550 979.920 1650.870 979.980 ;
        RECT 1650.090 979.580 1650.410 979.840 ;
        RECT 1650.090 531.320 1650.410 531.380 ;
        RECT 1651.010 531.320 1651.330 531.380 ;
        RECT 1650.090 531.180 1651.330 531.320 ;
        RECT 1650.090 531.120 1650.410 531.180 ;
        RECT 1651.010 531.120 1651.330 531.180 ;
        RECT 1650.090 427.960 1650.410 428.020 ;
        RECT 1650.550 427.960 1650.870 428.020 ;
        RECT 1650.090 427.820 1650.870 427.960 ;
        RECT 1650.090 427.760 1650.410 427.820 ;
        RECT 1650.550 427.760 1650.870 427.820 ;
        RECT 1650.090 380.360 1650.410 380.420 ;
        RECT 1650.090 380.220 1650.780 380.360 ;
        RECT 1650.090 380.160 1650.410 380.220 ;
        RECT 1650.640 379.740 1650.780 380.220 ;
        RECT 1650.550 379.480 1650.870 379.740 ;
        RECT 1650.090 331.400 1650.410 331.460 ;
        RECT 1649.895 331.260 1650.410 331.400 ;
        RECT 1650.090 331.200 1650.410 331.260 ;
        RECT 1650.090 324.940 1650.410 325.000 ;
        RECT 1649.895 324.800 1650.410 324.940 ;
        RECT 1650.090 324.740 1650.410 324.800 ;
        RECT 1649.645 317.460 1649.935 317.505 ;
        RECT 1650.090 317.460 1650.410 317.520 ;
        RECT 1649.645 317.320 1650.410 317.460 ;
        RECT 1649.645 317.275 1649.935 317.320 ;
        RECT 1650.090 317.260 1650.410 317.320 ;
        RECT 1649.630 269.180 1649.950 269.240 ;
        RECT 1649.435 269.040 1649.950 269.180 ;
        RECT 1649.630 268.980 1649.950 269.040 ;
        RECT 1649.630 72.660 1649.950 72.720 ;
        RECT 1650.550 72.660 1650.870 72.720 ;
        RECT 1649.630 72.520 1650.870 72.660 ;
        RECT 1649.630 72.460 1649.950 72.520 ;
        RECT 1650.550 72.460 1650.870 72.520 ;
        RECT 984.010 47.500 984.330 47.560 ;
        RECT 1650.090 47.500 1650.410 47.560 ;
        RECT 984.010 47.360 1650.410 47.500 ;
        RECT 984.010 47.300 984.330 47.360 ;
        RECT 1650.090 47.300 1650.410 47.360 ;
      LAYER via ;
        RECT 1650.120 1642.240 1650.380 1642.500 ;
        RECT 1652.880 1642.240 1653.140 1642.500 ;
        RECT 1650.120 1463.060 1650.380 1463.320 ;
        RECT 1650.120 1462.380 1650.380 1462.640 ;
        RECT 1650.120 1366.500 1650.380 1366.760 ;
        RECT 1650.120 1365.820 1650.380 1366.080 ;
        RECT 1650.120 1269.940 1650.380 1270.200 ;
        RECT 1650.120 1269.260 1650.380 1269.520 ;
        RECT 1650.580 1173.040 1650.840 1173.300 ;
        RECT 1650.120 1172.700 1650.380 1172.960 ;
        RECT 1650.580 1076.480 1650.840 1076.740 ;
        RECT 1650.120 1076.140 1650.380 1076.400 ;
        RECT 1650.580 979.920 1650.840 980.180 ;
        RECT 1650.120 979.580 1650.380 979.840 ;
        RECT 1650.120 531.120 1650.380 531.380 ;
        RECT 1651.040 531.120 1651.300 531.380 ;
        RECT 1650.120 427.760 1650.380 428.020 ;
        RECT 1650.580 427.760 1650.840 428.020 ;
        RECT 1650.120 380.160 1650.380 380.420 ;
        RECT 1650.580 379.480 1650.840 379.740 ;
        RECT 1650.120 331.200 1650.380 331.460 ;
        RECT 1650.120 324.740 1650.380 325.000 ;
        RECT 1650.120 317.260 1650.380 317.520 ;
        RECT 1649.660 268.980 1649.920 269.240 ;
        RECT 1649.660 72.460 1649.920 72.720 ;
        RECT 1650.580 72.460 1650.840 72.720 ;
        RECT 984.040 47.300 984.300 47.560 ;
        RECT 1650.120 47.300 1650.380 47.560 ;
      LAYER met2 ;
        RECT 1655.100 1700.410 1655.380 1702.400 ;
        RECT 1652.940 1700.270 1655.380 1700.410 ;
        RECT 1652.940 1642.530 1653.080 1700.270 ;
        RECT 1655.100 1700.000 1655.380 1700.270 ;
        RECT 1650.120 1642.210 1650.380 1642.530 ;
        RECT 1652.880 1642.210 1653.140 1642.530 ;
        RECT 1650.180 1463.350 1650.320 1642.210 ;
        RECT 1650.120 1463.030 1650.380 1463.350 ;
        RECT 1650.120 1462.350 1650.380 1462.670 ;
        RECT 1650.180 1366.790 1650.320 1462.350 ;
        RECT 1650.120 1366.470 1650.380 1366.790 ;
        RECT 1650.120 1365.790 1650.380 1366.110 ;
        RECT 1650.180 1270.230 1650.320 1365.790 ;
        RECT 1650.120 1269.910 1650.380 1270.230 ;
        RECT 1650.120 1269.230 1650.380 1269.550 ;
        RECT 1650.180 1207.410 1650.320 1269.230 ;
        RECT 1650.180 1207.270 1650.780 1207.410 ;
        RECT 1650.640 1173.330 1650.780 1207.270 ;
        RECT 1650.580 1173.010 1650.840 1173.330 ;
        RECT 1650.120 1172.670 1650.380 1172.990 ;
        RECT 1650.180 1110.850 1650.320 1172.670 ;
        RECT 1650.180 1110.710 1650.780 1110.850 ;
        RECT 1650.640 1076.770 1650.780 1110.710 ;
        RECT 1650.580 1076.450 1650.840 1076.770 ;
        RECT 1650.120 1076.110 1650.380 1076.430 ;
        RECT 1650.180 1014.290 1650.320 1076.110 ;
        RECT 1650.180 1014.150 1650.780 1014.290 ;
        RECT 1650.640 980.210 1650.780 1014.150 ;
        RECT 1650.580 979.890 1650.840 980.210 ;
        RECT 1650.120 979.550 1650.380 979.870 ;
        RECT 1650.180 787.170 1650.320 979.550 ;
        RECT 1649.720 787.030 1650.320 787.170 ;
        RECT 1649.720 786.490 1649.860 787.030 ;
        RECT 1649.720 786.350 1650.320 786.490 ;
        RECT 1650.180 686.530 1650.320 786.350 ;
        RECT 1650.180 686.390 1651.240 686.530 ;
        RECT 1651.100 676.445 1651.240 686.390 ;
        RECT 1651.030 676.075 1651.310 676.445 ;
        RECT 1649.650 675.395 1649.930 675.765 ;
        RECT 1649.720 628.050 1649.860 675.395 ;
        RECT 1649.720 627.910 1650.320 628.050 ;
        RECT 1650.180 593.880 1650.320 627.910 ;
        RECT 1650.180 593.740 1650.780 593.880 ;
        RECT 1650.640 592.690 1650.780 593.740 ;
        RECT 1650.180 592.550 1650.780 592.690 ;
        RECT 1650.180 531.410 1650.320 592.550 ;
        RECT 1650.120 531.090 1650.380 531.410 ;
        RECT 1651.040 531.090 1651.300 531.410 ;
        RECT 1651.100 476.410 1651.240 531.090 ;
        RECT 1650.640 476.270 1651.240 476.410 ;
        RECT 1650.640 428.050 1650.780 476.270 ;
        RECT 1650.120 427.730 1650.380 428.050 ;
        RECT 1650.580 427.730 1650.840 428.050 ;
        RECT 1650.180 380.450 1650.320 427.730 ;
        RECT 1650.120 380.130 1650.380 380.450 ;
        RECT 1650.580 379.450 1650.840 379.770 ;
        RECT 1650.640 379.170 1650.780 379.450 ;
        RECT 1650.180 379.030 1650.780 379.170 ;
        RECT 1650.180 331.490 1650.320 379.030 ;
        RECT 1650.120 331.170 1650.380 331.490 ;
        RECT 1650.120 324.710 1650.380 325.030 ;
        RECT 1650.180 317.550 1650.320 324.710 ;
        RECT 1650.120 317.230 1650.380 317.550 ;
        RECT 1649.660 268.950 1649.920 269.270 ;
        RECT 1649.720 228.325 1649.860 268.950 ;
        RECT 1649.650 227.955 1649.930 228.325 ;
        RECT 1650.570 227.275 1650.850 227.645 ;
        RECT 1650.640 72.750 1650.780 227.275 ;
        RECT 1649.660 72.430 1649.920 72.750 ;
        RECT 1650.580 72.430 1650.840 72.750 ;
        RECT 1649.720 48.010 1649.860 72.430 ;
        RECT 1649.720 47.870 1650.320 48.010 ;
        RECT 1650.180 47.590 1650.320 47.870 ;
        RECT 984.040 47.270 984.300 47.590 ;
        RECT 1650.120 47.270 1650.380 47.590 ;
        RECT 984.100 2.400 984.240 47.270 ;
        RECT 983.890 -4.800 984.450 2.400 ;
      LAYER via2 ;
        RECT 1651.030 676.120 1651.310 676.400 ;
        RECT 1649.650 675.440 1649.930 675.720 ;
        RECT 1649.650 228.000 1649.930 228.280 ;
        RECT 1650.570 227.320 1650.850 227.600 ;
      LAYER met3 ;
        RECT 1651.005 676.410 1651.335 676.425 ;
        RECT 1649.870 676.110 1651.335 676.410 ;
        RECT 1649.870 675.745 1650.170 676.110 ;
        RECT 1651.005 676.095 1651.335 676.110 ;
        RECT 1649.625 675.430 1650.170 675.745 ;
        RECT 1649.625 675.415 1649.955 675.430 ;
        RECT 1649.625 228.290 1649.955 228.305 ;
        RECT 1649.625 227.975 1650.170 228.290 ;
        RECT 1649.870 227.610 1650.170 227.975 ;
        RECT 1650.545 227.610 1650.875 227.625 ;
        RECT 1649.870 227.310 1650.875 227.610 ;
        RECT 1650.545 227.295 1650.875 227.310 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1484.030 1678.140 1484.350 1678.200 ;
        RECT 1487.710 1678.140 1488.030 1678.200 ;
        RECT 1484.030 1678.000 1488.030 1678.140 ;
        RECT 1484.030 1677.940 1484.350 1678.000 ;
        RECT 1487.710 1677.940 1488.030 1678.000 ;
        RECT 662.930 44.780 663.250 44.840 ;
        RECT 1484.030 44.780 1484.350 44.840 ;
        RECT 662.930 44.640 1484.350 44.780 ;
        RECT 662.930 44.580 663.250 44.640 ;
        RECT 1484.030 44.580 1484.350 44.640 ;
      LAYER via ;
        RECT 1484.060 1677.940 1484.320 1678.200 ;
        RECT 1487.740 1677.940 1488.000 1678.200 ;
        RECT 662.960 44.580 663.220 44.840 ;
        RECT 1484.060 44.580 1484.320 44.840 ;
      LAYER met2 ;
        RECT 1489.500 1700.410 1489.780 1702.400 ;
        RECT 1487.800 1700.270 1489.780 1700.410 ;
        RECT 1487.800 1678.230 1487.940 1700.270 ;
        RECT 1489.500 1700.000 1489.780 1700.270 ;
        RECT 1484.060 1677.910 1484.320 1678.230 ;
        RECT 1487.740 1677.910 1488.000 1678.230 ;
        RECT 1484.120 44.870 1484.260 1677.910 ;
        RECT 662.960 44.550 663.220 44.870 ;
        RECT 1484.060 44.550 1484.320 44.870 ;
        RECT 663.020 2.400 663.160 44.550 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1001.950 47.840 1002.270 47.900 ;
        RECT 1662.970 47.840 1663.290 47.900 ;
        RECT 1001.950 47.700 1663.290 47.840 ;
        RECT 1001.950 47.640 1002.270 47.700 ;
        RECT 1662.970 47.640 1663.290 47.700 ;
      LAYER via ;
        RECT 1001.980 47.640 1002.240 47.900 ;
        RECT 1663.000 47.640 1663.260 47.900 ;
      LAYER met2 ;
        RECT 1664.300 1700.410 1664.580 1702.400 ;
        RECT 1663.060 1700.270 1664.580 1700.410 ;
        RECT 1663.060 47.930 1663.200 1700.270 ;
        RECT 1664.300 1700.000 1664.580 1700.270 ;
        RECT 1001.980 47.610 1002.240 47.930 ;
        RECT 1663.000 47.610 1663.260 47.930 ;
        RECT 1002.040 2.400 1002.180 47.610 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1669.870 1658.080 1670.190 1658.140 ;
        RECT 1671.250 1658.080 1671.570 1658.140 ;
        RECT 1669.870 1657.940 1671.570 1658.080 ;
        RECT 1669.870 1657.880 1670.190 1657.940 ;
        RECT 1671.250 1657.880 1671.570 1657.940 ;
        RECT 1019.430 48.180 1019.750 48.240 ;
        RECT 1669.870 48.180 1670.190 48.240 ;
        RECT 1019.430 48.040 1670.190 48.180 ;
        RECT 1019.430 47.980 1019.750 48.040 ;
        RECT 1669.870 47.980 1670.190 48.040 ;
      LAYER via ;
        RECT 1669.900 1657.880 1670.160 1658.140 ;
        RECT 1671.280 1657.880 1671.540 1658.140 ;
        RECT 1019.460 47.980 1019.720 48.240 ;
        RECT 1669.900 47.980 1670.160 48.240 ;
      LAYER met2 ;
        RECT 1673.500 1700.410 1673.780 1702.400 ;
        RECT 1671.340 1700.270 1673.780 1700.410 ;
        RECT 1671.340 1658.170 1671.480 1700.270 ;
        RECT 1673.500 1700.000 1673.780 1700.270 ;
        RECT 1669.900 1657.850 1670.160 1658.170 ;
        RECT 1671.280 1657.850 1671.540 1658.170 ;
        RECT 1669.960 48.270 1670.100 1657.850 ;
        RECT 1019.460 47.950 1019.720 48.270 ;
        RECT 1669.900 47.950 1670.160 48.270 ;
        RECT 1019.520 2.400 1019.660 47.950 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1676.770 1678.140 1677.090 1678.200 ;
        RECT 1680.910 1678.140 1681.230 1678.200 ;
        RECT 1676.770 1678.000 1681.230 1678.140 ;
        RECT 1676.770 1677.940 1677.090 1678.000 ;
        RECT 1680.910 1677.940 1681.230 1678.000 ;
        RECT 1037.370 44.100 1037.690 44.160 ;
        RECT 1676.770 44.100 1677.090 44.160 ;
        RECT 1037.370 43.960 1677.090 44.100 ;
        RECT 1037.370 43.900 1037.690 43.960 ;
        RECT 1676.770 43.900 1677.090 43.960 ;
      LAYER via ;
        RECT 1676.800 1677.940 1677.060 1678.200 ;
        RECT 1680.940 1677.940 1681.200 1678.200 ;
        RECT 1037.400 43.900 1037.660 44.160 ;
        RECT 1676.800 43.900 1677.060 44.160 ;
      LAYER met2 ;
        RECT 1682.240 1700.410 1682.520 1702.400 ;
        RECT 1681.000 1700.270 1682.520 1700.410 ;
        RECT 1681.000 1678.230 1681.140 1700.270 ;
        RECT 1682.240 1700.000 1682.520 1700.270 ;
        RECT 1676.800 1677.910 1677.060 1678.230 ;
        RECT 1680.940 1677.910 1681.200 1678.230 ;
        RECT 1676.860 44.190 1677.000 1677.910 ;
        RECT 1037.400 43.870 1037.660 44.190 ;
        RECT 1676.800 43.870 1677.060 44.190 ;
        RECT 1037.460 2.400 1037.600 43.870 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1054.850 44.440 1055.170 44.500 ;
        RECT 1691.030 44.440 1691.350 44.500 ;
        RECT 1054.850 44.300 1691.350 44.440 ;
        RECT 1054.850 44.240 1055.170 44.300 ;
        RECT 1691.030 44.240 1691.350 44.300 ;
      LAYER via ;
        RECT 1054.880 44.240 1055.140 44.500 ;
        RECT 1691.060 44.240 1691.320 44.500 ;
      LAYER met2 ;
        RECT 1691.440 1700.410 1691.720 1702.400 ;
        RECT 1691.120 1700.270 1691.720 1700.410 ;
        RECT 1691.120 44.530 1691.260 1700.270 ;
        RECT 1691.440 1700.000 1691.720 1700.270 ;
        RECT 1054.880 44.210 1055.140 44.530 ;
        RECT 1691.060 44.210 1691.320 44.530 ;
        RECT 1054.940 17.410 1055.080 44.210 ;
        RECT 1054.940 17.270 1055.540 17.410 ;
        RECT 1055.400 2.400 1055.540 17.270 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1073.250 43.760 1073.570 43.820 ;
        RECT 1698.850 43.760 1699.170 43.820 ;
        RECT 1073.250 43.620 1699.170 43.760 ;
        RECT 1073.250 43.560 1073.570 43.620 ;
        RECT 1698.850 43.560 1699.170 43.620 ;
      LAYER via ;
        RECT 1073.280 43.560 1073.540 43.820 ;
        RECT 1698.880 43.560 1699.140 43.820 ;
      LAYER met2 ;
        RECT 1700.640 1700.410 1700.920 1702.400 ;
        RECT 1698.940 1700.270 1700.920 1700.410 ;
        RECT 1698.940 43.850 1699.080 1700.270 ;
        RECT 1700.640 1700.000 1700.920 1700.270 ;
        RECT 1073.280 43.530 1073.540 43.850 ;
        RECT 1698.880 43.530 1699.140 43.850 ;
        RECT 1073.340 2.400 1073.480 43.530 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1704.370 1673.040 1704.690 1673.100 ;
        RECT 1708.510 1673.040 1708.830 1673.100 ;
        RECT 1704.370 1672.900 1708.830 1673.040 ;
        RECT 1704.370 1672.840 1704.690 1672.900 ;
        RECT 1708.510 1672.840 1708.830 1672.900 ;
        RECT 1090.730 43.080 1091.050 43.140 ;
        RECT 1704.370 43.080 1704.690 43.140 ;
        RECT 1090.730 42.940 1704.690 43.080 ;
        RECT 1090.730 42.880 1091.050 42.940 ;
        RECT 1704.370 42.880 1704.690 42.940 ;
      LAYER via ;
        RECT 1704.400 1672.840 1704.660 1673.100 ;
        RECT 1708.540 1672.840 1708.800 1673.100 ;
        RECT 1090.760 42.880 1091.020 43.140 ;
        RECT 1704.400 42.880 1704.660 43.140 ;
      LAYER met2 ;
        RECT 1709.840 1700.410 1710.120 1702.400 ;
        RECT 1708.600 1700.270 1710.120 1700.410 ;
        RECT 1708.600 1673.130 1708.740 1700.270 ;
        RECT 1709.840 1700.000 1710.120 1700.270 ;
        RECT 1704.400 1672.810 1704.660 1673.130 ;
        RECT 1708.540 1672.810 1708.800 1673.130 ;
        RECT 1704.460 43.170 1704.600 1672.810 ;
        RECT 1090.760 42.850 1091.020 43.170 ;
        RECT 1704.400 42.850 1704.660 43.170 ;
        RECT 1090.820 2.400 1090.960 42.850 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1108.670 43.420 1108.990 43.480 ;
        RECT 1718.630 43.420 1718.950 43.480 ;
        RECT 1108.670 43.280 1718.950 43.420 ;
        RECT 1108.670 43.220 1108.990 43.280 ;
        RECT 1718.630 43.220 1718.950 43.280 ;
      LAYER via ;
        RECT 1108.700 43.220 1108.960 43.480 ;
        RECT 1718.660 43.220 1718.920 43.480 ;
      LAYER met2 ;
        RECT 1719.040 1700.410 1719.320 1702.400 ;
        RECT 1718.720 1700.270 1719.320 1700.410 ;
        RECT 1718.720 43.510 1718.860 1700.270 ;
        RECT 1719.040 1700.000 1719.320 1700.270 ;
        RECT 1108.700 43.190 1108.960 43.510 ;
        RECT 1718.660 43.190 1718.920 43.510 ;
        RECT 1108.760 2.400 1108.900 43.190 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1126.610 42.740 1126.930 42.800 ;
        RECT 1725.990 42.740 1726.310 42.800 ;
        RECT 1126.610 42.600 1726.310 42.740 ;
        RECT 1126.610 42.540 1126.930 42.600 ;
        RECT 1725.990 42.540 1726.310 42.600 ;
      LAYER via ;
        RECT 1126.640 42.540 1126.900 42.800 ;
        RECT 1726.020 42.540 1726.280 42.800 ;
      LAYER met2 ;
        RECT 1728.240 1700.410 1728.520 1702.400 ;
        RECT 1726.080 1700.270 1728.520 1700.410 ;
        RECT 1726.080 42.830 1726.220 1700.270 ;
        RECT 1728.240 1700.000 1728.520 1700.270 ;
        RECT 1126.640 42.510 1126.900 42.830 ;
        RECT 1726.020 42.510 1726.280 42.830 ;
        RECT 1126.700 2.400 1126.840 42.510 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1732.965 1545.725 1733.135 1559.155 ;
        RECT 1732.965 1449.165 1733.135 1497.275 ;
        RECT 1732.965 1352.605 1733.135 1400.715 ;
        RECT 1732.965 1256.045 1733.135 1304.155 ;
        RECT 1732.965 579.785 1733.135 627.895 ;
        RECT 1732.965 483.225 1733.135 531.335 ;
        RECT 1732.965 403.665 1733.135 434.775 ;
        RECT 1732.045 113.645 1732.215 137.955 ;
        RECT 1732.505 42.245 1732.675 48.195 ;
      LAYER mcon ;
        RECT 1732.965 1558.985 1733.135 1559.155 ;
        RECT 1732.965 1497.105 1733.135 1497.275 ;
        RECT 1732.965 1400.545 1733.135 1400.715 ;
        RECT 1732.965 1303.985 1733.135 1304.155 ;
        RECT 1732.965 627.725 1733.135 627.895 ;
        RECT 1732.965 531.165 1733.135 531.335 ;
        RECT 1732.965 434.605 1733.135 434.775 ;
        RECT 1732.045 137.785 1732.215 137.955 ;
        RECT 1732.505 48.025 1732.675 48.195 ;
      LAYER met1 ;
        RECT 1732.890 1559.140 1733.210 1559.200 ;
        RECT 1732.695 1559.000 1733.210 1559.140 ;
        RECT 1732.890 1558.940 1733.210 1559.000 ;
        RECT 1732.890 1545.880 1733.210 1545.940 ;
        RECT 1732.695 1545.740 1733.210 1545.880 ;
        RECT 1732.890 1545.680 1733.210 1545.740 ;
        RECT 1732.890 1497.260 1733.210 1497.320 ;
        RECT 1732.695 1497.120 1733.210 1497.260 ;
        RECT 1732.890 1497.060 1733.210 1497.120 ;
        RECT 1732.890 1449.320 1733.210 1449.380 ;
        RECT 1732.695 1449.180 1733.210 1449.320 ;
        RECT 1732.890 1449.120 1733.210 1449.180 ;
        RECT 1732.890 1400.700 1733.210 1400.760 ;
        RECT 1732.695 1400.560 1733.210 1400.700 ;
        RECT 1732.890 1400.500 1733.210 1400.560 ;
        RECT 1732.890 1352.760 1733.210 1352.820 ;
        RECT 1732.695 1352.620 1733.210 1352.760 ;
        RECT 1732.890 1352.560 1733.210 1352.620 ;
        RECT 1732.890 1304.140 1733.210 1304.200 ;
        RECT 1732.695 1304.000 1733.210 1304.140 ;
        RECT 1732.890 1303.940 1733.210 1304.000 ;
        RECT 1732.890 1256.200 1733.210 1256.260 ;
        RECT 1732.695 1256.060 1733.210 1256.200 ;
        RECT 1732.890 1256.000 1733.210 1256.060 ;
        RECT 1732.890 1159.300 1733.210 1159.360 ;
        RECT 1733.810 1159.300 1734.130 1159.360 ;
        RECT 1732.890 1159.160 1734.130 1159.300 ;
        RECT 1732.890 1159.100 1733.210 1159.160 ;
        RECT 1733.810 1159.100 1734.130 1159.160 ;
        RECT 1732.890 1062.740 1733.210 1062.800 ;
        RECT 1733.810 1062.740 1734.130 1062.800 ;
        RECT 1732.890 1062.600 1734.130 1062.740 ;
        RECT 1732.890 1062.540 1733.210 1062.600 ;
        RECT 1733.810 1062.540 1734.130 1062.600 ;
        RECT 1732.890 966.180 1733.210 966.240 ;
        RECT 1733.810 966.180 1734.130 966.240 ;
        RECT 1732.890 966.040 1734.130 966.180 ;
        RECT 1732.890 965.980 1733.210 966.040 ;
        RECT 1733.810 965.980 1734.130 966.040 ;
        RECT 1732.890 869.620 1733.210 869.680 ;
        RECT 1733.810 869.620 1734.130 869.680 ;
        RECT 1732.890 869.480 1734.130 869.620 ;
        RECT 1732.890 869.420 1733.210 869.480 ;
        RECT 1733.810 869.420 1734.130 869.480 ;
        RECT 1732.890 821.000 1733.210 821.060 ;
        RECT 1733.810 821.000 1734.130 821.060 ;
        RECT 1732.890 820.860 1734.130 821.000 ;
        RECT 1732.890 820.800 1733.210 820.860 ;
        RECT 1733.810 820.800 1734.130 820.860 ;
        RECT 1732.890 724.440 1733.210 724.500 ;
        RECT 1733.810 724.440 1734.130 724.500 ;
        RECT 1732.890 724.300 1734.130 724.440 ;
        RECT 1732.890 724.240 1733.210 724.300 ;
        RECT 1733.810 724.240 1734.130 724.300 ;
        RECT 1732.890 627.880 1733.210 627.940 ;
        RECT 1732.695 627.740 1733.210 627.880 ;
        RECT 1732.890 627.680 1733.210 627.740 ;
        RECT 1732.890 579.940 1733.210 580.000 ;
        RECT 1732.695 579.800 1733.210 579.940 ;
        RECT 1732.890 579.740 1733.210 579.800 ;
        RECT 1732.890 531.320 1733.210 531.380 ;
        RECT 1732.695 531.180 1733.210 531.320 ;
        RECT 1732.890 531.120 1733.210 531.180 ;
        RECT 1732.890 483.380 1733.210 483.440 ;
        RECT 1732.695 483.240 1733.210 483.380 ;
        RECT 1732.890 483.180 1733.210 483.240 ;
        RECT 1732.890 434.760 1733.210 434.820 ;
        RECT 1732.695 434.620 1733.210 434.760 ;
        RECT 1732.890 434.560 1733.210 434.620 ;
        RECT 1732.430 403.820 1732.750 403.880 ;
        RECT 1732.905 403.820 1733.195 403.865 ;
        RECT 1732.430 403.680 1733.195 403.820 ;
        RECT 1732.430 403.620 1732.750 403.680 ;
        RECT 1732.905 403.635 1733.195 403.680 ;
        RECT 1732.430 379.340 1732.750 379.400 ;
        RECT 1732.890 379.340 1733.210 379.400 ;
        RECT 1732.430 379.200 1733.210 379.340 ;
        RECT 1732.430 379.140 1732.750 379.200 ;
        RECT 1732.890 379.140 1733.210 379.200 ;
        RECT 1732.890 159.020 1733.210 159.080 ;
        RECT 1732.520 158.880 1733.210 159.020 ;
        RECT 1732.520 158.740 1732.660 158.880 ;
        RECT 1732.890 158.820 1733.210 158.880 ;
        RECT 1732.430 158.480 1732.750 158.740 ;
        RECT 1731.985 137.940 1732.275 137.985 ;
        RECT 1732.430 137.940 1732.750 138.000 ;
        RECT 1731.985 137.800 1732.750 137.940 ;
        RECT 1731.985 137.755 1732.275 137.800 ;
        RECT 1732.430 137.740 1732.750 137.800 ;
        RECT 1731.985 113.800 1732.275 113.845 ;
        RECT 1732.430 113.800 1732.750 113.860 ;
        RECT 1731.985 113.660 1732.750 113.800 ;
        RECT 1731.985 113.615 1732.275 113.660 ;
        RECT 1732.430 113.600 1732.750 113.660 ;
        RECT 1732.430 48.180 1732.750 48.240 ;
        RECT 1732.235 48.040 1732.750 48.180 ;
        RECT 1732.430 47.980 1732.750 48.040 ;
        RECT 1144.550 42.400 1144.870 42.460 ;
        RECT 1732.445 42.400 1732.735 42.445 ;
        RECT 1144.550 42.260 1732.735 42.400 ;
        RECT 1144.550 42.200 1144.870 42.260 ;
        RECT 1732.445 42.215 1732.735 42.260 ;
      LAYER via ;
        RECT 1732.920 1558.940 1733.180 1559.200 ;
        RECT 1732.920 1545.680 1733.180 1545.940 ;
        RECT 1732.920 1497.060 1733.180 1497.320 ;
        RECT 1732.920 1449.120 1733.180 1449.380 ;
        RECT 1732.920 1400.500 1733.180 1400.760 ;
        RECT 1732.920 1352.560 1733.180 1352.820 ;
        RECT 1732.920 1303.940 1733.180 1304.200 ;
        RECT 1732.920 1256.000 1733.180 1256.260 ;
        RECT 1732.920 1159.100 1733.180 1159.360 ;
        RECT 1733.840 1159.100 1734.100 1159.360 ;
        RECT 1732.920 1062.540 1733.180 1062.800 ;
        RECT 1733.840 1062.540 1734.100 1062.800 ;
        RECT 1732.920 965.980 1733.180 966.240 ;
        RECT 1733.840 965.980 1734.100 966.240 ;
        RECT 1732.920 869.420 1733.180 869.680 ;
        RECT 1733.840 869.420 1734.100 869.680 ;
        RECT 1732.920 820.800 1733.180 821.060 ;
        RECT 1733.840 820.800 1734.100 821.060 ;
        RECT 1732.920 724.240 1733.180 724.500 ;
        RECT 1733.840 724.240 1734.100 724.500 ;
        RECT 1732.920 627.680 1733.180 627.940 ;
        RECT 1732.920 579.740 1733.180 580.000 ;
        RECT 1732.920 531.120 1733.180 531.380 ;
        RECT 1732.920 483.180 1733.180 483.440 ;
        RECT 1732.920 434.560 1733.180 434.820 ;
        RECT 1732.460 403.620 1732.720 403.880 ;
        RECT 1732.460 379.140 1732.720 379.400 ;
        RECT 1732.920 379.140 1733.180 379.400 ;
        RECT 1732.920 158.820 1733.180 159.080 ;
        RECT 1732.460 158.480 1732.720 158.740 ;
        RECT 1732.460 137.740 1732.720 138.000 ;
        RECT 1732.460 113.600 1732.720 113.860 ;
        RECT 1732.460 47.980 1732.720 48.240 ;
        RECT 1144.580 42.200 1144.840 42.460 ;
      LAYER met2 ;
        RECT 1737.440 1700.410 1737.720 1702.400 ;
        RECT 1735.280 1700.270 1737.720 1700.410 ;
        RECT 1735.280 1678.650 1735.420 1700.270 ;
        RECT 1737.440 1700.000 1737.720 1700.270 ;
        RECT 1732.980 1678.510 1735.420 1678.650 ;
        RECT 1732.980 1559.230 1733.120 1678.510 ;
        RECT 1732.920 1558.910 1733.180 1559.230 ;
        RECT 1732.920 1545.650 1733.180 1545.970 ;
        RECT 1732.980 1497.350 1733.120 1545.650 ;
        RECT 1732.920 1497.030 1733.180 1497.350 ;
        RECT 1732.920 1449.090 1733.180 1449.410 ;
        RECT 1732.980 1400.790 1733.120 1449.090 ;
        RECT 1732.920 1400.470 1733.180 1400.790 ;
        RECT 1732.920 1352.530 1733.180 1352.850 ;
        RECT 1732.980 1304.230 1733.120 1352.530 ;
        RECT 1732.920 1303.910 1733.180 1304.230 ;
        RECT 1732.920 1255.970 1733.180 1256.290 ;
        RECT 1732.980 1207.525 1733.120 1255.970 ;
        RECT 1732.910 1207.155 1733.190 1207.525 ;
        RECT 1733.830 1207.155 1734.110 1207.525 ;
        RECT 1733.900 1159.390 1734.040 1207.155 ;
        RECT 1732.920 1159.070 1733.180 1159.390 ;
        RECT 1733.840 1159.070 1734.100 1159.390 ;
        RECT 1732.980 1110.965 1733.120 1159.070 ;
        RECT 1732.910 1110.595 1733.190 1110.965 ;
        RECT 1733.830 1110.595 1734.110 1110.965 ;
        RECT 1733.900 1062.830 1734.040 1110.595 ;
        RECT 1732.920 1062.510 1733.180 1062.830 ;
        RECT 1733.840 1062.510 1734.100 1062.830 ;
        RECT 1732.980 1014.405 1733.120 1062.510 ;
        RECT 1732.910 1014.035 1733.190 1014.405 ;
        RECT 1733.830 1014.035 1734.110 1014.405 ;
        RECT 1733.900 966.270 1734.040 1014.035 ;
        RECT 1732.920 965.950 1733.180 966.270 ;
        RECT 1733.840 965.950 1734.100 966.270 ;
        RECT 1732.980 917.845 1733.120 965.950 ;
        RECT 1732.910 917.475 1733.190 917.845 ;
        RECT 1733.830 917.475 1734.110 917.845 ;
        RECT 1733.900 869.710 1734.040 917.475 ;
        RECT 1732.920 869.390 1733.180 869.710 ;
        RECT 1733.840 869.390 1734.100 869.710 ;
        RECT 1732.980 821.090 1733.120 869.390 ;
        RECT 1732.920 820.770 1733.180 821.090 ;
        RECT 1733.840 820.770 1734.100 821.090 ;
        RECT 1733.900 773.005 1734.040 820.770 ;
        RECT 1732.910 772.635 1733.190 773.005 ;
        RECT 1733.830 772.635 1734.110 773.005 ;
        RECT 1732.980 724.530 1733.120 772.635 ;
        RECT 1732.920 724.210 1733.180 724.530 ;
        RECT 1733.840 724.210 1734.100 724.530 ;
        RECT 1733.900 676.445 1734.040 724.210 ;
        RECT 1732.910 676.075 1733.190 676.445 ;
        RECT 1733.830 676.075 1734.110 676.445 ;
        RECT 1732.980 627.970 1733.120 676.075 ;
        RECT 1732.920 627.650 1733.180 627.970 ;
        RECT 1732.920 579.710 1733.180 580.030 ;
        RECT 1732.980 531.410 1733.120 579.710 ;
        RECT 1732.920 531.090 1733.180 531.410 ;
        RECT 1732.920 483.150 1733.180 483.470 ;
        RECT 1732.980 434.850 1733.120 483.150 ;
        RECT 1732.920 434.530 1733.180 434.850 ;
        RECT 1732.460 403.590 1732.720 403.910 ;
        RECT 1732.520 379.850 1732.660 403.590 ;
        RECT 1732.520 379.710 1733.120 379.850 ;
        RECT 1732.980 379.430 1733.120 379.710 ;
        RECT 1732.460 379.110 1732.720 379.430 ;
        RECT 1732.920 379.110 1733.180 379.430 ;
        RECT 1732.520 331.570 1732.660 379.110 ;
        RECT 1732.520 331.430 1733.120 331.570 ;
        RECT 1732.980 159.110 1733.120 331.430 ;
        RECT 1732.920 158.790 1733.180 159.110 ;
        RECT 1732.460 158.450 1732.720 158.770 ;
        RECT 1732.520 138.030 1732.660 158.450 ;
        RECT 1732.460 137.710 1732.720 138.030 ;
        RECT 1732.460 113.570 1732.720 113.890 ;
        RECT 1732.520 48.270 1732.660 113.570 ;
        RECT 1732.460 47.950 1732.720 48.270 ;
        RECT 1144.580 42.170 1144.840 42.490 ;
        RECT 1144.640 2.400 1144.780 42.170 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
      LAYER via2 ;
        RECT 1732.910 1207.200 1733.190 1207.480 ;
        RECT 1733.830 1207.200 1734.110 1207.480 ;
        RECT 1732.910 1110.640 1733.190 1110.920 ;
        RECT 1733.830 1110.640 1734.110 1110.920 ;
        RECT 1732.910 1014.080 1733.190 1014.360 ;
        RECT 1733.830 1014.080 1734.110 1014.360 ;
        RECT 1732.910 917.520 1733.190 917.800 ;
        RECT 1733.830 917.520 1734.110 917.800 ;
        RECT 1732.910 772.680 1733.190 772.960 ;
        RECT 1733.830 772.680 1734.110 772.960 ;
        RECT 1732.910 676.120 1733.190 676.400 ;
        RECT 1733.830 676.120 1734.110 676.400 ;
      LAYER met3 ;
        RECT 1732.885 1207.490 1733.215 1207.505 ;
        RECT 1733.805 1207.490 1734.135 1207.505 ;
        RECT 1732.885 1207.190 1734.135 1207.490 ;
        RECT 1732.885 1207.175 1733.215 1207.190 ;
        RECT 1733.805 1207.175 1734.135 1207.190 ;
        RECT 1732.885 1110.930 1733.215 1110.945 ;
        RECT 1733.805 1110.930 1734.135 1110.945 ;
        RECT 1732.885 1110.630 1734.135 1110.930 ;
        RECT 1732.885 1110.615 1733.215 1110.630 ;
        RECT 1733.805 1110.615 1734.135 1110.630 ;
        RECT 1732.885 1014.370 1733.215 1014.385 ;
        RECT 1733.805 1014.370 1734.135 1014.385 ;
        RECT 1732.885 1014.070 1734.135 1014.370 ;
        RECT 1732.885 1014.055 1733.215 1014.070 ;
        RECT 1733.805 1014.055 1734.135 1014.070 ;
        RECT 1732.885 917.810 1733.215 917.825 ;
        RECT 1733.805 917.810 1734.135 917.825 ;
        RECT 1732.885 917.510 1734.135 917.810 ;
        RECT 1732.885 917.495 1733.215 917.510 ;
        RECT 1733.805 917.495 1734.135 917.510 ;
        RECT 1732.885 772.970 1733.215 772.985 ;
        RECT 1733.805 772.970 1734.135 772.985 ;
        RECT 1732.885 772.670 1734.135 772.970 ;
        RECT 1732.885 772.655 1733.215 772.670 ;
        RECT 1733.805 772.655 1734.135 772.670 ;
        RECT 1732.885 676.410 1733.215 676.425 ;
        RECT 1733.805 676.410 1734.135 676.425 ;
        RECT 1732.885 676.110 1734.135 676.410 ;
        RECT 1732.885 676.095 1733.215 676.110 ;
        RECT 1733.805 676.095 1734.135 676.110 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1162.490 42.060 1162.810 42.120 ;
        RECT 1746.230 42.060 1746.550 42.120 ;
        RECT 1162.490 41.920 1746.550 42.060 ;
        RECT 1162.490 41.860 1162.810 41.920 ;
        RECT 1746.230 41.860 1746.550 41.920 ;
      LAYER via ;
        RECT 1162.520 41.860 1162.780 42.120 ;
        RECT 1746.260 41.860 1746.520 42.120 ;
      LAYER met2 ;
        RECT 1746.640 1700.410 1746.920 1702.400 ;
        RECT 1746.320 1700.270 1746.920 1700.410 ;
        RECT 1746.320 42.150 1746.460 1700.270 ;
        RECT 1746.640 1700.000 1746.920 1700.270 ;
        RECT 1162.520 41.830 1162.780 42.150 ;
        RECT 1746.260 41.830 1746.520 42.150 ;
        RECT 1162.580 2.400 1162.720 41.830 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1498.700 1700.410 1498.980 1702.400 ;
        RECT 1497.920 1700.270 1498.980 1700.410 ;
        RECT 1497.920 44.725 1498.060 1700.270 ;
        RECT 1498.700 1700.000 1498.980 1700.270 ;
        RECT 680.430 44.355 680.710 44.725 ;
        RECT 1497.850 44.355 1498.130 44.725 ;
        RECT 680.500 2.400 680.640 44.355 ;
        RECT 680.290 -4.800 680.850 2.400 ;
      LAYER via2 ;
        RECT 680.430 44.400 680.710 44.680 ;
        RECT 1497.850 44.400 1498.130 44.680 ;
      LAYER met3 ;
        RECT 680.405 44.690 680.735 44.705 ;
        RECT 1497.825 44.690 1498.155 44.705 ;
        RECT 680.405 44.390 1498.155 44.690 ;
        RECT 680.405 44.375 680.735 44.390 ;
        RECT 1497.825 44.375 1498.155 44.390 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 41.720 1180.290 41.780 ;
        RECT 1753.590 41.720 1753.910 41.780 ;
        RECT 1179.970 41.580 1753.910 41.720 ;
        RECT 1179.970 41.520 1180.290 41.580 ;
        RECT 1753.590 41.520 1753.910 41.580 ;
      LAYER via ;
        RECT 1180.000 41.520 1180.260 41.780 ;
        RECT 1753.620 41.520 1753.880 41.780 ;
      LAYER met2 ;
        RECT 1755.840 1700.410 1756.120 1702.400 ;
        RECT 1753.680 1700.270 1756.120 1700.410 ;
        RECT 1753.680 41.810 1753.820 1700.270 ;
        RECT 1755.840 1700.000 1756.120 1700.270 ;
        RECT 1180.000 41.490 1180.260 41.810 ;
        RECT 1753.620 41.490 1753.880 41.810 ;
        RECT 1180.060 2.400 1180.200 41.490 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1760.105 1151.665 1760.275 1173.255 ;
        RECT 1760.105 772.565 1760.275 814.215 ;
        RECT 1760.105 269.025 1760.275 290.615 ;
      LAYER mcon ;
        RECT 1760.105 1173.085 1760.275 1173.255 ;
        RECT 1760.105 814.045 1760.275 814.215 ;
        RECT 1760.105 290.445 1760.275 290.615 ;
      LAYER met1 ;
        RECT 1760.030 1593.620 1760.350 1593.880 ;
        RECT 1760.120 1593.480 1760.260 1593.620 ;
        RECT 1760.490 1593.480 1760.810 1593.540 ;
        RECT 1760.120 1593.340 1760.810 1593.480 ;
        RECT 1760.490 1593.280 1760.810 1593.340 ;
        RECT 1760.490 1490.460 1760.810 1490.520 ;
        RECT 1760.490 1490.320 1761.180 1490.460 ;
        RECT 1760.490 1490.260 1760.810 1490.320 ;
        RECT 1761.040 1490.180 1761.180 1490.320 ;
        RECT 1760.950 1489.920 1761.270 1490.180 ;
        RECT 1760.030 1435.380 1760.350 1435.440 ;
        RECT 1760.490 1435.380 1760.810 1435.440 ;
        RECT 1760.030 1435.240 1760.810 1435.380 ;
        RECT 1760.030 1435.180 1760.350 1435.240 ;
        RECT 1760.490 1435.180 1760.810 1435.240 ;
        RECT 1760.030 1401.040 1760.350 1401.100 ;
        RECT 1760.030 1400.900 1760.720 1401.040 ;
        RECT 1760.030 1400.840 1760.350 1400.900 ;
        RECT 1760.580 1400.760 1760.720 1400.900 ;
        RECT 1760.490 1400.500 1760.810 1400.760 ;
        RECT 1760.030 1317.400 1760.350 1317.460 ;
        RECT 1761.410 1317.400 1761.730 1317.460 ;
        RECT 1760.030 1317.260 1761.730 1317.400 ;
        RECT 1760.030 1317.200 1760.350 1317.260 ;
        RECT 1761.410 1317.200 1761.730 1317.260 ;
        RECT 1760.030 1173.240 1760.350 1173.300 ;
        RECT 1759.835 1173.100 1760.350 1173.240 ;
        RECT 1760.030 1173.040 1760.350 1173.100 ;
        RECT 1760.045 1151.820 1760.335 1151.865 ;
        RECT 1760.950 1151.820 1761.270 1151.880 ;
        RECT 1760.045 1151.680 1761.270 1151.820 ;
        RECT 1760.045 1151.635 1760.335 1151.680 ;
        RECT 1760.950 1151.620 1761.270 1151.680 ;
        RECT 1760.030 1104.220 1760.350 1104.280 ;
        RECT 1760.950 1104.220 1761.270 1104.280 ;
        RECT 1760.030 1104.080 1761.270 1104.220 ;
        RECT 1760.030 1104.020 1760.350 1104.080 ;
        RECT 1760.950 1104.020 1761.270 1104.080 ;
        RECT 1760.030 1062.740 1760.350 1062.800 ;
        RECT 1760.490 1062.740 1760.810 1062.800 ;
        RECT 1760.030 1062.600 1760.810 1062.740 ;
        RECT 1760.030 1062.540 1760.350 1062.600 ;
        RECT 1760.490 1062.540 1760.810 1062.600 ;
        RECT 1760.030 1014.460 1760.350 1014.520 ;
        RECT 1760.490 1014.460 1760.810 1014.520 ;
        RECT 1760.030 1014.320 1760.810 1014.460 ;
        RECT 1760.030 1014.260 1760.350 1014.320 ;
        RECT 1760.490 1014.260 1760.810 1014.320 ;
        RECT 1760.490 932.180 1760.810 932.240 ;
        RECT 1760.120 932.040 1760.810 932.180 ;
        RECT 1760.120 931.560 1760.260 932.040 ;
        RECT 1760.490 931.980 1760.810 932.040 ;
        RECT 1760.030 931.300 1760.350 931.560 ;
        RECT 1760.030 869.620 1760.350 869.680 ;
        RECT 1760.490 869.620 1760.810 869.680 ;
        RECT 1760.030 869.480 1760.810 869.620 ;
        RECT 1760.030 869.420 1760.350 869.480 ;
        RECT 1760.490 869.420 1760.810 869.480 ;
        RECT 1760.030 814.200 1760.350 814.260 ;
        RECT 1759.835 814.060 1760.350 814.200 ;
        RECT 1760.030 814.000 1760.350 814.060 ;
        RECT 1760.030 772.720 1760.350 772.780 ;
        RECT 1759.835 772.580 1760.350 772.720 ;
        RECT 1760.030 772.520 1760.350 772.580 ;
        RECT 1759.110 748.580 1759.430 748.640 ;
        RECT 1760.030 748.580 1760.350 748.640 ;
        RECT 1759.110 748.440 1760.350 748.580 ;
        RECT 1759.110 748.380 1759.430 748.440 ;
        RECT 1760.030 748.380 1760.350 748.440 ;
        RECT 1760.030 724.440 1760.350 724.500 ;
        RECT 1760.950 724.440 1761.270 724.500 ;
        RECT 1760.030 724.300 1761.270 724.440 ;
        RECT 1760.030 724.240 1760.350 724.300 ;
        RECT 1760.950 724.240 1761.270 724.300 ;
        RECT 1760.490 676.160 1760.810 676.220 ;
        RECT 1760.950 676.160 1761.270 676.220 ;
        RECT 1760.490 676.020 1761.270 676.160 ;
        RECT 1760.490 675.960 1760.810 676.020 ;
        RECT 1760.950 675.960 1761.270 676.020 ;
        RECT 1760.030 627.880 1760.350 627.940 ;
        RECT 1760.950 627.880 1761.270 627.940 ;
        RECT 1760.030 627.740 1761.270 627.880 ;
        RECT 1760.030 627.680 1760.350 627.740 ;
        RECT 1760.950 627.680 1761.270 627.740 ;
        RECT 1760.030 531.320 1760.350 531.380 ;
        RECT 1760.950 531.320 1761.270 531.380 ;
        RECT 1760.030 531.180 1761.270 531.320 ;
        RECT 1760.030 531.120 1760.350 531.180 ;
        RECT 1760.950 531.120 1761.270 531.180 ;
        RECT 1760.030 434.560 1760.350 434.820 ;
        RECT 1760.120 434.420 1760.260 434.560 ;
        RECT 1760.490 434.420 1760.810 434.480 ;
        RECT 1760.120 434.280 1760.810 434.420 ;
        RECT 1760.490 434.220 1760.810 434.280 ;
        RECT 1760.030 290.600 1760.350 290.660 ;
        RECT 1759.835 290.460 1760.350 290.600 ;
        RECT 1760.030 290.400 1760.350 290.460 ;
        RECT 1760.030 269.180 1760.350 269.240 ;
        RECT 1759.835 269.040 1760.350 269.180 ;
        RECT 1760.030 268.980 1760.350 269.040 ;
        RECT 1760.030 227.700 1760.350 227.760 ;
        RECT 1761.870 227.700 1762.190 227.760 ;
        RECT 1760.030 227.560 1762.190 227.700 ;
        RECT 1760.030 227.500 1760.350 227.560 ;
        RECT 1761.870 227.500 1762.190 227.560 ;
        RECT 1760.030 96.800 1760.350 96.860 ;
        RECT 1760.950 96.800 1761.270 96.860 ;
        RECT 1760.030 96.660 1761.270 96.800 ;
        RECT 1760.030 96.600 1760.350 96.660 ;
        RECT 1760.950 96.600 1761.270 96.660 ;
        RECT 1200.210 70.280 1200.530 70.340 ;
        RECT 1760.030 70.280 1760.350 70.340 ;
        RECT 1200.210 70.140 1760.350 70.280 ;
        RECT 1200.210 70.080 1200.530 70.140 ;
        RECT 1760.030 70.080 1760.350 70.140 ;
        RECT 1197.910 18.260 1198.230 18.320 ;
        RECT 1200.210 18.260 1200.530 18.320 ;
        RECT 1197.910 18.120 1200.530 18.260 ;
        RECT 1197.910 18.060 1198.230 18.120 ;
        RECT 1200.210 18.060 1200.530 18.120 ;
      LAYER via ;
        RECT 1760.060 1593.620 1760.320 1593.880 ;
        RECT 1760.520 1593.280 1760.780 1593.540 ;
        RECT 1760.520 1490.260 1760.780 1490.520 ;
        RECT 1760.980 1489.920 1761.240 1490.180 ;
        RECT 1760.060 1435.180 1760.320 1435.440 ;
        RECT 1760.520 1435.180 1760.780 1435.440 ;
        RECT 1760.060 1400.840 1760.320 1401.100 ;
        RECT 1760.520 1400.500 1760.780 1400.760 ;
        RECT 1760.060 1317.200 1760.320 1317.460 ;
        RECT 1761.440 1317.200 1761.700 1317.460 ;
        RECT 1760.060 1173.040 1760.320 1173.300 ;
        RECT 1760.980 1151.620 1761.240 1151.880 ;
        RECT 1760.060 1104.020 1760.320 1104.280 ;
        RECT 1760.980 1104.020 1761.240 1104.280 ;
        RECT 1760.060 1062.540 1760.320 1062.800 ;
        RECT 1760.520 1062.540 1760.780 1062.800 ;
        RECT 1760.060 1014.260 1760.320 1014.520 ;
        RECT 1760.520 1014.260 1760.780 1014.520 ;
        RECT 1760.520 931.980 1760.780 932.240 ;
        RECT 1760.060 931.300 1760.320 931.560 ;
        RECT 1760.060 869.420 1760.320 869.680 ;
        RECT 1760.520 869.420 1760.780 869.680 ;
        RECT 1760.060 814.000 1760.320 814.260 ;
        RECT 1760.060 772.520 1760.320 772.780 ;
        RECT 1759.140 748.380 1759.400 748.640 ;
        RECT 1760.060 748.380 1760.320 748.640 ;
        RECT 1760.060 724.240 1760.320 724.500 ;
        RECT 1760.980 724.240 1761.240 724.500 ;
        RECT 1760.520 675.960 1760.780 676.220 ;
        RECT 1760.980 675.960 1761.240 676.220 ;
        RECT 1760.060 627.680 1760.320 627.940 ;
        RECT 1760.980 627.680 1761.240 627.940 ;
        RECT 1760.060 531.120 1760.320 531.380 ;
        RECT 1760.980 531.120 1761.240 531.380 ;
        RECT 1760.060 434.560 1760.320 434.820 ;
        RECT 1760.520 434.220 1760.780 434.480 ;
        RECT 1760.060 290.400 1760.320 290.660 ;
        RECT 1760.060 268.980 1760.320 269.240 ;
        RECT 1760.060 227.500 1760.320 227.760 ;
        RECT 1761.900 227.500 1762.160 227.760 ;
        RECT 1760.060 96.600 1760.320 96.860 ;
        RECT 1760.980 96.600 1761.240 96.860 ;
        RECT 1200.240 70.080 1200.500 70.340 ;
        RECT 1760.060 70.080 1760.320 70.340 ;
        RECT 1197.940 18.060 1198.200 18.320 ;
        RECT 1200.240 18.060 1200.500 18.320 ;
      LAYER met2 ;
        RECT 1765.040 1700.410 1765.320 1702.400 ;
        RECT 1763.340 1700.270 1765.320 1700.410 ;
        RECT 1763.340 1678.140 1763.480 1700.270 ;
        RECT 1765.040 1700.000 1765.320 1700.270 ;
        RECT 1760.580 1678.000 1763.480 1678.140 ;
        RECT 1760.580 1594.330 1760.720 1678.000 ;
        RECT 1760.120 1594.190 1760.720 1594.330 ;
        RECT 1760.120 1593.910 1760.260 1594.190 ;
        RECT 1760.060 1593.590 1760.320 1593.910 ;
        RECT 1760.520 1593.250 1760.780 1593.570 ;
        RECT 1760.580 1490.550 1760.720 1593.250 ;
        RECT 1760.520 1490.230 1760.780 1490.550 ;
        RECT 1760.980 1489.890 1761.240 1490.210 ;
        RECT 1761.040 1483.490 1761.180 1489.890 ;
        RECT 1760.580 1483.350 1761.180 1483.490 ;
        RECT 1760.580 1435.470 1760.720 1483.350 ;
        RECT 1760.060 1435.150 1760.320 1435.470 ;
        RECT 1760.520 1435.150 1760.780 1435.470 ;
        RECT 1760.120 1401.130 1760.260 1435.150 ;
        RECT 1760.060 1400.810 1760.320 1401.130 ;
        RECT 1760.520 1400.470 1760.780 1400.790 ;
        RECT 1760.580 1345.565 1760.720 1400.470 ;
        RECT 1760.510 1345.195 1760.790 1345.565 ;
        RECT 1761.430 1345.195 1761.710 1345.565 ;
        RECT 1761.500 1317.490 1761.640 1345.195 ;
        RECT 1760.060 1317.170 1760.320 1317.490 ;
        RECT 1761.440 1317.170 1761.700 1317.490 ;
        RECT 1760.120 1173.330 1760.260 1317.170 ;
        RECT 1760.060 1173.010 1760.320 1173.330 ;
        RECT 1760.980 1151.590 1761.240 1151.910 ;
        RECT 1761.040 1104.310 1761.180 1151.590 ;
        RECT 1760.060 1103.990 1760.320 1104.310 ;
        RECT 1760.980 1103.990 1761.240 1104.310 ;
        RECT 1760.120 1062.830 1760.260 1103.990 ;
        RECT 1760.060 1062.510 1760.320 1062.830 ;
        RECT 1760.520 1062.510 1760.780 1062.830 ;
        RECT 1760.580 1014.550 1760.720 1062.510 ;
        RECT 1760.060 1014.405 1760.320 1014.550 ;
        RECT 1760.050 1014.035 1760.330 1014.405 ;
        RECT 1760.520 1014.230 1760.780 1014.550 ;
        RECT 1760.510 1013.355 1760.790 1013.725 ;
        RECT 1760.580 932.270 1760.720 1013.355 ;
        RECT 1760.520 931.950 1760.780 932.270 ;
        RECT 1760.060 931.270 1760.320 931.590 ;
        RECT 1760.120 869.710 1760.260 931.270 ;
        RECT 1760.060 869.390 1760.320 869.710 ;
        RECT 1760.520 869.390 1760.780 869.710 ;
        RECT 1760.580 821.285 1760.720 869.390 ;
        RECT 1760.510 820.915 1760.790 821.285 ;
        RECT 1760.050 820.235 1760.330 820.605 ;
        RECT 1760.120 814.290 1760.260 820.235 ;
        RECT 1760.060 813.970 1760.320 814.290 ;
        RECT 1760.060 772.490 1760.320 772.810 ;
        RECT 1760.120 748.670 1760.260 772.490 ;
        RECT 1759.140 748.350 1759.400 748.670 ;
        RECT 1760.060 748.350 1760.320 748.670 ;
        RECT 1759.200 724.725 1759.340 748.350 ;
        RECT 1759.130 724.355 1759.410 724.725 ;
        RECT 1760.050 724.355 1760.330 724.725 ;
        RECT 1760.060 724.210 1760.320 724.355 ;
        RECT 1760.980 724.210 1761.240 724.530 ;
        RECT 1761.040 688.570 1761.180 724.210 ;
        RECT 1760.580 688.430 1761.180 688.570 ;
        RECT 1760.580 676.250 1760.720 688.430 ;
        RECT 1760.520 675.930 1760.780 676.250 ;
        RECT 1760.980 675.930 1761.240 676.250 ;
        RECT 1761.040 628.165 1761.180 675.930 ;
        RECT 1760.050 627.795 1760.330 628.165 ;
        RECT 1760.970 627.795 1761.250 628.165 ;
        RECT 1760.060 627.650 1760.320 627.795 ;
        RECT 1760.980 627.650 1761.240 627.795 ;
        RECT 1761.040 592.010 1761.180 627.650 ;
        RECT 1760.580 591.870 1761.180 592.010 ;
        RECT 1760.580 545.770 1760.720 591.870 ;
        RECT 1760.580 545.630 1761.180 545.770 ;
        RECT 1761.040 544.410 1761.180 545.630 ;
        RECT 1760.120 544.270 1761.180 544.410 ;
        RECT 1760.120 531.410 1760.260 544.270 ;
        RECT 1760.060 531.090 1760.320 531.410 ;
        RECT 1760.980 531.090 1761.240 531.410 ;
        RECT 1761.040 495.450 1761.180 531.090 ;
        RECT 1760.580 495.310 1761.180 495.450 ;
        RECT 1760.580 435.725 1760.720 495.310 ;
        RECT 1760.510 435.355 1760.790 435.725 ;
        RECT 1760.050 434.675 1760.330 435.045 ;
        RECT 1760.060 434.530 1760.320 434.675 ;
        RECT 1760.520 434.190 1760.780 434.510 ;
        RECT 1760.580 362.170 1760.720 434.190 ;
        RECT 1760.120 362.030 1760.720 362.170 ;
        RECT 1760.120 290.690 1760.260 362.030 ;
        RECT 1760.060 290.370 1760.320 290.690 ;
        RECT 1760.060 268.950 1760.320 269.270 ;
        RECT 1760.120 227.790 1760.260 268.950 ;
        RECT 1760.060 227.470 1760.320 227.790 ;
        RECT 1761.900 227.470 1762.160 227.790 ;
        RECT 1761.960 161.570 1762.100 227.470 ;
        RECT 1760.580 161.430 1762.100 161.570 ;
        RECT 1760.580 121.450 1760.720 161.430 ;
        RECT 1760.580 121.310 1761.180 121.450 ;
        RECT 1761.040 96.890 1761.180 121.310 ;
        RECT 1760.060 96.570 1760.320 96.890 ;
        RECT 1760.980 96.570 1761.240 96.890 ;
        RECT 1760.120 70.370 1760.260 96.570 ;
        RECT 1200.240 70.050 1200.500 70.370 ;
        RECT 1760.060 70.050 1760.320 70.370 ;
        RECT 1200.300 18.350 1200.440 70.050 ;
        RECT 1197.940 18.030 1198.200 18.350 ;
        RECT 1200.240 18.030 1200.500 18.350 ;
        RECT 1198.000 2.400 1198.140 18.030 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
      LAYER via2 ;
        RECT 1760.510 1345.240 1760.790 1345.520 ;
        RECT 1761.430 1345.240 1761.710 1345.520 ;
        RECT 1760.050 1014.080 1760.330 1014.360 ;
        RECT 1760.510 1013.400 1760.790 1013.680 ;
        RECT 1760.510 820.960 1760.790 821.240 ;
        RECT 1760.050 820.280 1760.330 820.560 ;
        RECT 1759.130 724.400 1759.410 724.680 ;
        RECT 1760.050 724.400 1760.330 724.680 ;
        RECT 1760.050 627.840 1760.330 628.120 ;
        RECT 1760.970 627.840 1761.250 628.120 ;
        RECT 1760.510 435.400 1760.790 435.680 ;
        RECT 1760.050 434.720 1760.330 435.000 ;
      LAYER met3 ;
        RECT 1760.485 1345.530 1760.815 1345.545 ;
        RECT 1761.405 1345.530 1761.735 1345.545 ;
        RECT 1760.485 1345.230 1761.735 1345.530 ;
        RECT 1760.485 1345.215 1760.815 1345.230 ;
        RECT 1761.405 1345.215 1761.735 1345.230 ;
        RECT 1760.025 1014.370 1760.355 1014.385 ;
        RECT 1760.025 1014.055 1760.570 1014.370 ;
        RECT 1760.270 1013.705 1760.570 1014.055 ;
        RECT 1760.270 1013.390 1760.815 1013.705 ;
        RECT 1760.485 1013.375 1760.815 1013.390 ;
        RECT 1760.485 821.250 1760.815 821.265 ;
        RECT 1759.350 820.950 1760.815 821.250 ;
        RECT 1759.350 820.570 1759.650 820.950 ;
        RECT 1760.485 820.935 1760.815 820.950 ;
        RECT 1760.025 820.570 1760.355 820.585 ;
        RECT 1759.350 820.270 1760.355 820.570 ;
        RECT 1760.025 820.255 1760.355 820.270 ;
        RECT 1759.105 724.690 1759.435 724.705 ;
        RECT 1760.025 724.690 1760.355 724.705 ;
        RECT 1759.105 724.390 1760.355 724.690 ;
        RECT 1759.105 724.375 1759.435 724.390 ;
        RECT 1760.025 724.375 1760.355 724.390 ;
        RECT 1760.025 628.130 1760.355 628.145 ;
        RECT 1760.945 628.130 1761.275 628.145 ;
        RECT 1760.025 627.830 1761.275 628.130 ;
        RECT 1760.025 627.815 1760.355 627.830 ;
        RECT 1760.945 627.815 1761.275 627.830 ;
        RECT 1760.485 435.690 1760.815 435.705 ;
        RECT 1760.270 435.375 1760.815 435.690 ;
        RECT 1760.270 435.025 1760.570 435.375 ;
        RECT 1760.025 434.710 1760.570 435.025 ;
        RECT 1760.025 434.695 1760.355 434.710 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1220.910 72.320 1221.230 72.380 ;
        RECT 1773.830 72.320 1774.150 72.380 ;
        RECT 1220.910 72.180 1774.150 72.320 ;
        RECT 1220.910 72.120 1221.230 72.180 ;
        RECT 1773.830 72.120 1774.150 72.180 ;
        RECT 1215.850 18.260 1216.170 18.320 ;
        RECT 1220.910 18.260 1221.230 18.320 ;
        RECT 1215.850 18.120 1221.230 18.260 ;
        RECT 1215.850 18.060 1216.170 18.120 ;
        RECT 1220.910 18.060 1221.230 18.120 ;
      LAYER via ;
        RECT 1220.940 72.120 1221.200 72.380 ;
        RECT 1773.860 72.120 1774.120 72.380 ;
        RECT 1215.880 18.060 1216.140 18.320 ;
        RECT 1220.940 18.060 1221.200 18.320 ;
      LAYER met2 ;
        RECT 1774.240 1700.410 1774.520 1702.400 ;
        RECT 1773.920 1700.270 1774.520 1700.410 ;
        RECT 1773.920 72.410 1774.060 1700.270 ;
        RECT 1774.240 1700.000 1774.520 1700.270 ;
        RECT 1220.940 72.090 1221.200 72.410 ;
        RECT 1773.860 72.090 1774.120 72.410 ;
        RECT 1221.000 18.350 1221.140 72.090 ;
        RECT 1215.880 18.030 1216.140 18.350 ;
        RECT 1220.940 18.030 1221.200 18.350 ;
        RECT 1215.940 2.400 1216.080 18.030 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 49.540 1234.110 49.600 ;
        RECT 1781.190 49.540 1781.510 49.600 ;
        RECT 1233.790 49.400 1781.510 49.540 ;
        RECT 1233.790 49.340 1234.110 49.400 ;
        RECT 1781.190 49.340 1781.510 49.400 ;
      LAYER via ;
        RECT 1233.820 49.340 1234.080 49.600 ;
        RECT 1781.220 49.340 1781.480 49.600 ;
      LAYER met2 ;
        RECT 1783.440 1700.410 1783.720 1702.400 ;
        RECT 1781.280 1700.270 1783.720 1700.410 ;
        RECT 1781.280 49.630 1781.420 1700.270 ;
        RECT 1783.440 1700.000 1783.720 1700.270 ;
        RECT 1233.820 49.310 1234.080 49.630 ;
        RECT 1781.220 49.310 1781.480 49.630 ;
        RECT 1233.880 2.400 1234.020 49.310 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1788.165 1629.025 1788.335 1676.455 ;
        RECT 1787.705 917.745 1787.875 932.195 ;
        RECT 1788.165 772.905 1788.335 821.015 ;
        RECT 1787.705 324.445 1787.875 372.555 ;
      LAYER mcon ;
        RECT 1788.165 1676.285 1788.335 1676.455 ;
        RECT 1787.705 932.025 1787.875 932.195 ;
        RECT 1788.165 820.845 1788.335 821.015 ;
        RECT 1787.705 372.385 1787.875 372.555 ;
      LAYER met1 ;
        RECT 1788.090 1678.140 1788.410 1678.200 ;
        RECT 1791.310 1678.140 1791.630 1678.200 ;
        RECT 1788.090 1678.000 1791.630 1678.140 ;
        RECT 1788.090 1677.940 1788.410 1678.000 ;
        RECT 1791.310 1677.940 1791.630 1678.000 ;
        RECT 1788.090 1676.440 1788.410 1676.500 ;
        RECT 1787.895 1676.300 1788.410 1676.440 ;
        RECT 1788.090 1676.240 1788.410 1676.300 ;
        RECT 1788.090 1629.180 1788.410 1629.240 ;
        RECT 1787.895 1629.040 1788.410 1629.180 ;
        RECT 1788.090 1628.980 1788.410 1629.040 ;
        RECT 1787.630 1580.220 1787.950 1580.280 ;
        RECT 1789.010 1580.220 1789.330 1580.280 ;
        RECT 1787.630 1580.080 1789.330 1580.220 ;
        RECT 1787.630 1580.020 1787.950 1580.080 ;
        RECT 1789.010 1580.020 1789.330 1580.080 ;
        RECT 1787.630 1531.940 1787.950 1532.000 ;
        RECT 1788.090 1531.940 1788.410 1532.000 ;
        RECT 1787.630 1531.800 1788.410 1531.940 ;
        RECT 1787.630 1531.740 1787.950 1531.800 ;
        RECT 1788.090 1531.740 1788.410 1531.800 ;
        RECT 1788.090 1459.520 1788.410 1459.580 ;
        RECT 1789.010 1459.520 1789.330 1459.580 ;
        RECT 1788.090 1459.380 1789.330 1459.520 ;
        RECT 1788.090 1459.320 1788.410 1459.380 ;
        RECT 1789.010 1459.320 1789.330 1459.380 ;
        RECT 1788.090 1366.500 1788.410 1366.760 ;
        RECT 1788.180 1366.080 1788.320 1366.500 ;
        RECT 1788.090 1365.820 1788.410 1366.080 ;
        RECT 1788.090 1269.940 1788.410 1270.200 ;
        RECT 1788.180 1269.520 1788.320 1269.940 ;
        RECT 1788.090 1269.260 1788.410 1269.520 ;
        RECT 1788.550 1173.240 1788.870 1173.300 ;
        RECT 1788.180 1173.100 1788.870 1173.240 ;
        RECT 1788.180 1172.960 1788.320 1173.100 ;
        RECT 1788.550 1173.040 1788.870 1173.100 ;
        RECT 1788.090 1172.700 1788.410 1172.960 ;
        RECT 1788.550 1076.680 1788.870 1076.740 ;
        RECT 1788.180 1076.540 1788.870 1076.680 ;
        RECT 1788.180 1076.400 1788.320 1076.540 ;
        RECT 1788.550 1076.480 1788.870 1076.540 ;
        RECT 1788.090 1076.140 1788.410 1076.400 ;
        RECT 1787.645 932.180 1787.935 932.225 ;
        RECT 1788.090 932.180 1788.410 932.240 ;
        RECT 1787.645 932.040 1788.410 932.180 ;
        RECT 1787.645 931.995 1787.935 932.040 ;
        RECT 1788.090 931.980 1788.410 932.040 ;
        RECT 1787.630 917.900 1787.950 917.960 ;
        RECT 1787.435 917.760 1787.950 917.900 ;
        RECT 1787.630 917.700 1787.950 917.760 ;
        RECT 1788.090 821.000 1788.410 821.060 ;
        RECT 1787.895 820.860 1788.410 821.000 ;
        RECT 1788.090 820.800 1788.410 820.860 ;
        RECT 1788.090 773.060 1788.410 773.120 ;
        RECT 1787.895 772.920 1788.410 773.060 ;
        RECT 1788.090 772.860 1788.410 772.920 ;
        RECT 1788.090 724.780 1788.410 724.840 ;
        RECT 1788.550 724.780 1788.870 724.840 ;
        RECT 1788.090 724.640 1788.870 724.780 ;
        RECT 1788.090 724.580 1788.410 724.640 ;
        RECT 1788.550 724.580 1788.870 724.640 ;
        RECT 1787.630 717.640 1787.950 717.700 ;
        RECT 1788.090 717.640 1788.410 717.700 ;
        RECT 1787.630 717.500 1788.410 717.640 ;
        RECT 1787.630 717.440 1787.950 717.500 ;
        RECT 1788.090 717.440 1788.410 717.500 ;
        RECT 1788.090 627.880 1788.410 627.940 ;
        RECT 1788.550 627.880 1788.870 627.940 ;
        RECT 1788.090 627.740 1788.870 627.880 ;
        RECT 1788.090 627.680 1788.410 627.740 ;
        RECT 1788.550 627.680 1788.870 627.740 ;
        RECT 1788.090 434.760 1788.410 434.820 ;
        RECT 1789.010 434.760 1789.330 434.820 ;
        RECT 1788.090 434.620 1789.330 434.760 ;
        RECT 1788.090 434.560 1788.410 434.620 ;
        RECT 1789.010 434.560 1789.330 434.620 ;
        RECT 1787.645 372.540 1787.935 372.585 ;
        RECT 1788.090 372.540 1788.410 372.600 ;
        RECT 1787.645 372.400 1788.410 372.540 ;
        RECT 1787.645 372.355 1787.935 372.400 ;
        RECT 1788.090 372.340 1788.410 372.400 ;
        RECT 1787.630 324.600 1787.950 324.660 ;
        RECT 1787.435 324.460 1787.950 324.600 ;
        RECT 1787.630 324.400 1787.950 324.460 ;
        RECT 1787.630 96.800 1787.950 96.860 ;
        RECT 1788.090 96.800 1788.410 96.860 ;
        RECT 1787.630 96.660 1788.410 96.800 ;
        RECT 1787.630 96.600 1787.950 96.660 ;
        RECT 1788.090 96.600 1788.410 96.660 ;
        RECT 1251.730 49.200 1252.050 49.260 ;
        RECT 1788.090 49.200 1788.410 49.260 ;
        RECT 1251.730 49.060 1788.410 49.200 ;
        RECT 1251.730 49.000 1252.050 49.060 ;
        RECT 1788.090 49.000 1788.410 49.060 ;
      LAYER via ;
        RECT 1788.120 1677.940 1788.380 1678.200 ;
        RECT 1791.340 1677.940 1791.600 1678.200 ;
        RECT 1788.120 1676.240 1788.380 1676.500 ;
        RECT 1788.120 1628.980 1788.380 1629.240 ;
        RECT 1787.660 1580.020 1787.920 1580.280 ;
        RECT 1789.040 1580.020 1789.300 1580.280 ;
        RECT 1787.660 1531.740 1787.920 1532.000 ;
        RECT 1788.120 1531.740 1788.380 1532.000 ;
        RECT 1788.120 1459.320 1788.380 1459.580 ;
        RECT 1789.040 1459.320 1789.300 1459.580 ;
        RECT 1788.120 1366.500 1788.380 1366.760 ;
        RECT 1788.120 1365.820 1788.380 1366.080 ;
        RECT 1788.120 1269.940 1788.380 1270.200 ;
        RECT 1788.120 1269.260 1788.380 1269.520 ;
        RECT 1788.580 1173.040 1788.840 1173.300 ;
        RECT 1788.120 1172.700 1788.380 1172.960 ;
        RECT 1788.580 1076.480 1788.840 1076.740 ;
        RECT 1788.120 1076.140 1788.380 1076.400 ;
        RECT 1788.120 931.980 1788.380 932.240 ;
        RECT 1787.660 917.700 1787.920 917.960 ;
        RECT 1788.120 820.800 1788.380 821.060 ;
        RECT 1788.120 772.860 1788.380 773.120 ;
        RECT 1788.120 724.580 1788.380 724.840 ;
        RECT 1788.580 724.580 1788.840 724.840 ;
        RECT 1787.660 717.440 1787.920 717.700 ;
        RECT 1788.120 717.440 1788.380 717.700 ;
        RECT 1788.120 627.680 1788.380 627.940 ;
        RECT 1788.580 627.680 1788.840 627.940 ;
        RECT 1788.120 434.560 1788.380 434.820 ;
        RECT 1789.040 434.560 1789.300 434.820 ;
        RECT 1788.120 372.340 1788.380 372.600 ;
        RECT 1787.660 324.400 1787.920 324.660 ;
        RECT 1787.660 96.600 1787.920 96.860 ;
        RECT 1788.120 96.600 1788.380 96.860 ;
        RECT 1251.760 49.000 1252.020 49.260 ;
        RECT 1788.120 49.000 1788.380 49.260 ;
      LAYER met2 ;
        RECT 1792.640 1700.410 1792.920 1702.400 ;
        RECT 1791.400 1700.270 1792.920 1700.410 ;
        RECT 1791.400 1678.230 1791.540 1700.270 ;
        RECT 1792.640 1700.000 1792.920 1700.270 ;
        RECT 1788.120 1677.910 1788.380 1678.230 ;
        RECT 1791.340 1677.910 1791.600 1678.230 ;
        RECT 1788.180 1676.530 1788.320 1677.910 ;
        RECT 1788.120 1676.210 1788.380 1676.530 ;
        RECT 1788.120 1628.950 1788.380 1629.270 ;
        RECT 1788.180 1628.445 1788.320 1628.950 ;
        RECT 1788.110 1628.075 1788.390 1628.445 ;
        RECT 1789.030 1628.075 1789.310 1628.445 ;
        RECT 1787.720 1580.310 1787.860 1580.465 ;
        RECT 1789.100 1580.310 1789.240 1628.075 ;
        RECT 1787.660 1580.050 1787.920 1580.310 ;
        RECT 1787.660 1579.990 1788.320 1580.050 ;
        RECT 1789.040 1579.990 1789.300 1580.310 ;
        RECT 1787.720 1579.910 1788.320 1579.990 ;
        RECT 1788.180 1532.030 1788.320 1579.910 ;
        RECT 1787.660 1531.710 1787.920 1532.030 ;
        RECT 1788.120 1531.710 1788.380 1532.030 ;
        RECT 1787.720 1514.770 1787.860 1531.710 ;
        RECT 1787.720 1514.630 1788.780 1514.770 ;
        RECT 1788.640 1491.765 1788.780 1514.630 ;
        RECT 1788.570 1491.395 1788.850 1491.765 ;
        RECT 1788.110 1490.715 1788.390 1491.085 ;
        RECT 1788.180 1483.605 1788.320 1490.715 ;
        RECT 1788.110 1483.235 1788.390 1483.605 ;
        RECT 1789.030 1483.235 1789.310 1483.605 ;
        RECT 1789.100 1459.610 1789.240 1483.235 ;
        RECT 1788.120 1459.290 1788.380 1459.610 ;
        RECT 1789.040 1459.290 1789.300 1459.610 ;
        RECT 1788.180 1366.790 1788.320 1459.290 ;
        RECT 1788.120 1366.470 1788.380 1366.790 ;
        RECT 1788.120 1365.790 1788.380 1366.110 ;
        RECT 1788.180 1270.230 1788.320 1365.790 ;
        RECT 1788.120 1269.910 1788.380 1270.230 ;
        RECT 1788.120 1269.230 1788.380 1269.550 ;
        RECT 1788.180 1207.410 1788.320 1269.230 ;
        RECT 1788.180 1207.270 1788.780 1207.410 ;
        RECT 1788.640 1173.330 1788.780 1207.270 ;
        RECT 1788.580 1173.010 1788.840 1173.330 ;
        RECT 1788.120 1172.670 1788.380 1172.990 ;
        RECT 1788.180 1110.850 1788.320 1172.670 ;
        RECT 1788.180 1110.710 1788.780 1110.850 ;
        RECT 1788.640 1076.770 1788.780 1110.710 ;
        RECT 1788.580 1076.450 1788.840 1076.770 ;
        RECT 1788.120 1076.110 1788.380 1076.430 ;
        RECT 1788.180 980.290 1788.320 1076.110 ;
        RECT 1787.720 980.150 1788.320 980.290 ;
        RECT 1787.720 979.610 1787.860 980.150 ;
        RECT 1787.720 979.470 1788.320 979.610 ;
        RECT 1788.180 932.270 1788.320 979.470 ;
        RECT 1788.120 931.950 1788.380 932.270 ;
        RECT 1787.720 917.990 1787.860 918.145 ;
        RECT 1787.660 917.730 1787.920 917.990 ;
        RECT 1787.660 917.670 1788.320 917.730 ;
        RECT 1787.720 917.590 1788.320 917.670 ;
        RECT 1788.180 821.090 1788.320 917.590 ;
        RECT 1788.120 820.770 1788.380 821.090 ;
        RECT 1788.120 772.830 1788.380 773.150 ;
        RECT 1788.180 738.210 1788.320 772.830 ;
        RECT 1788.180 738.070 1788.780 738.210 ;
        RECT 1788.640 724.870 1788.780 738.070 ;
        RECT 1788.120 724.610 1788.380 724.870 ;
        RECT 1787.720 724.550 1788.380 724.610 ;
        RECT 1788.580 724.550 1788.840 724.870 ;
        RECT 1787.720 724.470 1788.320 724.550 ;
        RECT 1787.720 717.730 1787.860 724.470 ;
        RECT 1787.660 717.410 1787.920 717.730 ;
        RECT 1788.120 717.410 1788.380 717.730 ;
        RECT 1788.180 627.970 1788.320 717.410 ;
        RECT 1788.120 627.650 1788.380 627.970 ;
        RECT 1788.580 627.650 1788.840 627.970 ;
        RECT 1788.640 579.885 1788.780 627.650 ;
        RECT 1788.570 579.515 1788.850 579.885 ;
        RECT 1789.030 578.835 1789.310 579.205 ;
        RECT 1789.100 531.605 1789.240 578.835 ;
        RECT 1788.110 531.235 1788.390 531.605 ;
        RECT 1789.030 531.235 1789.310 531.605 ;
        RECT 1788.180 434.850 1788.320 531.235 ;
        RECT 1788.120 434.530 1788.380 434.850 ;
        RECT 1789.040 434.530 1789.300 434.850 ;
        RECT 1789.100 386.765 1789.240 434.530 ;
        RECT 1788.110 386.395 1788.390 386.765 ;
        RECT 1789.030 386.395 1789.310 386.765 ;
        RECT 1788.180 372.630 1788.320 386.395 ;
        RECT 1788.120 372.310 1788.380 372.630 ;
        RECT 1787.660 324.370 1787.920 324.690 ;
        RECT 1787.720 234.330 1787.860 324.370 ;
        RECT 1787.720 234.190 1788.320 234.330 ;
        RECT 1788.180 169.050 1788.320 234.190 ;
        RECT 1787.720 168.910 1788.320 169.050 ;
        RECT 1787.720 96.890 1787.860 168.910 ;
        RECT 1787.660 96.570 1787.920 96.890 ;
        RECT 1788.120 96.570 1788.380 96.890 ;
        RECT 1788.180 49.290 1788.320 96.570 ;
        RECT 1251.760 48.970 1252.020 49.290 ;
        RECT 1788.120 48.970 1788.380 49.290 ;
        RECT 1251.820 2.400 1251.960 48.970 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
      LAYER via2 ;
        RECT 1788.110 1628.120 1788.390 1628.400 ;
        RECT 1789.030 1628.120 1789.310 1628.400 ;
        RECT 1788.570 1491.440 1788.850 1491.720 ;
        RECT 1788.110 1490.760 1788.390 1491.040 ;
        RECT 1788.110 1483.280 1788.390 1483.560 ;
        RECT 1789.030 1483.280 1789.310 1483.560 ;
        RECT 1788.570 579.560 1788.850 579.840 ;
        RECT 1789.030 578.880 1789.310 579.160 ;
        RECT 1788.110 531.280 1788.390 531.560 ;
        RECT 1789.030 531.280 1789.310 531.560 ;
        RECT 1788.110 386.440 1788.390 386.720 ;
        RECT 1789.030 386.440 1789.310 386.720 ;
      LAYER met3 ;
        RECT 1788.085 1628.410 1788.415 1628.425 ;
        RECT 1789.005 1628.410 1789.335 1628.425 ;
        RECT 1788.085 1628.110 1789.335 1628.410 ;
        RECT 1788.085 1628.095 1788.415 1628.110 ;
        RECT 1789.005 1628.095 1789.335 1628.110 ;
        RECT 1788.545 1491.730 1788.875 1491.745 ;
        RECT 1788.545 1491.415 1789.090 1491.730 ;
        RECT 1788.085 1491.050 1788.415 1491.065 ;
        RECT 1788.790 1491.050 1789.090 1491.415 ;
        RECT 1788.085 1490.750 1789.090 1491.050 ;
        RECT 1788.085 1490.735 1788.415 1490.750 ;
        RECT 1788.085 1483.570 1788.415 1483.585 ;
        RECT 1789.005 1483.570 1789.335 1483.585 ;
        RECT 1788.085 1483.270 1789.335 1483.570 ;
        RECT 1788.085 1483.255 1788.415 1483.270 ;
        RECT 1789.005 1483.255 1789.335 1483.270 ;
        RECT 1788.545 579.850 1788.875 579.865 ;
        RECT 1787.870 579.550 1788.875 579.850 ;
        RECT 1787.870 579.170 1788.170 579.550 ;
        RECT 1788.545 579.535 1788.875 579.550 ;
        RECT 1789.005 579.170 1789.335 579.185 ;
        RECT 1787.870 578.870 1789.335 579.170 ;
        RECT 1789.005 578.855 1789.335 578.870 ;
        RECT 1788.085 531.570 1788.415 531.585 ;
        RECT 1789.005 531.570 1789.335 531.585 ;
        RECT 1788.085 531.270 1789.335 531.570 ;
        RECT 1788.085 531.255 1788.415 531.270 ;
        RECT 1789.005 531.255 1789.335 531.270 ;
        RECT 1788.085 386.730 1788.415 386.745 ;
        RECT 1789.005 386.730 1789.335 386.745 ;
        RECT 1788.085 386.430 1789.335 386.730 ;
        RECT 1788.085 386.415 1788.415 386.430 ;
        RECT 1789.005 386.415 1789.335 386.430 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 48.860 1269.530 48.920 ;
        RECT 1801.430 48.860 1801.750 48.920 ;
        RECT 1269.210 48.720 1801.750 48.860 ;
        RECT 1269.210 48.660 1269.530 48.720 ;
        RECT 1801.430 48.660 1801.750 48.720 ;
      LAYER via ;
        RECT 1269.240 48.660 1269.500 48.920 ;
        RECT 1801.460 48.660 1801.720 48.920 ;
      LAYER met2 ;
        RECT 1801.840 1700.410 1802.120 1702.400 ;
        RECT 1801.520 1700.270 1802.120 1700.410 ;
        RECT 1801.520 48.950 1801.660 1700.270 ;
        RECT 1801.840 1700.000 1802.120 1700.270 ;
        RECT 1269.240 48.630 1269.500 48.950 ;
        RECT 1801.460 48.630 1801.720 48.950 ;
        RECT 1269.300 2.400 1269.440 48.630 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1287.150 48.520 1287.470 48.580 ;
        RECT 1808.790 48.520 1809.110 48.580 ;
        RECT 1287.150 48.380 1809.110 48.520 ;
        RECT 1287.150 48.320 1287.470 48.380 ;
        RECT 1808.790 48.320 1809.110 48.380 ;
      LAYER via ;
        RECT 1287.180 48.320 1287.440 48.580 ;
        RECT 1808.820 48.320 1809.080 48.580 ;
      LAYER met2 ;
        RECT 1811.040 1700.410 1811.320 1702.400 ;
        RECT 1808.880 1700.270 1811.320 1700.410 ;
        RECT 1808.880 48.610 1809.020 1700.270 ;
        RECT 1811.040 1700.000 1811.320 1700.270 ;
        RECT 1287.180 48.290 1287.440 48.610 ;
        RECT 1808.820 48.290 1809.080 48.610 ;
        RECT 1287.240 2.400 1287.380 48.290 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1814.770 1672.020 1815.090 1672.080 ;
        RECT 1818.910 1672.020 1819.230 1672.080 ;
        RECT 1814.770 1671.880 1819.230 1672.020 ;
        RECT 1814.770 1671.820 1815.090 1671.880 ;
        RECT 1818.910 1671.820 1819.230 1671.880 ;
        RECT 1780.270 23.020 1780.590 23.080 ;
        RECT 1814.770 23.020 1815.090 23.080 ;
        RECT 1780.270 22.880 1815.090 23.020 ;
        RECT 1780.270 22.820 1780.590 22.880 ;
        RECT 1814.770 22.820 1815.090 22.880 ;
        RECT 1305.090 17.240 1305.410 17.300 ;
        RECT 1780.270 17.240 1780.590 17.300 ;
        RECT 1305.090 17.100 1780.590 17.240 ;
        RECT 1305.090 17.040 1305.410 17.100 ;
        RECT 1780.270 17.040 1780.590 17.100 ;
      LAYER via ;
        RECT 1814.800 1671.820 1815.060 1672.080 ;
        RECT 1818.940 1671.820 1819.200 1672.080 ;
        RECT 1780.300 22.820 1780.560 23.080 ;
        RECT 1814.800 22.820 1815.060 23.080 ;
        RECT 1305.120 17.040 1305.380 17.300 ;
        RECT 1780.300 17.040 1780.560 17.300 ;
      LAYER met2 ;
        RECT 1820.240 1700.410 1820.520 1702.400 ;
        RECT 1819.000 1700.270 1820.520 1700.410 ;
        RECT 1819.000 1672.110 1819.140 1700.270 ;
        RECT 1820.240 1700.000 1820.520 1700.270 ;
        RECT 1814.800 1671.790 1815.060 1672.110 ;
        RECT 1818.940 1671.790 1819.200 1672.110 ;
        RECT 1814.860 23.110 1815.000 1671.790 ;
        RECT 1780.300 22.790 1780.560 23.110 ;
        RECT 1814.800 22.790 1815.060 23.110 ;
        RECT 1780.360 17.330 1780.500 22.790 ;
        RECT 1305.120 17.010 1305.380 17.330 ;
        RECT 1780.300 17.010 1780.560 17.330 ;
        RECT 1305.180 2.400 1305.320 17.010 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1390.265 18.445 1390.435 19.975 ;
      LAYER mcon ;
        RECT 1390.265 19.805 1390.435 19.975 ;
      LAYER met1 ;
        RECT 1417.790 1688.340 1418.110 1688.400 ;
        RECT 1829.490 1688.340 1829.810 1688.400 ;
        RECT 1417.790 1688.200 1829.810 1688.340 ;
        RECT 1417.790 1688.140 1418.110 1688.200 ;
        RECT 1829.490 1688.140 1829.810 1688.200 ;
        RECT 1390.205 19.960 1390.495 20.005 ;
        RECT 1417.330 19.960 1417.650 20.020 ;
        RECT 1390.205 19.820 1417.650 19.960 ;
        RECT 1390.205 19.775 1390.495 19.820 ;
        RECT 1417.330 19.760 1417.650 19.820 ;
        RECT 1323.030 18.600 1323.350 18.660 ;
        RECT 1390.205 18.600 1390.495 18.645 ;
        RECT 1323.030 18.460 1390.495 18.600 ;
        RECT 1323.030 18.400 1323.350 18.460 ;
        RECT 1390.205 18.415 1390.495 18.460 ;
      LAYER via ;
        RECT 1417.820 1688.140 1418.080 1688.400 ;
        RECT 1829.520 1688.140 1829.780 1688.400 ;
        RECT 1417.360 19.760 1417.620 20.020 ;
        RECT 1323.060 18.400 1323.320 18.660 ;
      LAYER met2 ;
        RECT 1829.440 1700.000 1829.720 1702.400 ;
        RECT 1829.580 1688.430 1829.720 1700.000 ;
        RECT 1417.820 1688.110 1418.080 1688.430 ;
        RECT 1829.520 1688.110 1829.780 1688.430 ;
        RECT 1417.880 40.530 1418.020 1688.110 ;
        RECT 1417.420 40.390 1418.020 40.530 ;
        RECT 1417.420 20.050 1417.560 40.390 ;
        RECT 1417.360 19.730 1417.620 20.050 ;
        RECT 1323.060 18.370 1323.320 18.690 ;
        RECT 1323.120 2.400 1323.260 18.370 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1390.265 16.745 1390.435 17.935 ;
      LAYER mcon ;
        RECT 1390.265 17.765 1390.435 17.935 ;
      LAYER met1 ;
        RECT 1449.530 52.940 1449.850 53.000 ;
        RECT 1836.390 52.940 1836.710 53.000 ;
        RECT 1449.530 52.800 1836.710 52.940 ;
        RECT 1449.530 52.740 1449.850 52.800 ;
        RECT 1836.390 52.740 1836.710 52.800 ;
        RECT 1390.205 17.920 1390.495 17.965 ;
        RECT 1390.205 17.780 1438.720 17.920 ;
        RECT 1390.205 17.735 1390.495 17.780 ;
        RECT 1438.580 17.580 1438.720 17.780 ;
        RECT 1449.530 17.580 1449.850 17.640 ;
        RECT 1438.580 17.440 1449.850 17.580 ;
        RECT 1449.530 17.380 1449.850 17.440 ;
        RECT 1340.510 16.900 1340.830 16.960 ;
        RECT 1390.205 16.900 1390.495 16.945 ;
        RECT 1340.510 16.760 1390.495 16.900 ;
        RECT 1340.510 16.700 1340.830 16.760 ;
        RECT 1390.205 16.715 1390.495 16.760 ;
      LAYER via ;
        RECT 1449.560 52.740 1449.820 53.000 ;
        RECT 1836.420 52.740 1836.680 53.000 ;
        RECT 1449.560 17.380 1449.820 17.640 ;
        RECT 1340.540 16.700 1340.800 16.960 ;
      LAYER met2 ;
        RECT 1838.640 1700.410 1838.920 1702.400 ;
        RECT 1836.480 1700.270 1838.920 1700.410 ;
        RECT 1836.480 53.030 1836.620 1700.270 ;
        RECT 1838.640 1700.000 1838.920 1700.270 ;
        RECT 1449.560 52.710 1449.820 53.030 ;
        RECT 1836.420 52.710 1836.680 53.030 ;
        RECT 1449.620 17.670 1449.760 52.710 ;
        RECT 1449.560 17.350 1449.820 17.670 ;
        RECT 1340.540 16.670 1340.800 16.990 ;
        RECT 1340.600 2.400 1340.740 16.670 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 54.640 703.730 54.700 ;
        RECT 1505.190 54.640 1505.510 54.700 ;
        RECT 703.410 54.500 1505.510 54.640 ;
        RECT 703.410 54.440 703.730 54.500 ;
        RECT 1505.190 54.440 1505.510 54.500 ;
        RECT 698.350 2.960 698.670 3.020 ;
        RECT 703.410 2.960 703.730 3.020 ;
        RECT 698.350 2.820 703.730 2.960 ;
        RECT 698.350 2.760 698.670 2.820 ;
        RECT 703.410 2.760 703.730 2.820 ;
      LAYER via ;
        RECT 703.440 54.440 703.700 54.700 ;
        RECT 1505.220 54.440 1505.480 54.700 ;
        RECT 698.380 2.760 698.640 3.020 ;
        RECT 703.440 2.760 703.700 3.020 ;
      LAYER met2 ;
        RECT 1507.900 1700.410 1508.180 1702.400 ;
        RECT 1505.280 1700.270 1508.180 1700.410 ;
        RECT 1505.280 54.730 1505.420 1700.270 ;
        RECT 1507.900 1700.000 1508.180 1700.270 ;
        RECT 703.440 54.410 703.700 54.730 ;
        RECT 1505.220 54.410 1505.480 54.730 ;
        RECT 703.500 3.050 703.640 54.410 ;
        RECT 698.380 2.730 698.640 3.050 ;
        RECT 703.440 2.730 703.700 3.050 ;
        RECT 698.440 2.400 698.580 2.730 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1816.225 1686.995 1816.395 1688.695 ;
        RECT 1817.145 1686.995 1817.315 1687.335 ;
        RECT 1816.225 1686.825 1817.315 1686.995 ;
        RECT 1389.805 18.275 1389.975 19.975 ;
        RECT 1390.725 18.275 1390.895 18.615 ;
        RECT 1389.805 18.105 1390.895 18.275 ;
      LAYER mcon ;
        RECT 1816.225 1688.525 1816.395 1688.695 ;
        RECT 1817.145 1687.165 1817.315 1687.335 ;
        RECT 1389.805 19.805 1389.975 19.975 ;
        RECT 1390.725 18.445 1390.895 18.615 ;
      LAYER met1 ;
        RECT 1438.490 1688.680 1438.810 1688.740 ;
        RECT 1816.165 1688.680 1816.455 1688.725 ;
        RECT 1438.490 1688.540 1816.455 1688.680 ;
        RECT 1438.490 1688.480 1438.810 1688.540 ;
        RECT 1816.165 1688.495 1816.455 1688.540 ;
        RECT 1817.085 1687.320 1817.375 1687.365 ;
        RECT 1847.890 1687.320 1848.210 1687.380 ;
        RECT 1817.085 1687.180 1848.210 1687.320 ;
        RECT 1817.085 1687.135 1817.375 1687.180 ;
        RECT 1847.890 1687.120 1848.210 1687.180 ;
        RECT 1358.450 19.960 1358.770 20.020 ;
        RECT 1389.745 19.960 1390.035 20.005 ;
        RECT 1358.450 19.820 1390.035 19.960 ;
        RECT 1358.450 19.760 1358.770 19.820 ;
        RECT 1389.745 19.775 1390.035 19.820 ;
        RECT 1390.665 18.600 1390.955 18.645 ;
        RECT 1438.490 18.600 1438.810 18.660 ;
        RECT 1390.665 18.460 1438.810 18.600 ;
        RECT 1390.665 18.415 1390.955 18.460 ;
        RECT 1438.490 18.400 1438.810 18.460 ;
      LAYER via ;
        RECT 1438.520 1688.480 1438.780 1688.740 ;
        RECT 1847.920 1687.120 1848.180 1687.380 ;
        RECT 1358.480 19.760 1358.740 20.020 ;
        RECT 1438.520 18.400 1438.780 18.660 ;
      LAYER met2 ;
        RECT 1847.840 1700.000 1848.120 1702.400 ;
        RECT 1438.520 1688.450 1438.780 1688.770 ;
        RECT 1358.480 19.730 1358.740 20.050 ;
        RECT 1358.540 2.400 1358.680 19.730 ;
        RECT 1438.580 18.690 1438.720 1688.450 ;
        RECT 1847.980 1687.410 1848.120 1700.000 ;
        RECT 1847.920 1687.090 1848.180 1687.410 ;
        RECT 1438.520 18.370 1438.780 18.690 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1383.290 1686.980 1383.610 1687.040 ;
        RECT 1857.090 1686.980 1857.410 1687.040 ;
        RECT 1383.290 1686.840 1857.410 1686.980 ;
        RECT 1383.290 1686.780 1383.610 1686.840 ;
        RECT 1857.090 1686.780 1857.410 1686.840 ;
        RECT 1376.390 20.640 1376.710 20.700 ;
        RECT 1383.290 20.640 1383.610 20.700 ;
        RECT 1376.390 20.500 1383.610 20.640 ;
        RECT 1376.390 20.440 1376.710 20.500 ;
        RECT 1383.290 20.440 1383.610 20.500 ;
      LAYER via ;
        RECT 1383.320 1686.780 1383.580 1687.040 ;
        RECT 1857.120 1686.780 1857.380 1687.040 ;
        RECT 1376.420 20.440 1376.680 20.700 ;
        RECT 1383.320 20.440 1383.580 20.700 ;
      LAYER met2 ;
        RECT 1857.040 1700.000 1857.320 1702.400 ;
        RECT 1857.180 1687.070 1857.320 1700.000 ;
        RECT 1383.320 1686.750 1383.580 1687.070 ;
        RECT 1857.120 1686.750 1857.380 1687.070 ;
        RECT 1383.380 20.730 1383.520 1686.750 ;
        RECT 1376.420 20.410 1376.680 20.730 ;
        RECT 1383.320 20.410 1383.580 20.730 ;
        RECT 1376.480 2.400 1376.620 20.410 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1816.685 1687.165 1816.855 1688.695 ;
      LAYER mcon ;
        RECT 1816.685 1688.525 1816.855 1688.695 ;
      LAYER met1 ;
        RECT 1816.625 1688.680 1816.915 1688.725 ;
        RECT 1866.290 1688.680 1866.610 1688.740 ;
        RECT 1816.625 1688.540 1866.610 1688.680 ;
        RECT 1816.625 1688.495 1816.915 1688.540 ;
        RECT 1866.290 1688.480 1866.610 1688.540 ;
        RECT 1400.310 1687.320 1400.630 1687.380 ;
        RECT 1816.625 1687.320 1816.915 1687.365 ;
        RECT 1400.310 1687.180 1816.915 1687.320 ;
        RECT 1400.310 1687.120 1400.630 1687.180 ;
        RECT 1816.625 1687.135 1816.915 1687.180 ;
        RECT 1400.310 850.720 1400.630 850.980 ;
        RECT 1400.400 849.960 1400.540 850.720 ;
        RECT 1400.310 849.700 1400.630 849.960 ;
        RECT 1394.330 20.640 1394.650 20.700 ;
        RECT 1400.310 20.640 1400.630 20.700 ;
        RECT 1394.330 20.500 1400.630 20.640 ;
        RECT 1394.330 20.440 1394.650 20.500 ;
        RECT 1400.310 20.440 1400.630 20.500 ;
      LAYER via ;
        RECT 1866.320 1688.480 1866.580 1688.740 ;
        RECT 1400.340 1687.120 1400.600 1687.380 ;
        RECT 1400.340 850.720 1400.600 850.980 ;
        RECT 1400.340 849.700 1400.600 849.960 ;
        RECT 1394.360 20.440 1394.620 20.700 ;
        RECT 1400.340 20.440 1400.600 20.700 ;
      LAYER met2 ;
        RECT 1866.240 1700.000 1866.520 1702.400 ;
        RECT 1866.380 1688.770 1866.520 1700.000 ;
        RECT 1866.320 1688.450 1866.580 1688.770 ;
        RECT 1400.340 1687.090 1400.600 1687.410 ;
        RECT 1400.400 851.010 1400.540 1687.090 ;
        RECT 1400.340 850.690 1400.600 851.010 ;
        RECT 1400.340 849.670 1400.600 849.990 ;
        RECT 1400.400 20.730 1400.540 849.670 ;
        RECT 1394.360 20.410 1394.620 20.730 ;
        RECT 1400.340 20.410 1400.600 20.730 ;
        RECT 1394.420 2.400 1394.560 20.410 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1472.990 1689.020 1473.310 1689.080 ;
        RECT 1875.490 1689.020 1875.810 1689.080 ;
        RECT 1472.990 1688.880 1875.810 1689.020 ;
        RECT 1472.990 1688.820 1473.310 1688.880 ;
        RECT 1875.490 1688.820 1875.810 1688.880 ;
        RECT 1412.270 16.900 1412.590 16.960 ;
        RECT 1472.990 16.900 1473.310 16.960 ;
        RECT 1412.270 16.760 1473.310 16.900 ;
        RECT 1412.270 16.700 1412.590 16.760 ;
        RECT 1472.990 16.700 1473.310 16.760 ;
      LAYER via ;
        RECT 1473.020 1688.820 1473.280 1689.080 ;
        RECT 1875.520 1688.820 1875.780 1689.080 ;
        RECT 1412.300 16.700 1412.560 16.960 ;
        RECT 1473.020 16.700 1473.280 16.960 ;
      LAYER met2 ;
        RECT 1875.440 1700.000 1875.720 1702.400 ;
        RECT 1875.580 1689.110 1875.720 1700.000 ;
        RECT 1473.020 1688.790 1473.280 1689.110 ;
        RECT 1875.520 1688.790 1875.780 1689.110 ;
        RECT 1473.080 16.990 1473.220 1688.790 ;
        RECT 1412.300 16.670 1412.560 16.990 ;
        RECT 1473.020 16.670 1473.280 16.990 ;
        RECT 1412.360 2.400 1412.500 16.670 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1434.810 1687.660 1435.130 1687.720 ;
        RECT 1884.690 1687.660 1885.010 1687.720 ;
        RECT 1434.810 1687.520 1885.010 1687.660 ;
        RECT 1434.810 1687.460 1435.130 1687.520 ;
        RECT 1884.690 1687.460 1885.010 1687.520 ;
        RECT 1429.750 15.880 1430.070 15.940 ;
        RECT 1434.810 15.880 1435.130 15.940 ;
        RECT 1429.750 15.740 1435.130 15.880 ;
        RECT 1429.750 15.680 1430.070 15.740 ;
        RECT 1434.810 15.680 1435.130 15.740 ;
      LAYER via ;
        RECT 1434.840 1687.460 1435.100 1687.720 ;
        RECT 1884.720 1687.460 1884.980 1687.720 ;
        RECT 1429.780 15.680 1430.040 15.940 ;
        RECT 1434.840 15.680 1435.100 15.940 ;
      LAYER met2 ;
        RECT 1884.640 1700.000 1884.920 1702.400 ;
        RECT 1884.780 1687.750 1884.920 1700.000 ;
        RECT 1434.840 1687.430 1435.100 1687.750 ;
        RECT 1884.720 1687.430 1884.980 1687.750 ;
        RECT 1434.900 15.970 1435.040 1687.430 ;
        RECT 1429.780 15.650 1430.040 15.970 ;
        RECT 1434.840 15.650 1435.100 15.970 ;
        RECT 1429.840 2.400 1429.980 15.650 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1462.945 16.405 1463.115 17.935 ;
        RECT 1510.785 16.405 1510.955 17.595 ;
      LAYER mcon ;
        RECT 1462.945 17.765 1463.115 17.935 ;
        RECT 1510.785 17.425 1510.955 17.595 ;
      LAYER met1 ;
        RECT 1447.690 17.920 1448.010 17.980 ;
        RECT 1462.885 17.920 1463.175 17.965 ;
        RECT 1447.690 17.780 1463.175 17.920 ;
        RECT 1447.690 17.720 1448.010 17.780 ;
        RECT 1462.885 17.735 1463.175 17.780 ;
        RECT 1510.725 17.580 1511.015 17.625 ;
        RECT 1892.050 17.580 1892.370 17.640 ;
        RECT 1510.725 17.440 1892.370 17.580 ;
        RECT 1510.725 17.395 1511.015 17.440 ;
        RECT 1892.050 17.380 1892.370 17.440 ;
        RECT 1462.885 16.560 1463.175 16.605 ;
        RECT 1510.725 16.560 1511.015 16.605 ;
        RECT 1462.885 16.420 1511.015 16.560 ;
        RECT 1462.885 16.375 1463.175 16.420 ;
        RECT 1510.725 16.375 1511.015 16.420 ;
      LAYER via ;
        RECT 1447.720 17.720 1447.980 17.980 ;
        RECT 1892.080 17.380 1892.340 17.640 ;
      LAYER met2 ;
        RECT 1893.840 1700.410 1894.120 1702.400 ;
        RECT 1892.140 1700.270 1894.120 1700.410 ;
        RECT 1447.720 17.690 1447.980 18.010 ;
        RECT 1447.780 2.400 1447.920 17.690 ;
        RECT 1892.140 17.670 1892.280 1700.270 ;
        RECT 1893.840 1700.000 1894.120 1700.270 ;
        RECT 1892.080 17.350 1892.340 17.670 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.310 1688.000 1469.630 1688.060 ;
        RECT 1903.090 1688.000 1903.410 1688.060 ;
        RECT 1469.310 1687.860 1903.410 1688.000 ;
        RECT 1469.310 1687.800 1469.630 1687.860 ;
        RECT 1903.090 1687.800 1903.410 1687.860 ;
        RECT 1465.630 15.880 1465.950 15.940 ;
        RECT 1469.310 15.880 1469.630 15.940 ;
        RECT 1465.630 15.740 1469.630 15.880 ;
        RECT 1465.630 15.680 1465.950 15.740 ;
        RECT 1469.310 15.680 1469.630 15.740 ;
      LAYER via ;
        RECT 1469.340 1687.800 1469.600 1688.060 ;
        RECT 1903.120 1687.800 1903.380 1688.060 ;
        RECT 1465.660 15.680 1465.920 15.940 ;
        RECT 1469.340 15.680 1469.600 15.940 ;
      LAYER met2 ;
        RECT 1903.040 1700.000 1903.320 1702.400 ;
        RECT 1903.180 1688.090 1903.320 1700.000 ;
        RECT 1469.340 1687.770 1469.600 1688.090 ;
        RECT 1903.120 1687.770 1903.380 1688.090 ;
        RECT 1469.400 15.970 1469.540 1687.770 ;
        RECT 1465.660 15.650 1465.920 15.970 ;
        RECT 1469.340 15.650 1469.600 15.970 ;
        RECT 1465.720 2.400 1465.860 15.650 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1907.690 1683.920 1908.010 1683.980 ;
        RECT 1912.290 1683.920 1912.610 1683.980 ;
        RECT 1907.690 1683.780 1912.610 1683.920 ;
        RECT 1907.690 1683.720 1908.010 1683.780 ;
        RECT 1912.290 1683.720 1912.610 1683.780 ;
        RECT 1483.570 17.920 1483.890 17.980 ;
        RECT 1907.690 17.920 1908.010 17.980 ;
        RECT 1483.570 17.780 1908.010 17.920 ;
        RECT 1483.570 17.720 1483.890 17.780 ;
        RECT 1907.690 17.720 1908.010 17.780 ;
      LAYER via ;
        RECT 1907.720 1683.720 1907.980 1683.980 ;
        RECT 1912.320 1683.720 1912.580 1683.980 ;
        RECT 1483.600 17.720 1483.860 17.980 ;
        RECT 1907.720 17.720 1907.980 17.980 ;
      LAYER met2 ;
        RECT 1912.240 1700.000 1912.520 1702.400 ;
        RECT 1912.380 1684.010 1912.520 1700.000 ;
        RECT 1907.720 1683.690 1907.980 1684.010 ;
        RECT 1912.320 1683.690 1912.580 1684.010 ;
        RECT 1907.780 18.010 1907.920 1683.690 ;
        RECT 1483.600 17.690 1483.860 18.010 ;
        RECT 1907.720 17.690 1907.980 18.010 ;
        RECT 1483.660 2.400 1483.800 17.690 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1872.805 1683.765 1872.975 1687.335 ;
      LAYER mcon ;
        RECT 1872.805 1687.165 1872.975 1687.335 ;
      LAYER met1 ;
        RECT 1920.110 1687.660 1920.430 1687.720 ;
        RECT 1885.240 1687.520 1920.430 1687.660 ;
        RECT 1872.745 1687.320 1873.035 1687.365 ;
        RECT 1885.240 1687.320 1885.380 1687.520 ;
        RECT 1920.110 1687.460 1920.430 1687.520 ;
        RECT 1872.745 1687.180 1885.380 1687.320 ;
        RECT 1872.745 1687.135 1873.035 1687.180 ;
        RECT 1817.990 1683.920 1818.310 1683.980 ;
        RECT 1872.745 1683.920 1873.035 1683.965 ;
        RECT 1817.990 1683.780 1873.035 1683.920 ;
        RECT 1817.990 1683.720 1818.310 1683.780 ;
        RECT 1872.745 1683.735 1873.035 1683.780 ;
        RECT 1501.510 19.960 1501.830 20.020 ;
        RECT 1817.990 19.960 1818.310 20.020 ;
        RECT 1501.510 19.820 1818.310 19.960 ;
        RECT 1501.510 19.760 1501.830 19.820 ;
        RECT 1817.990 19.760 1818.310 19.820 ;
      LAYER via ;
        RECT 1920.140 1687.460 1920.400 1687.720 ;
        RECT 1818.020 1683.720 1818.280 1683.980 ;
        RECT 1501.540 19.760 1501.800 20.020 ;
        RECT 1818.020 19.760 1818.280 20.020 ;
      LAYER met2 ;
        RECT 1921.440 1700.410 1921.720 1702.400 ;
        RECT 1920.200 1700.270 1921.720 1700.410 ;
        RECT 1920.200 1687.750 1920.340 1700.270 ;
        RECT 1921.440 1700.000 1921.720 1700.270 ;
        RECT 1920.140 1687.430 1920.400 1687.750 ;
        RECT 1818.020 1683.690 1818.280 1684.010 ;
        RECT 1818.080 20.050 1818.220 1683.690 ;
        RECT 1501.540 19.730 1501.800 20.050 ;
        RECT 1818.020 19.730 1818.280 20.050 ;
        RECT 1501.600 2.400 1501.740 19.730 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1914.590 1683.920 1914.910 1683.980 ;
        RECT 1930.690 1683.920 1931.010 1683.980 ;
        RECT 1914.590 1683.780 1931.010 1683.920 ;
        RECT 1914.590 1683.720 1914.910 1683.780 ;
        RECT 1930.690 1683.720 1931.010 1683.780 ;
        RECT 1518.990 18.260 1519.310 18.320 ;
        RECT 1914.590 18.260 1914.910 18.320 ;
        RECT 1518.990 18.120 1914.910 18.260 ;
        RECT 1518.990 18.060 1519.310 18.120 ;
        RECT 1914.590 18.060 1914.910 18.120 ;
      LAYER via ;
        RECT 1914.620 1683.720 1914.880 1683.980 ;
        RECT 1930.720 1683.720 1930.980 1683.980 ;
        RECT 1519.020 18.060 1519.280 18.320 ;
        RECT 1914.620 18.060 1914.880 18.320 ;
      LAYER met2 ;
        RECT 1930.640 1700.000 1930.920 1702.400 ;
        RECT 1930.780 1684.010 1930.920 1700.000 ;
        RECT 1914.620 1683.690 1914.880 1684.010 ;
        RECT 1930.720 1683.690 1930.980 1684.010 ;
        RECT 1914.680 18.350 1914.820 1683.690 ;
        RECT 1519.020 18.030 1519.280 18.350 ;
        RECT 1914.620 18.030 1914.880 18.350 ;
        RECT 1519.080 2.400 1519.220 18.030 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1511.630 1678.140 1511.950 1678.200 ;
        RECT 1515.310 1678.140 1515.630 1678.200 ;
        RECT 1511.630 1678.000 1515.630 1678.140 ;
        RECT 1511.630 1677.940 1511.950 1678.000 ;
        RECT 1515.310 1677.940 1515.630 1678.000 ;
        RECT 717.210 54.980 717.530 55.040 ;
        RECT 1511.630 54.980 1511.950 55.040 ;
        RECT 717.210 54.840 1511.950 54.980 ;
        RECT 717.210 54.780 717.530 54.840 ;
        RECT 1511.630 54.780 1511.950 54.840 ;
      LAYER via ;
        RECT 1511.660 1677.940 1511.920 1678.200 ;
        RECT 1515.340 1677.940 1515.600 1678.200 ;
        RECT 717.240 54.780 717.500 55.040 ;
        RECT 1511.660 54.780 1511.920 55.040 ;
      LAYER met2 ;
        RECT 1517.100 1700.410 1517.380 1702.400 ;
        RECT 1515.400 1700.270 1517.380 1700.410 ;
        RECT 1515.400 1678.230 1515.540 1700.270 ;
        RECT 1517.100 1700.000 1517.380 1700.270 ;
        RECT 1511.660 1677.910 1511.920 1678.230 ;
        RECT 1515.340 1677.910 1515.600 1678.230 ;
        RECT 1511.720 55.070 1511.860 1677.910 ;
        RECT 717.240 54.750 717.500 55.070 ;
        RECT 1511.660 54.750 1511.920 55.070 ;
        RECT 717.300 16.730 717.440 54.750 ;
        RECT 716.380 16.590 717.440 16.730 ;
        RECT 716.380 2.400 716.520 16.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1548.890 1689.700 1549.210 1689.760 ;
        RECT 1548.890 1689.560 1577.640 1689.700 ;
        RECT 1548.890 1689.500 1549.210 1689.560 ;
        RECT 1577.500 1689.360 1577.640 1689.560 ;
        RECT 1939.890 1689.360 1940.210 1689.420 ;
        RECT 1577.500 1689.220 1940.210 1689.360 ;
        RECT 1939.890 1689.160 1940.210 1689.220 ;
        RECT 1536.930 18.600 1537.250 18.660 ;
        RECT 1548.890 18.600 1549.210 18.660 ;
        RECT 1536.930 18.460 1549.210 18.600 ;
        RECT 1536.930 18.400 1537.250 18.460 ;
        RECT 1548.890 18.400 1549.210 18.460 ;
      LAYER via ;
        RECT 1548.920 1689.500 1549.180 1689.760 ;
        RECT 1939.920 1689.160 1940.180 1689.420 ;
        RECT 1536.960 18.400 1537.220 18.660 ;
        RECT 1548.920 18.400 1549.180 18.660 ;
      LAYER met2 ;
        RECT 1939.840 1700.000 1940.120 1702.400 ;
        RECT 1548.920 1689.470 1549.180 1689.790 ;
        RECT 1548.980 18.690 1549.120 1689.470 ;
        RECT 1939.980 1689.450 1940.120 1700.000 ;
        RECT 1939.920 1689.130 1940.180 1689.450 ;
        RECT 1536.960 18.370 1537.220 18.690 ;
        RECT 1548.920 18.370 1549.180 18.690 ;
        RECT 1537.020 2.400 1537.160 18.370 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1928.390 1689.700 1928.710 1689.760 ;
        RECT 1948.630 1689.700 1948.950 1689.760 ;
        RECT 1928.390 1689.560 1948.950 1689.700 ;
        RECT 1928.390 1689.500 1928.710 1689.560 ;
        RECT 1948.630 1689.500 1948.950 1689.560 ;
        RECT 1554.870 14.180 1555.190 14.240 ;
        RECT 1928.390 14.180 1928.710 14.240 ;
        RECT 1554.870 14.040 1928.710 14.180 ;
        RECT 1554.870 13.980 1555.190 14.040 ;
        RECT 1928.390 13.980 1928.710 14.040 ;
      LAYER via ;
        RECT 1928.420 1689.500 1928.680 1689.760 ;
        RECT 1948.660 1689.500 1948.920 1689.760 ;
        RECT 1554.900 13.980 1555.160 14.240 ;
        RECT 1928.420 13.980 1928.680 14.240 ;
      LAYER met2 ;
        RECT 1948.580 1700.000 1948.860 1702.400 ;
        RECT 1948.720 1689.790 1948.860 1700.000 ;
        RECT 1928.420 1689.470 1928.680 1689.790 ;
        RECT 1948.660 1689.470 1948.920 1689.790 ;
        RECT 1928.480 14.270 1928.620 1689.470 ;
        RECT 1554.900 13.950 1555.160 14.270 ;
        RECT 1928.420 13.950 1928.680 14.270 ;
        RECT 1554.960 2.400 1555.100 13.950 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1631.765 1685.805 1631.935 1689.715 ;
        RECT 1921.565 1687.845 1921.735 1689.715 ;
      LAYER mcon ;
        RECT 1631.765 1689.545 1631.935 1689.715 ;
        RECT 1921.565 1689.545 1921.735 1689.715 ;
      LAYER met1 ;
        RECT 1631.705 1689.700 1631.995 1689.745 ;
        RECT 1921.505 1689.700 1921.795 1689.745 ;
        RECT 1631.705 1689.560 1921.795 1689.700 ;
        RECT 1631.705 1689.515 1631.995 1689.560 ;
        RECT 1921.505 1689.515 1921.795 1689.560 ;
        RECT 1921.505 1688.000 1921.795 1688.045 ;
        RECT 1957.830 1688.000 1958.150 1688.060 ;
        RECT 1921.505 1687.860 1958.150 1688.000 ;
        RECT 1921.505 1687.815 1921.795 1687.860 ;
        RECT 1957.830 1687.800 1958.150 1687.860 ;
        RECT 1583.390 1685.960 1583.710 1686.020 ;
        RECT 1631.705 1685.960 1631.995 1686.005 ;
        RECT 1583.390 1685.820 1631.995 1685.960 ;
        RECT 1583.390 1685.760 1583.710 1685.820 ;
        RECT 1631.705 1685.775 1631.995 1685.820 ;
        RECT 1572.810 20.640 1573.130 20.700 ;
        RECT 1583.390 20.640 1583.710 20.700 ;
        RECT 1572.810 20.500 1583.710 20.640 ;
        RECT 1572.810 20.440 1573.130 20.500 ;
        RECT 1583.390 20.440 1583.710 20.500 ;
      LAYER via ;
        RECT 1957.860 1687.800 1958.120 1688.060 ;
        RECT 1583.420 1685.760 1583.680 1686.020 ;
        RECT 1572.840 20.440 1573.100 20.700 ;
        RECT 1583.420 20.440 1583.680 20.700 ;
      LAYER met2 ;
        RECT 1957.780 1700.000 1958.060 1702.400 ;
        RECT 1957.920 1688.090 1958.060 1700.000 ;
        RECT 1957.860 1687.770 1958.120 1688.090 ;
        RECT 1583.420 1685.730 1583.680 1686.050 ;
        RECT 1583.480 20.730 1583.620 1685.730 ;
        RECT 1572.840 20.410 1573.100 20.730 ;
        RECT 1583.420 20.410 1583.680 20.730 ;
        RECT 1572.900 2.400 1573.040 20.410 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1949.550 1683.920 1949.870 1683.980 ;
        RECT 1967.030 1683.920 1967.350 1683.980 ;
        RECT 1949.550 1683.780 1967.350 1683.920 ;
        RECT 1949.550 1683.720 1949.870 1683.780 ;
        RECT 1967.030 1683.720 1967.350 1683.780 ;
        RECT 1590.290 18.940 1590.610 19.000 ;
        RECT 1949.090 18.940 1949.410 19.000 ;
        RECT 1590.290 18.800 1949.410 18.940 ;
        RECT 1590.290 18.740 1590.610 18.800 ;
        RECT 1949.090 18.740 1949.410 18.800 ;
      LAYER via ;
        RECT 1949.580 1683.720 1949.840 1683.980 ;
        RECT 1967.060 1683.720 1967.320 1683.980 ;
        RECT 1590.320 18.740 1590.580 19.000 ;
        RECT 1949.120 18.740 1949.380 19.000 ;
      LAYER met2 ;
        RECT 1966.980 1700.000 1967.260 1702.400 ;
        RECT 1967.120 1684.010 1967.260 1700.000 ;
        RECT 1949.580 1683.690 1949.840 1684.010 ;
        RECT 1967.060 1683.690 1967.320 1684.010 ;
        RECT 1949.640 1677.970 1949.780 1683.690 ;
        RECT 1949.180 1677.830 1949.780 1677.970 ;
        RECT 1949.180 19.030 1949.320 1677.830 ;
        RECT 1590.320 18.710 1590.580 19.030 ;
        RECT 1949.120 18.710 1949.380 19.030 ;
        RECT 1590.380 2.400 1590.520 18.710 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1613.750 1690.040 1614.070 1690.100 ;
        RECT 1976.230 1690.040 1976.550 1690.100 ;
        RECT 1613.750 1689.900 1976.550 1690.040 ;
        RECT 1613.750 1689.840 1614.070 1689.900 ;
        RECT 1976.230 1689.840 1976.550 1689.900 ;
        RECT 1608.230 20.640 1608.550 20.700 ;
        RECT 1613.750 20.640 1614.070 20.700 ;
        RECT 1608.230 20.500 1614.070 20.640 ;
        RECT 1608.230 20.440 1608.550 20.500 ;
        RECT 1613.750 20.440 1614.070 20.500 ;
      LAYER via ;
        RECT 1613.780 1689.840 1614.040 1690.100 ;
        RECT 1976.260 1689.840 1976.520 1690.100 ;
        RECT 1608.260 20.440 1608.520 20.700 ;
        RECT 1613.780 20.440 1614.040 20.700 ;
      LAYER met2 ;
        RECT 1976.180 1700.000 1976.460 1702.400 ;
        RECT 1976.320 1690.130 1976.460 1700.000 ;
        RECT 1613.780 1689.810 1614.040 1690.130 ;
        RECT 1976.260 1689.810 1976.520 1690.130 ;
        RECT 1613.840 20.730 1613.980 1689.810 ;
        RECT 1608.260 20.410 1608.520 20.730 ;
        RECT 1613.780 20.410 1614.040 20.730 ;
        RECT 1608.320 2.400 1608.460 20.410 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1955.990 1689.360 1956.310 1689.420 ;
        RECT 1985.430 1689.360 1985.750 1689.420 ;
        RECT 1955.990 1689.220 1985.750 1689.360 ;
        RECT 1955.990 1689.160 1956.310 1689.220 ;
        RECT 1985.430 1689.160 1985.750 1689.220 ;
        RECT 1626.170 19.620 1626.490 19.680 ;
        RECT 1955.530 19.620 1955.850 19.680 ;
        RECT 1626.170 19.480 1955.850 19.620 ;
        RECT 1626.170 19.420 1626.490 19.480 ;
        RECT 1955.530 19.420 1955.850 19.480 ;
      LAYER via ;
        RECT 1956.020 1689.160 1956.280 1689.420 ;
        RECT 1985.460 1689.160 1985.720 1689.420 ;
        RECT 1626.200 19.420 1626.460 19.680 ;
        RECT 1955.560 19.420 1955.820 19.680 ;
      LAYER met2 ;
        RECT 1985.380 1700.000 1985.660 1702.400 ;
        RECT 1985.520 1689.450 1985.660 1700.000 ;
        RECT 1956.020 1689.130 1956.280 1689.450 ;
        RECT 1985.460 1689.130 1985.720 1689.450 ;
        RECT 1956.080 20.130 1956.220 1689.130 ;
        RECT 1955.620 19.990 1956.220 20.130 ;
        RECT 1955.620 19.710 1955.760 19.990 ;
        RECT 1626.200 19.390 1626.460 19.710 ;
        RECT 1955.560 19.390 1955.820 19.710 ;
        RECT 1626.260 2.400 1626.400 19.390 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1818.450 1684.600 1818.770 1684.660 ;
        RECT 1818.450 1684.460 1970.020 1684.600 ;
        RECT 1818.450 1684.400 1818.770 1684.460 ;
        RECT 1969.880 1684.260 1970.020 1684.460 ;
        RECT 1994.630 1684.260 1994.950 1684.320 ;
        RECT 1969.880 1684.120 1994.950 1684.260 ;
        RECT 1994.630 1684.060 1994.950 1684.120 ;
        RECT 1644.110 16.220 1644.430 16.280 ;
        RECT 1818.450 16.220 1818.770 16.280 ;
        RECT 1644.110 16.080 1818.770 16.220 ;
        RECT 1644.110 16.020 1644.430 16.080 ;
        RECT 1818.450 16.020 1818.770 16.080 ;
      LAYER via ;
        RECT 1818.480 1684.400 1818.740 1684.660 ;
        RECT 1994.660 1684.060 1994.920 1684.320 ;
        RECT 1644.140 16.020 1644.400 16.280 ;
        RECT 1818.480 16.020 1818.740 16.280 ;
      LAYER met2 ;
        RECT 1994.580 1700.000 1994.860 1702.400 ;
        RECT 1818.480 1684.370 1818.740 1684.690 ;
        RECT 1818.540 16.310 1818.680 1684.370 ;
        RECT 1994.720 1684.350 1994.860 1700.000 ;
        RECT 1994.660 1684.030 1994.920 1684.350 ;
        RECT 1644.140 15.990 1644.400 16.310 ;
        RECT 1818.480 15.990 1818.740 16.310 ;
        RECT 1644.200 2.400 1644.340 15.990 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1977.150 1684.600 1977.470 1684.660 ;
        RECT 2003.830 1684.600 2004.150 1684.660 ;
        RECT 1977.150 1684.460 2004.150 1684.600 ;
        RECT 1977.150 1684.400 1977.470 1684.460 ;
        RECT 2003.830 1684.400 2004.150 1684.460 ;
        RECT 1662.050 19.280 1662.370 19.340 ;
        RECT 1662.050 19.140 1961.280 19.280 ;
        RECT 1662.050 19.080 1662.370 19.140 ;
        RECT 1961.140 18.940 1961.280 19.140 ;
        RECT 1976.690 18.940 1977.010 19.000 ;
        RECT 1961.140 18.800 1977.010 18.940 ;
        RECT 1976.690 18.740 1977.010 18.800 ;
      LAYER via ;
        RECT 1977.180 1684.400 1977.440 1684.660 ;
        RECT 2003.860 1684.400 2004.120 1684.660 ;
        RECT 1662.080 19.080 1662.340 19.340 ;
        RECT 1976.720 18.740 1976.980 19.000 ;
      LAYER met2 ;
        RECT 2003.780 1700.000 2004.060 1702.400 ;
        RECT 2003.920 1684.690 2004.060 1700.000 ;
        RECT 1977.180 1684.370 1977.440 1684.690 ;
        RECT 2003.860 1684.370 2004.120 1684.690 ;
        RECT 1977.240 1670.490 1977.380 1684.370 ;
        RECT 1976.780 1670.350 1977.380 1670.490 ;
        RECT 1662.080 19.050 1662.340 19.370 ;
        RECT 1662.140 2.400 1662.280 19.050 ;
        RECT 1976.780 19.030 1976.920 1670.350 ;
        RECT 1976.720 18.710 1976.980 19.030 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1969.405 1684.105 1969.575 1689.715 ;
        RECT 1816.225 15.385 1816.395 16.575 ;
      LAYER mcon ;
        RECT 1969.405 1689.545 1969.575 1689.715 ;
        RECT 1816.225 16.405 1816.395 16.575 ;
      LAYER met1 ;
        RECT 2013.030 1690.040 2013.350 1690.100 ;
        RECT 1976.780 1689.900 2013.350 1690.040 ;
        RECT 1969.345 1689.700 1969.635 1689.745 ;
        RECT 1976.780 1689.700 1976.920 1689.900 ;
        RECT 2013.030 1689.840 2013.350 1689.900 ;
        RECT 1969.345 1689.560 1976.920 1689.700 ;
        RECT 1969.345 1689.515 1969.635 1689.560 ;
        RECT 1832.250 1684.260 1832.570 1684.320 ;
        RECT 1969.345 1684.260 1969.635 1684.305 ;
        RECT 1832.250 1684.120 1969.635 1684.260 ;
        RECT 1832.250 1684.060 1832.570 1684.120 ;
        RECT 1969.345 1684.075 1969.635 1684.120 ;
        RECT 1816.165 16.560 1816.455 16.605 ;
        RECT 1832.250 16.560 1832.570 16.620 ;
        RECT 1816.165 16.420 1832.570 16.560 ;
        RECT 1816.165 16.375 1816.455 16.420 ;
        RECT 1832.250 16.360 1832.570 16.420 ;
        RECT 1679.530 15.540 1679.850 15.600 ;
        RECT 1816.165 15.540 1816.455 15.585 ;
        RECT 1679.530 15.400 1816.455 15.540 ;
        RECT 1679.530 15.340 1679.850 15.400 ;
        RECT 1816.165 15.355 1816.455 15.400 ;
      LAYER via ;
        RECT 2013.060 1689.840 2013.320 1690.100 ;
        RECT 1832.280 1684.060 1832.540 1684.320 ;
        RECT 1832.280 16.360 1832.540 16.620 ;
        RECT 1679.560 15.340 1679.820 15.600 ;
      LAYER met2 ;
        RECT 2012.980 1700.000 2013.260 1702.400 ;
        RECT 2013.120 1690.130 2013.260 1700.000 ;
        RECT 2013.060 1689.810 2013.320 1690.130 ;
        RECT 1832.280 1684.030 1832.540 1684.350 ;
        RECT 1832.340 16.650 1832.480 1684.030 ;
        RECT 1832.280 16.330 1832.540 16.650 ;
        RECT 1679.560 15.310 1679.820 15.630 ;
        RECT 1679.620 2.400 1679.760 15.310 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1964.805 19.125 1964.975 20.315 ;
      LAYER mcon ;
        RECT 1964.805 20.145 1964.975 20.315 ;
      LAYER met1 ;
        RECT 2022.230 1684.260 2022.550 1684.320 ;
        RECT 2004.380 1684.120 2022.550 1684.260 ;
        RECT 1983.590 1683.920 1983.910 1683.980 ;
        RECT 2004.380 1683.920 2004.520 1684.120 ;
        RECT 2022.230 1684.060 2022.550 1684.120 ;
        RECT 1983.590 1683.780 2004.520 1683.920 ;
        RECT 1983.590 1683.720 1983.910 1683.780 ;
        RECT 1697.470 20.300 1697.790 20.360 ;
        RECT 1964.745 20.300 1965.035 20.345 ;
        RECT 1697.470 20.160 1965.035 20.300 ;
        RECT 1697.470 20.100 1697.790 20.160 ;
        RECT 1964.745 20.115 1965.035 20.160 ;
        RECT 1964.745 19.280 1965.035 19.325 ;
        RECT 1983.590 19.280 1983.910 19.340 ;
        RECT 1964.745 19.140 1983.910 19.280 ;
        RECT 1964.745 19.095 1965.035 19.140 ;
        RECT 1983.590 19.080 1983.910 19.140 ;
      LAYER via ;
        RECT 1983.620 1683.720 1983.880 1683.980 ;
        RECT 2022.260 1684.060 2022.520 1684.320 ;
        RECT 1697.500 20.100 1697.760 20.360 ;
        RECT 1983.620 19.080 1983.880 19.340 ;
      LAYER met2 ;
        RECT 2022.180 1700.000 2022.460 1702.400 ;
        RECT 2022.320 1684.350 2022.460 1700.000 ;
        RECT 2022.260 1684.030 2022.520 1684.350 ;
        RECT 1983.620 1683.690 1983.880 1684.010 ;
        RECT 1697.500 20.070 1697.760 20.390 ;
        RECT 1697.560 2.400 1697.700 20.070 ;
        RECT 1983.680 19.370 1983.820 1683.690 ;
        RECT 1983.620 19.050 1983.880 19.370 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 51.240 738.230 51.300 ;
        RECT 1524.970 51.240 1525.290 51.300 ;
        RECT 737.910 51.100 1525.290 51.240 ;
        RECT 737.910 51.040 738.230 51.100 ;
        RECT 1524.970 51.040 1525.290 51.100 ;
      LAYER via ;
        RECT 737.940 51.040 738.200 51.300 ;
        RECT 1525.000 51.040 1525.260 51.300 ;
      LAYER met2 ;
        RECT 1526.300 1700.410 1526.580 1702.400 ;
        RECT 1525.060 1700.270 1526.580 1700.410 ;
        RECT 1525.060 51.330 1525.200 1700.270 ;
        RECT 1526.300 1700.000 1526.580 1700.270 ;
        RECT 737.940 51.010 738.200 51.330 ;
        RECT 1525.000 51.010 1525.260 51.330 ;
        RECT 738.000 16.730 738.140 51.010 ;
        RECT 734.320 16.590 738.140 16.730 ;
        RECT 734.320 2.400 734.460 16.590 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1849.345 14.365 1849.515 15.895 ;
      LAYER mcon ;
        RECT 1849.345 15.725 1849.515 15.895 ;
      LAYER met1 ;
        RECT 2031.430 1689.020 2031.750 1689.080 ;
        RECT 1921.580 1688.880 2031.750 1689.020 ;
        RECT 1880.090 1688.680 1880.410 1688.740 ;
        RECT 1921.580 1688.680 1921.720 1688.880 ;
        RECT 2031.430 1688.820 2031.750 1688.880 ;
        RECT 1880.090 1688.540 1921.720 1688.680 ;
        RECT 1880.090 1688.480 1880.410 1688.540 ;
        RECT 1715.410 15.880 1715.730 15.940 ;
        RECT 1849.285 15.880 1849.575 15.925 ;
        RECT 1715.410 15.740 1849.575 15.880 ;
        RECT 1715.410 15.680 1715.730 15.740 ;
        RECT 1849.285 15.695 1849.575 15.740 ;
        RECT 1849.285 14.520 1849.575 14.565 ;
        RECT 1880.090 14.520 1880.410 14.580 ;
        RECT 1849.285 14.380 1880.410 14.520 ;
        RECT 1849.285 14.335 1849.575 14.380 ;
        RECT 1880.090 14.320 1880.410 14.380 ;
      LAYER via ;
        RECT 1880.120 1688.480 1880.380 1688.740 ;
        RECT 2031.460 1688.820 2031.720 1689.080 ;
        RECT 1715.440 15.680 1715.700 15.940 ;
        RECT 1880.120 14.320 1880.380 14.580 ;
      LAYER met2 ;
        RECT 2031.380 1700.000 2031.660 1702.400 ;
        RECT 2031.520 1689.110 2031.660 1700.000 ;
        RECT 2031.460 1688.790 2031.720 1689.110 ;
        RECT 1880.120 1688.450 1880.380 1688.770 ;
        RECT 1715.440 15.650 1715.700 15.970 ;
        RECT 1715.500 2.400 1715.640 15.650 ;
        RECT 1880.180 14.610 1880.320 1688.450 ;
        RECT 1880.120 14.290 1880.380 14.610 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1956.065 19.465 1956.235 20.655 ;
      LAYER mcon ;
        RECT 1956.065 20.485 1956.235 20.655 ;
      LAYER met1 ;
        RECT 2005.210 1683.920 2005.530 1683.980 ;
        RECT 2040.630 1683.920 2040.950 1683.980 ;
        RECT 2005.210 1683.780 2040.950 1683.920 ;
        RECT 2005.210 1683.720 2005.530 1683.780 ;
        RECT 2040.630 1683.720 2040.950 1683.780 ;
        RECT 1733.350 20.640 1733.670 20.700 ;
        RECT 1956.005 20.640 1956.295 20.685 ;
        RECT 1733.350 20.500 1956.295 20.640 ;
        RECT 1733.350 20.440 1733.670 20.500 ;
        RECT 1956.005 20.455 1956.295 20.500 ;
        RECT 1956.005 19.620 1956.295 19.665 ;
        RECT 2004.290 19.620 2004.610 19.680 ;
        RECT 1956.005 19.480 2004.610 19.620 ;
        RECT 1956.005 19.435 1956.295 19.480 ;
        RECT 2004.290 19.420 2004.610 19.480 ;
      LAYER via ;
        RECT 2005.240 1683.720 2005.500 1683.980 ;
        RECT 2040.660 1683.720 2040.920 1683.980 ;
        RECT 1733.380 20.440 1733.640 20.700 ;
        RECT 2004.320 19.420 2004.580 19.680 ;
      LAYER met2 ;
        RECT 2040.580 1700.000 2040.860 1702.400 ;
        RECT 2040.720 1684.010 2040.860 1700.000 ;
        RECT 2005.240 1683.690 2005.500 1684.010 ;
        RECT 2040.660 1683.690 2040.920 1684.010 ;
        RECT 2005.300 1677.290 2005.440 1683.690 ;
        RECT 2004.380 1677.150 2005.440 1677.290 ;
        RECT 1733.380 20.410 1733.640 20.730 ;
        RECT 1733.440 2.400 1733.580 20.410 ;
        RECT 2004.380 19.710 2004.520 1677.150 ;
        RECT 2004.320 19.390 2004.580 19.710 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1922.025 1687.505 1922.195 1688.695 ;
        RECT 1907.305 1683.765 1907.475 1687.335 ;
      LAYER mcon ;
        RECT 1922.025 1688.525 1922.195 1688.695 ;
        RECT 1907.305 1687.165 1907.475 1687.335 ;
      LAYER met1 ;
        RECT 1921.965 1688.680 1922.255 1688.725 ;
        RECT 2049.830 1688.680 2050.150 1688.740 ;
        RECT 1921.965 1688.540 2050.150 1688.680 ;
        RECT 1921.965 1688.495 1922.255 1688.540 ;
        RECT 2049.830 1688.480 2050.150 1688.540 ;
        RECT 1921.965 1687.660 1922.255 1687.705 ;
        RECT 1920.660 1687.520 1922.255 1687.660 ;
        RECT 1907.245 1687.320 1907.535 1687.365 ;
        RECT 1920.660 1687.320 1920.800 1687.520 ;
        RECT 1921.965 1687.475 1922.255 1687.520 ;
        RECT 1907.245 1687.180 1920.800 1687.320 ;
        RECT 1907.245 1687.135 1907.535 1687.180 ;
        RECT 1873.190 1683.920 1873.510 1683.980 ;
        RECT 1907.245 1683.920 1907.535 1683.965 ;
        RECT 1873.190 1683.780 1907.535 1683.920 ;
        RECT 1873.190 1683.720 1873.510 1683.780 ;
        RECT 1907.245 1683.735 1907.535 1683.780 ;
        RECT 1873.190 15.540 1873.510 15.600 ;
        RECT 1861.320 15.400 1873.510 15.540 ;
        RECT 1751.290 15.200 1751.610 15.260 ;
        RECT 1861.320 15.200 1861.460 15.400 ;
        RECT 1873.190 15.340 1873.510 15.400 ;
        RECT 1751.290 15.060 1861.460 15.200 ;
        RECT 1751.290 15.000 1751.610 15.060 ;
      LAYER via ;
        RECT 2049.860 1688.480 2050.120 1688.740 ;
        RECT 1873.220 1683.720 1873.480 1683.980 ;
        RECT 1751.320 15.000 1751.580 15.260 ;
        RECT 1873.220 15.340 1873.480 15.600 ;
      LAYER met2 ;
        RECT 2049.780 1700.000 2050.060 1702.400 ;
        RECT 2049.920 1688.770 2050.060 1700.000 ;
        RECT 2049.860 1688.450 2050.120 1688.770 ;
        RECT 1873.220 1683.690 1873.480 1684.010 ;
        RECT 1873.280 15.630 1873.420 1683.690 ;
        RECT 1873.220 15.310 1873.480 15.630 ;
        RECT 1751.320 14.970 1751.580 15.290 ;
        RECT 1751.380 2.400 1751.520 14.970 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1969.865 16.745 1970.035 20.315 ;
        RECT 2000.225 19.125 2000.395 20.315 ;
        RECT 2016.785 19.125 2016.955 20.995 ;
      LAYER mcon ;
        RECT 2016.785 20.825 2016.955 20.995 ;
        RECT 1969.865 20.145 1970.035 20.315 ;
        RECT 2000.225 20.145 2000.395 20.315 ;
      LAYER met1 ;
        RECT 2024.990 1690.380 2025.310 1690.440 ;
        RECT 2059.030 1690.380 2059.350 1690.440 ;
        RECT 2024.990 1690.240 2059.350 1690.380 ;
        RECT 2024.990 1690.180 2025.310 1690.240 ;
        RECT 2059.030 1690.180 2059.350 1690.240 ;
        RECT 2016.725 20.980 2017.015 21.025 ;
        RECT 2024.990 20.980 2025.310 21.040 ;
        RECT 2016.725 20.840 2025.310 20.980 ;
        RECT 2016.725 20.795 2017.015 20.840 ;
        RECT 2024.990 20.780 2025.310 20.840 ;
        RECT 1969.805 20.300 1970.095 20.345 ;
        RECT 2000.165 20.300 2000.455 20.345 ;
        RECT 1969.805 20.160 2000.455 20.300 ;
        RECT 1969.805 20.115 1970.095 20.160 ;
        RECT 2000.165 20.115 2000.455 20.160 ;
        RECT 2000.165 19.280 2000.455 19.325 ;
        RECT 2016.725 19.280 2017.015 19.325 ;
        RECT 2000.165 19.140 2017.015 19.280 ;
        RECT 2000.165 19.095 2000.455 19.140 ;
        RECT 2016.725 19.095 2017.015 19.140 ;
        RECT 1768.770 16.900 1769.090 16.960 ;
        RECT 1969.805 16.900 1970.095 16.945 ;
        RECT 1768.770 16.760 1970.095 16.900 ;
        RECT 1768.770 16.700 1769.090 16.760 ;
        RECT 1969.805 16.715 1970.095 16.760 ;
      LAYER via ;
        RECT 2025.020 1690.180 2025.280 1690.440 ;
        RECT 2059.060 1690.180 2059.320 1690.440 ;
        RECT 2025.020 20.780 2025.280 21.040 ;
        RECT 1768.800 16.700 1769.060 16.960 ;
      LAYER met2 ;
        RECT 2058.980 1700.000 2059.260 1702.400 ;
        RECT 2059.120 1690.470 2059.260 1700.000 ;
        RECT 2025.020 1690.150 2025.280 1690.470 ;
        RECT 2059.060 1690.150 2059.320 1690.470 ;
        RECT 2025.080 21.070 2025.220 1690.150 ;
        RECT 2025.020 20.750 2025.280 21.070 ;
        RECT 1768.800 16.670 1769.060 16.990 ;
        RECT 1768.860 2.400 1769.000 16.670 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1786.710 1685.620 1787.030 1685.680 ;
        RECT 2068.230 1685.620 2068.550 1685.680 ;
        RECT 1786.710 1685.480 2068.550 1685.620 ;
        RECT 1786.710 1685.420 1787.030 1685.480 ;
        RECT 2068.230 1685.420 2068.550 1685.480 ;
      LAYER via ;
        RECT 1786.740 1685.420 1787.000 1685.680 ;
        RECT 2068.260 1685.420 2068.520 1685.680 ;
      LAYER met2 ;
        RECT 2068.180 1700.000 2068.460 1702.400 ;
        RECT 2068.320 1685.710 2068.460 1700.000 ;
        RECT 1786.740 1685.390 1787.000 1685.710 ;
        RECT 2068.260 1685.390 2068.520 1685.710 ;
        RECT 1786.800 2.400 1786.940 1685.390 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1873.725 14.705 1873.895 17.255 ;
        RECT 2012.185 16.065 2012.355 17.255 ;
        RECT 2017.705 16.405 2019.255 16.575 ;
        RECT 2017.705 16.235 2017.875 16.405 ;
        RECT 2016.785 16.065 2017.875 16.235 ;
      LAYER mcon ;
        RECT 1873.725 17.085 1873.895 17.255 ;
        RECT 2012.185 17.085 2012.355 17.255 ;
        RECT 2019.085 16.405 2019.255 16.575 ;
      LAYER met1 ;
        RECT 2038.790 1689.700 2039.110 1689.760 ;
        RECT 2077.430 1689.700 2077.750 1689.760 ;
        RECT 2038.790 1689.560 2077.750 1689.700 ;
        RECT 2038.790 1689.500 2039.110 1689.560 ;
        RECT 2077.430 1689.500 2077.750 1689.560 ;
        RECT 1873.665 17.240 1873.955 17.285 ;
        RECT 2012.125 17.240 2012.415 17.285 ;
        RECT 1873.665 17.100 2012.415 17.240 ;
        RECT 1873.665 17.055 1873.955 17.100 ;
        RECT 2012.125 17.055 2012.415 17.100 ;
        RECT 2019.025 16.560 2019.315 16.605 ;
        RECT 2035.570 16.560 2035.890 16.620 ;
        RECT 2019.025 16.420 2035.890 16.560 ;
        RECT 2019.025 16.375 2019.315 16.420 ;
        RECT 2035.570 16.360 2035.890 16.420 ;
        RECT 2012.125 16.220 2012.415 16.265 ;
        RECT 2016.725 16.220 2017.015 16.265 ;
        RECT 2012.125 16.080 2017.015 16.220 ;
        RECT 2012.125 16.035 2012.415 16.080 ;
        RECT 2016.725 16.035 2017.015 16.080 ;
        RECT 1804.650 14.860 1804.970 14.920 ;
        RECT 1873.665 14.860 1873.955 14.905 ;
        RECT 1804.650 14.720 1873.955 14.860 ;
        RECT 1804.650 14.660 1804.970 14.720 ;
        RECT 1873.665 14.675 1873.955 14.720 ;
      LAYER via ;
        RECT 2038.820 1689.500 2039.080 1689.760 ;
        RECT 2077.460 1689.500 2077.720 1689.760 ;
        RECT 2035.600 16.360 2035.860 16.620 ;
        RECT 1804.680 14.660 1804.940 14.920 ;
      LAYER met2 ;
        RECT 2077.380 1700.000 2077.660 1702.400 ;
        RECT 2077.520 1689.790 2077.660 1700.000 ;
        RECT 2038.820 1689.470 2039.080 1689.790 ;
        RECT 2077.460 1689.470 2077.720 1689.790 ;
        RECT 2038.880 24.380 2039.020 1689.470 ;
        RECT 2037.040 24.240 2039.020 24.380 ;
        RECT 2037.040 17.240 2037.180 24.240 ;
        RECT 2035.660 17.100 2037.180 17.240 ;
        RECT 2035.660 16.650 2035.800 17.100 ;
        RECT 2035.600 16.330 2035.860 16.650 ;
        RECT 1804.680 14.630 1804.940 14.950 ;
        RECT 1804.740 2.400 1804.880 14.630 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2042.545 1684.785 2042.715 1686.315 ;
      LAYER mcon ;
        RECT 2042.545 1686.145 2042.715 1686.315 ;
      LAYER met1 ;
        RECT 2042.485 1686.300 2042.775 1686.345 ;
        RECT 2042.485 1686.160 2056.500 1686.300 ;
        RECT 2042.485 1686.115 2042.775 1686.160 ;
        RECT 2056.360 1685.960 2056.500 1686.160 ;
        RECT 2086.630 1685.960 2086.950 1686.020 ;
        RECT 2056.360 1685.820 2086.950 1685.960 ;
        RECT 2086.630 1685.760 2086.950 1685.820 ;
        RECT 1831.790 1684.940 1832.110 1685.000 ;
        RECT 2042.485 1684.940 2042.775 1684.985 ;
        RECT 1831.790 1684.800 2042.775 1684.940 ;
        RECT 1831.790 1684.740 1832.110 1684.800 ;
        RECT 2042.485 1684.755 2042.775 1684.800 ;
        RECT 1822.590 19.960 1822.910 20.020 ;
        RECT 1831.790 19.960 1832.110 20.020 ;
        RECT 1822.590 19.820 1832.110 19.960 ;
        RECT 1822.590 19.760 1822.910 19.820 ;
        RECT 1831.790 19.760 1832.110 19.820 ;
      LAYER via ;
        RECT 2086.660 1685.760 2086.920 1686.020 ;
        RECT 1831.820 1684.740 1832.080 1685.000 ;
        RECT 1822.620 19.760 1822.880 20.020 ;
        RECT 1831.820 19.760 1832.080 20.020 ;
      LAYER met2 ;
        RECT 2086.580 1700.000 2086.860 1702.400 ;
        RECT 2086.720 1686.050 2086.860 1700.000 ;
        RECT 2086.660 1685.730 2086.920 1686.050 ;
        RECT 1831.820 1684.710 1832.080 1685.030 ;
        RECT 1831.880 20.050 1832.020 1684.710 ;
        RECT 1822.620 19.730 1822.880 20.050 ;
        RECT 1831.820 19.730 1832.080 20.050 ;
        RECT 1822.680 2.400 1822.820 19.730 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2042.545 20.145 2046.395 20.315 ;
        RECT 1873.265 17.085 1873.435 18.615 ;
        RECT 1921.565 18.445 1921.735 19.975 ;
      LAYER mcon ;
        RECT 2046.225 20.145 2046.395 20.315 ;
        RECT 1921.565 19.805 1921.735 19.975 ;
        RECT 1873.265 18.445 1873.435 18.615 ;
      LAYER met1 ;
        RECT 2060.410 1690.380 2060.730 1690.440 ;
        RECT 2095.830 1690.380 2096.150 1690.440 ;
        RECT 2060.410 1690.240 2096.150 1690.380 ;
        RECT 2060.410 1690.180 2060.730 1690.240 ;
        RECT 2095.830 1690.180 2096.150 1690.240 ;
        RECT 2059.490 20.640 2059.810 20.700 ;
        RECT 2053.140 20.500 2059.810 20.640 ;
        RECT 2042.485 20.300 2042.775 20.345 ;
        RECT 2018.180 20.160 2042.775 20.300 ;
        RECT 1921.505 19.960 1921.795 20.005 ;
        RECT 2018.180 19.960 2018.320 20.160 ;
        RECT 2042.485 20.115 2042.775 20.160 ;
        RECT 2046.165 20.300 2046.455 20.345 ;
        RECT 2053.140 20.300 2053.280 20.500 ;
        RECT 2059.490 20.440 2059.810 20.500 ;
        RECT 2046.165 20.160 2053.280 20.300 ;
        RECT 2046.165 20.115 2046.455 20.160 ;
        RECT 1921.505 19.820 2018.320 19.960 ;
        RECT 1921.505 19.775 1921.795 19.820 ;
        RECT 1873.205 18.600 1873.495 18.645 ;
        RECT 1921.505 18.600 1921.795 18.645 ;
        RECT 1873.205 18.460 1921.795 18.600 ;
        RECT 1873.205 18.415 1873.495 18.460 ;
        RECT 1921.505 18.415 1921.795 18.460 ;
        RECT 1840.070 17.240 1840.390 17.300 ;
        RECT 1873.205 17.240 1873.495 17.285 ;
        RECT 1840.070 17.100 1873.495 17.240 ;
        RECT 1840.070 17.040 1840.390 17.100 ;
        RECT 1873.205 17.055 1873.495 17.100 ;
      LAYER via ;
        RECT 2060.440 1690.180 2060.700 1690.440 ;
        RECT 2095.860 1690.180 2096.120 1690.440 ;
        RECT 2059.520 20.440 2059.780 20.700 ;
        RECT 1840.100 17.040 1840.360 17.300 ;
      LAYER met2 ;
        RECT 2095.780 1700.000 2096.060 1702.400 ;
        RECT 2095.920 1690.470 2096.060 1700.000 ;
        RECT 2060.440 1690.150 2060.700 1690.470 ;
        RECT 2095.860 1690.150 2096.120 1690.470 ;
        RECT 2060.500 1656.210 2060.640 1690.150 ;
        RECT 2059.580 1656.070 2060.640 1656.210 ;
        RECT 2059.580 20.730 2059.720 1656.070 ;
        RECT 2059.520 20.410 2059.780 20.730 ;
        RECT 1840.100 17.010 1840.360 17.330 ;
        RECT 1840.160 2.400 1840.300 17.010 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1896.740 1687.180 1898.260 1687.320 ;
        RECT 1862.610 1686.980 1862.930 1687.040 ;
        RECT 1896.740 1686.980 1896.880 1687.180 ;
        RECT 1862.610 1686.840 1896.880 1686.980 ;
        RECT 1898.120 1686.980 1898.260 1687.180 ;
        RECT 2105.030 1686.980 2105.350 1687.040 ;
        RECT 1898.120 1686.840 2105.350 1686.980 ;
        RECT 1862.610 1686.780 1862.930 1686.840 ;
        RECT 2105.030 1686.780 2105.350 1686.840 ;
        RECT 1858.010 19.960 1858.330 20.020 ;
        RECT 1862.610 19.960 1862.930 20.020 ;
        RECT 1858.010 19.820 1862.930 19.960 ;
        RECT 1858.010 19.760 1858.330 19.820 ;
        RECT 1862.610 19.760 1862.930 19.820 ;
      LAYER via ;
        RECT 1862.640 1686.780 1862.900 1687.040 ;
        RECT 2105.060 1686.780 2105.320 1687.040 ;
        RECT 1858.040 19.760 1858.300 20.020 ;
        RECT 1862.640 19.760 1862.900 20.020 ;
      LAYER met2 ;
        RECT 2104.980 1700.000 2105.260 1702.400 ;
        RECT 2105.120 1687.070 2105.260 1700.000 ;
        RECT 1862.640 1686.750 1862.900 1687.070 ;
        RECT 2105.060 1686.750 2105.320 1687.070 ;
        RECT 1862.700 20.050 1862.840 1686.750 ;
        RECT 1858.040 19.730 1858.300 20.050 ;
        RECT 1862.640 19.730 1862.900 20.050 ;
        RECT 1858.100 2.400 1858.240 19.730 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2047.605 15.385 2047.775 16.915 ;
      LAYER mcon ;
        RECT 2047.605 16.745 2047.775 16.915 ;
      LAYER met1 ;
        RECT 2073.290 1685.620 2073.610 1685.680 ;
        RECT 2114.230 1685.620 2114.550 1685.680 ;
        RECT 2073.290 1685.480 2114.550 1685.620 ;
        RECT 2073.290 1685.420 2073.610 1685.480 ;
        RECT 2114.230 1685.420 2114.550 1685.480 ;
        RECT 2047.545 16.900 2047.835 16.945 ;
        RECT 2018.640 16.760 2047.835 16.900 ;
        RECT 2018.640 16.560 2018.780 16.760 ;
        RECT 2047.545 16.715 2047.835 16.760 ;
        RECT 2017.720 16.420 2018.780 16.560 ;
        RECT 2017.720 16.220 2017.860 16.420 ;
        RECT 2017.260 16.080 2017.860 16.220 ;
        RECT 1875.950 15.540 1876.270 15.600 ;
        RECT 2017.260 15.540 2017.400 16.080 ;
        RECT 1875.950 15.400 2017.400 15.540 ;
        RECT 2047.545 15.540 2047.835 15.585 ;
        RECT 2073.290 15.540 2073.610 15.600 ;
        RECT 2047.545 15.400 2073.610 15.540 ;
        RECT 1875.950 15.340 1876.270 15.400 ;
        RECT 2047.545 15.355 2047.835 15.400 ;
        RECT 2073.290 15.340 2073.610 15.400 ;
      LAYER via ;
        RECT 2073.320 1685.420 2073.580 1685.680 ;
        RECT 2114.260 1685.420 2114.520 1685.680 ;
        RECT 1875.980 15.340 1876.240 15.600 ;
        RECT 2073.320 15.340 2073.580 15.600 ;
      LAYER met2 ;
        RECT 2114.180 1700.000 2114.460 1702.400 ;
        RECT 2114.320 1685.710 2114.460 1700.000 ;
        RECT 2073.320 1685.390 2073.580 1685.710 ;
        RECT 2114.260 1685.390 2114.520 1685.710 ;
        RECT 2073.380 15.630 2073.520 1685.390 ;
        RECT 1875.980 15.310 1876.240 15.630 ;
        RECT 2073.320 15.310 2073.580 15.630 ;
        RECT 1876.040 2.400 1876.180 15.310 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1531.870 1678.140 1532.190 1678.200 ;
        RECT 1533.710 1678.140 1534.030 1678.200 ;
        RECT 1531.870 1678.000 1534.030 1678.140 ;
        RECT 1531.870 1677.940 1532.190 1678.000 ;
        RECT 1533.710 1677.940 1534.030 1678.000 ;
        RECT 758.150 50.900 758.470 50.960 ;
        RECT 1531.870 50.900 1532.190 50.960 ;
        RECT 758.150 50.760 1532.190 50.900 ;
        RECT 758.150 50.700 758.470 50.760 ;
        RECT 1531.870 50.700 1532.190 50.760 ;
        RECT 752.170 20.980 752.490 21.040 ;
        RECT 758.150 20.980 758.470 21.040 ;
        RECT 752.170 20.840 758.470 20.980 ;
        RECT 752.170 20.780 752.490 20.840 ;
        RECT 758.150 20.780 758.470 20.840 ;
      LAYER via ;
        RECT 1531.900 1677.940 1532.160 1678.200 ;
        RECT 1533.740 1677.940 1534.000 1678.200 ;
        RECT 758.180 50.700 758.440 50.960 ;
        RECT 1531.900 50.700 1532.160 50.960 ;
        RECT 752.200 20.780 752.460 21.040 ;
        RECT 758.180 20.780 758.440 21.040 ;
      LAYER met2 ;
        RECT 1535.500 1700.410 1535.780 1702.400 ;
        RECT 1533.800 1700.270 1535.780 1700.410 ;
        RECT 1533.800 1678.230 1533.940 1700.270 ;
        RECT 1535.500 1700.000 1535.780 1700.270 ;
        RECT 1531.900 1677.910 1532.160 1678.230 ;
        RECT 1533.740 1677.910 1534.000 1678.230 ;
        RECT 1531.960 50.990 1532.100 1677.910 ;
        RECT 758.180 50.670 758.440 50.990 ;
        RECT 1531.900 50.670 1532.160 50.990 ;
        RECT 758.240 21.070 758.380 50.670 ;
        RECT 752.200 20.750 752.460 21.070 ;
        RECT 758.180 20.750 758.440 21.070 ;
        RECT 752.260 2.400 752.400 20.750 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2123.430 1684.260 2123.750 1684.320 ;
        RECT 2115.240 1684.120 2123.750 1684.260 ;
        RECT 2080.650 1683.920 2080.970 1683.980 ;
        RECT 2115.240 1683.920 2115.380 1684.120 ;
        RECT 2123.430 1684.060 2123.750 1684.120 ;
        RECT 2080.650 1683.780 2115.380 1683.920 ;
        RECT 2080.650 1683.720 2080.970 1683.780 ;
        RECT 1894.350 15.200 1894.670 15.260 ;
        RECT 1894.350 15.060 2046.840 15.200 ;
        RECT 1894.350 15.000 1894.670 15.060 ;
        RECT 2046.700 14.520 2046.840 15.060 ;
        RECT 2080.190 14.520 2080.510 14.580 ;
        RECT 2046.700 14.380 2080.510 14.520 ;
        RECT 2080.190 14.320 2080.510 14.380 ;
      LAYER via ;
        RECT 2080.680 1683.720 2080.940 1683.980 ;
        RECT 2123.460 1684.060 2123.720 1684.320 ;
        RECT 1894.380 15.000 1894.640 15.260 ;
        RECT 2080.220 14.320 2080.480 14.580 ;
      LAYER met2 ;
        RECT 2123.380 1700.000 2123.660 1702.400 ;
        RECT 2123.520 1684.350 2123.660 1700.000 ;
        RECT 2123.460 1684.030 2123.720 1684.350 ;
        RECT 2080.680 1683.690 2080.940 1684.010 ;
        RECT 1894.380 14.970 1894.640 15.290 ;
        RECT 1894.440 7.890 1894.580 14.970 ;
        RECT 2080.740 14.690 2080.880 1683.690 ;
        RECT 2080.280 14.610 2080.880 14.690 ;
        RECT 2080.220 14.550 2080.880 14.610 ;
        RECT 2080.220 14.290 2080.480 14.550 ;
        RECT 1893.980 7.750 1894.580 7.890 ;
        RECT 1893.980 2.400 1894.120 7.750 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2094.525 14.705 2094.695 17.595 ;
      LAYER mcon ;
        RECT 2094.525 17.425 2094.695 17.595 ;
      LAYER met1 ;
        RECT 1911.830 17.580 1912.150 17.640 ;
        RECT 2094.465 17.580 2094.755 17.625 ;
        RECT 1911.830 17.440 2094.755 17.580 ;
        RECT 1911.830 17.380 1912.150 17.440 ;
        RECT 2094.465 17.395 2094.755 17.440 ;
        RECT 2094.465 14.860 2094.755 14.905 ;
        RECT 2133.090 14.860 2133.410 14.920 ;
        RECT 2094.465 14.720 2133.410 14.860 ;
        RECT 2094.465 14.675 2094.755 14.720 ;
        RECT 2133.090 14.660 2133.410 14.720 ;
      LAYER via ;
        RECT 1911.860 17.380 1912.120 17.640 ;
        RECT 2133.120 14.660 2133.380 14.920 ;
      LAYER met2 ;
        RECT 2132.580 1700.410 2132.860 1702.400 ;
        RECT 2132.580 1700.270 2133.320 1700.410 ;
        RECT 2132.580 1700.000 2132.860 1700.270 ;
        RECT 1911.860 17.350 1912.120 17.670 ;
        RECT 1911.920 2.400 1912.060 17.350 ;
        RECT 2133.180 14.950 2133.320 1700.270 ;
        RECT 2133.120 14.630 2133.380 14.950 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2016.325 18.445 2016.495 21.675 ;
        RECT 2042.085 19.805 2042.255 21.675 ;
      LAYER mcon ;
        RECT 2016.325 21.505 2016.495 21.675 ;
        RECT 2042.085 21.505 2042.255 21.675 ;
      LAYER met1 ;
        RECT 2045.690 1686.640 2046.010 1686.700 ;
        RECT 2141.830 1686.640 2142.150 1686.700 ;
        RECT 2045.690 1686.500 2142.150 1686.640 ;
        RECT 2045.690 1686.440 2046.010 1686.500 ;
        RECT 2141.830 1686.440 2142.150 1686.500 ;
        RECT 2016.265 21.660 2016.555 21.705 ;
        RECT 2042.025 21.660 2042.315 21.705 ;
        RECT 2016.265 21.520 2042.315 21.660 ;
        RECT 2016.265 21.475 2016.555 21.520 ;
        RECT 2042.025 21.475 2042.315 21.520 ;
        RECT 2045.690 20.300 2046.010 20.360 ;
        RECT 2043.020 20.160 2046.010 20.300 ;
        RECT 2042.025 19.960 2042.315 20.005 ;
        RECT 2043.020 19.960 2043.160 20.160 ;
        RECT 2045.690 20.100 2046.010 20.160 ;
        RECT 2042.025 19.820 2043.160 19.960 ;
        RECT 2042.025 19.775 2042.315 19.820 ;
        RECT 1929.310 18.600 1929.630 18.660 ;
        RECT 2016.265 18.600 2016.555 18.645 ;
        RECT 1929.310 18.460 2016.555 18.600 ;
        RECT 1929.310 18.400 1929.630 18.460 ;
        RECT 2016.265 18.415 2016.555 18.460 ;
      LAYER via ;
        RECT 2045.720 1686.440 2045.980 1686.700 ;
        RECT 2141.860 1686.440 2142.120 1686.700 ;
        RECT 2045.720 20.100 2045.980 20.360 ;
        RECT 1929.340 18.400 1929.600 18.660 ;
      LAYER met2 ;
        RECT 2141.780 1700.000 2142.060 1702.400 ;
        RECT 2141.920 1686.730 2142.060 1700.000 ;
        RECT 2045.720 1686.410 2045.980 1686.730 ;
        RECT 2141.860 1686.410 2142.120 1686.730 ;
        RECT 2045.780 20.390 2045.920 1686.410 ;
        RECT 2045.720 20.070 2045.980 20.390 ;
        RECT 1929.340 18.370 1929.600 18.690 ;
        RECT 1929.400 2.400 1929.540 18.370 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2125.345 17.425 2125.515 20.655 ;
      LAYER mcon ;
        RECT 2125.345 20.485 2125.515 20.655 ;
      LAYER met1 ;
        RECT 2125.285 20.640 2125.575 20.685 ;
        RECT 2146.430 20.640 2146.750 20.700 ;
        RECT 2125.285 20.500 2146.750 20.640 ;
        RECT 2125.285 20.455 2125.575 20.500 ;
        RECT 2146.430 20.440 2146.750 20.500 ;
        RECT 1947.250 17.920 1947.570 17.980 ;
        RECT 1947.250 17.780 2114.460 17.920 ;
        RECT 1947.250 17.720 1947.570 17.780 ;
        RECT 2114.320 17.580 2114.460 17.780 ;
        RECT 2125.285 17.580 2125.575 17.625 ;
        RECT 2114.320 17.440 2125.575 17.580 ;
        RECT 2125.285 17.395 2125.575 17.440 ;
      LAYER via ;
        RECT 2146.460 20.440 2146.720 20.700 ;
        RECT 1947.280 17.720 1947.540 17.980 ;
      LAYER met2 ;
        RECT 2150.980 1700.410 2151.260 1702.400 ;
        RECT 2148.820 1700.270 2151.260 1700.410 ;
        RECT 2148.820 1656.210 2148.960 1700.270 ;
        RECT 2150.980 1700.000 2151.260 1700.270 ;
        RECT 2146.520 1656.070 2148.960 1656.210 ;
        RECT 2146.520 20.730 2146.660 1656.070 ;
        RECT 2146.460 20.410 2146.720 20.730 ;
        RECT 1947.280 17.690 1947.540 18.010 ;
        RECT 1947.340 2.400 1947.480 17.690 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1965.725 1635.485 1965.895 1656.395 ;
        RECT 1966.185 1545.725 1966.355 1621.035 ;
        RECT 1966.185 1352.605 1966.355 1400.715 ;
        RECT 1966.185 676.345 1966.355 724.455 ;
        RECT 1966.185 579.785 1966.355 627.895 ;
        RECT 1966.185 427.805 1966.355 475.915 ;
        RECT 1966.185 289.765 1966.355 337.875 ;
        RECT 1966.185 96.645 1966.355 144.755 ;
        RECT 1965.265 2.805 1965.435 48.195 ;
      LAYER mcon ;
        RECT 1965.725 1656.225 1965.895 1656.395 ;
        RECT 1966.185 1620.865 1966.355 1621.035 ;
        RECT 1966.185 1400.545 1966.355 1400.715 ;
        RECT 1966.185 724.285 1966.355 724.455 ;
        RECT 1966.185 627.725 1966.355 627.895 ;
        RECT 1966.185 475.745 1966.355 475.915 ;
        RECT 1966.185 337.705 1966.355 337.875 ;
        RECT 1966.185 144.585 1966.355 144.755 ;
        RECT 1965.265 48.025 1965.435 48.195 ;
      LAYER met1 ;
        RECT 1965.650 1688.000 1965.970 1688.060 ;
        RECT 2160.230 1688.000 2160.550 1688.060 ;
        RECT 1965.650 1687.860 2160.550 1688.000 ;
        RECT 1965.650 1687.800 1965.970 1687.860 ;
        RECT 2160.230 1687.800 2160.550 1687.860 ;
        RECT 1965.650 1656.380 1965.970 1656.440 ;
        RECT 1965.455 1656.240 1965.970 1656.380 ;
        RECT 1965.650 1656.180 1965.970 1656.240 ;
        RECT 1965.190 1635.640 1965.510 1635.700 ;
        RECT 1965.665 1635.640 1965.955 1635.685 ;
        RECT 1965.190 1635.500 1965.955 1635.640 ;
        RECT 1965.190 1635.440 1965.510 1635.500 ;
        RECT 1965.665 1635.455 1965.955 1635.500 ;
        RECT 1965.190 1621.020 1965.510 1621.080 ;
        RECT 1966.125 1621.020 1966.415 1621.065 ;
        RECT 1965.190 1620.880 1966.415 1621.020 ;
        RECT 1965.190 1620.820 1965.510 1620.880 ;
        RECT 1966.125 1620.835 1966.415 1620.880 ;
        RECT 1966.110 1545.880 1966.430 1545.940 ;
        RECT 1965.915 1545.740 1966.430 1545.880 ;
        RECT 1966.110 1545.680 1966.430 1545.740 ;
        RECT 1966.110 1400.700 1966.430 1400.760 ;
        RECT 1965.915 1400.560 1966.430 1400.700 ;
        RECT 1966.110 1400.500 1966.430 1400.560 ;
        RECT 1966.110 1352.760 1966.430 1352.820 ;
        RECT 1965.915 1352.620 1966.430 1352.760 ;
        RECT 1966.110 1352.560 1966.430 1352.620 ;
        RECT 1965.650 1159.300 1965.970 1159.360 ;
        RECT 1966.110 1159.300 1966.430 1159.360 ;
        RECT 1965.650 1159.160 1966.430 1159.300 ;
        RECT 1965.650 1159.100 1965.970 1159.160 ;
        RECT 1966.110 1159.100 1966.430 1159.160 ;
        RECT 1966.110 1111.020 1966.430 1111.080 ;
        RECT 1967.030 1111.020 1967.350 1111.080 ;
        RECT 1966.110 1110.880 1967.350 1111.020 ;
        RECT 1966.110 1110.820 1966.430 1110.880 ;
        RECT 1967.030 1110.820 1967.350 1110.880 ;
        RECT 1965.650 1062.740 1965.970 1062.800 ;
        RECT 1966.110 1062.740 1966.430 1062.800 ;
        RECT 1965.650 1062.600 1966.430 1062.740 ;
        RECT 1965.650 1062.540 1965.970 1062.600 ;
        RECT 1966.110 1062.540 1966.430 1062.600 ;
        RECT 1966.110 1014.460 1966.430 1014.520 ;
        RECT 1967.030 1014.460 1967.350 1014.520 ;
        RECT 1966.110 1014.320 1967.350 1014.460 ;
        RECT 1966.110 1014.260 1966.430 1014.320 ;
        RECT 1967.030 1014.260 1967.350 1014.320 ;
        RECT 1965.650 966.180 1965.970 966.240 ;
        RECT 1966.110 966.180 1966.430 966.240 ;
        RECT 1965.650 966.040 1966.430 966.180 ;
        RECT 1965.650 965.980 1965.970 966.040 ;
        RECT 1966.110 965.980 1966.430 966.040 ;
        RECT 1966.110 917.900 1966.430 917.960 ;
        RECT 1967.030 917.900 1967.350 917.960 ;
        RECT 1966.110 917.760 1967.350 917.900 ;
        RECT 1966.110 917.700 1966.430 917.760 ;
        RECT 1967.030 917.700 1967.350 917.760 ;
        RECT 1966.110 772.720 1966.430 772.780 ;
        RECT 1967.030 772.720 1967.350 772.780 ;
        RECT 1966.110 772.580 1967.350 772.720 ;
        RECT 1966.110 772.520 1966.430 772.580 ;
        RECT 1967.030 772.520 1967.350 772.580 ;
        RECT 1966.110 724.440 1966.430 724.500 ;
        RECT 1965.915 724.300 1966.430 724.440 ;
        RECT 1966.110 724.240 1966.430 724.300 ;
        RECT 1966.110 676.500 1966.430 676.560 ;
        RECT 1965.915 676.360 1966.430 676.500 ;
        RECT 1966.110 676.300 1966.430 676.360 ;
        RECT 1966.110 627.880 1966.430 627.940 ;
        RECT 1965.915 627.740 1966.430 627.880 ;
        RECT 1966.110 627.680 1966.430 627.740 ;
        RECT 1966.110 579.940 1966.430 580.000 ;
        RECT 1965.915 579.800 1966.430 579.940 ;
        RECT 1966.110 579.740 1966.430 579.800 ;
        RECT 1966.110 579.260 1966.430 579.320 ;
        RECT 1966.570 579.260 1966.890 579.320 ;
        RECT 1966.110 579.120 1966.890 579.260 ;
        RECT 1966.110 579.060 1966.430 579.120 ;
        RECT 1966.570 579.060 1966.890 579.120 ;
        RECT 1966.110 531.320 1966.430 531.380 ;
        RECT 1967.030 531.320 1967.350 531.380 ;
        RECT 1966.110 531.180 1967.350 531.320 ;
        RECT 1966.110 531.120 1966.430 531.180 ;
        RECT 1967.030 531.120 1967.350 531.180 ;
        RECT 1966.110 475.900 1966.430 475.960 ;
        RECT 1965.915 475.760 1966.430 475.900 ;
        RECT 1966.110 475.700 1966.430 475.760 ;
        RECT 1966.125 427.960 1966.415 428.005 ;
        RECT 1967.030 427.960 1967.350 428.020 ;
        RECT 1966.125 427.820 1967.350 427.960 ;
        RECT 1966.125 427.775 1966.415 427.820 ;
        RECT 1967.030 427.760 1967.350 427.820 ;
        RECT 1966.110 337.860 1966.430 337.920 ;
        RECT 1965.915 337.720 1966.430 337.860 ;
        RECT 1966.110 337.660 1966.430 337.720 ;
        RECT 1966.110 289.920 1966.430 289.980 ;
        RECT 1965.915 289.780 1966.430 289.920 ;
        RECT 1966.110 289.720 1966.430 289.780 ;
        RECT 1966.110 144.740 1966.430 144.800 ;
        RECT 1965.915 144.600 1966.430 144.740 ;
        RECT 1966.110 144.540 1966.430 144.600 ;
        RECT 1966.110 96.800 1966.430 96.860 ;
        RECT 1965.915 96.660 1966.430 96.800 ;
        RECT 1966.110 96.600 1966.430 96.660 ;
        RECT 1965.190 48.180 1965.510 48.240 ;
        RECT 1964.995 48.040 1965.510 48.180 ;
        RECT 1965.190 47.980 1965.510 48.040 ;
        RECT 1965.190 2.960 1965.510 3.020 ;
        RECT 1964.995 2.820 1965.510 2.960 ;
        RECT 1965.190 2.760 1965.510 2.820 ;
      LAYER via ;
        RECT 1965.680 1687.800 1965.940 1688.060 ;
        RECT 2160.260 1687.800 2160.520 1688.060 ;
        RECT 1965.680 1656.180 1965.940 1656.440 ;
        RECT 1965.220 1635.440 1965.480 1635.700 ;
        RECT 1965.220 1620.820 1965.480 1621.080 ;
        RECT 1966.140 1545.680 1966.400 1545.940 ;
        RECT 1966.140 1400.500 1966.400 1400.760 ;
        RECT 1966.140 1352.560 1966.400 1352.820 ;
        RECT 1965.680 1159.100 1965.940 1159.360 ;
        RECT 1966.140 1159.100 1966.400 1159.360 ;
        RECT 1966.140 1110.820 1966.400 1111.080 ;
        RECT 1967.060 1110.820 1967.320 1111.080 ;
        RECT 1965.680 1062.540 1965.940 1062.800 ;
        RECT 1966.140 1062.540 1966.400 1062.800 ;
        RECT 1966.140 1014.260 1966.400 1014.520 ;
        RECT 1967.060 1014.260 1967.320 1014.520 ;
        RECT 1965.680 965.980 1965.940 966.240 ;
        RECT 1966.140 965.980 1966.400 966.240 ;
        RECT 1966.140 917.700 1966.400 917.960 ;
        RECT 1967.060 917.700 1967.320 917.960 ;
        RECT 1966.140 772.520 1966.400 772.780 ;
        RECT 1967.060 772.520 1967.320 772.780 ;
        RECT 1966.140 724.240 1966.400 724.500 ;
        RECT 1966.140 676.300 1966.400 676.560 ;
        RECT 1966.140 627.680 1966.400 627.940 ;
        RECT 1966.140 579.740 1966.400 580.000 ;
        RECT 1966.140 579.060 1966.400 579.320 ;
        RECT 1966.600 579.060 1966.860 579.320 ;
        RECT 1966.140 531.120 1966.400 531.380 ;
        RECT 1967.060 531.120 1967.320 531.380 ;
        RECT 1966.140 475.700 1966.400 475.960 ;
        RECT 1967.060 427.760 1967.320 428.020 ;
        RECT 1966.140 337.660 1966.400 337.920 ;
        RECT 1966.140 289.720 1966.400 289.980 ;
        RECT 1966.140 144.540 1966.400 144.800 ;
        RECT 1966.140 96.600 1966.400 96.860 ;
        RECT 1965.220 47.980 1965.480 48.240 ;
        RECT 1965.220 2.760 1965.480 3.020 ;
      LAYER met2 ;
        RECT 2160.180 1700.000 2160.460 1702.400 ;
        RECT 2160.320 1688.090 2160.460 1700.000 ;
        RECT 1965.680 1687.770 1965.940 1688.090 ;
        RECT 2160.260 1687.770 2160.520 1688.090 ;
        RECT 1965.740 1656.470 1965.880 1687.770 ;
        RECT 1965.680 1656.150 1965.940 1656.470 ;
        RECT 1965.220 1635.410 1965.480 1635.730 ;
        RECT 1965.280 1621.110 1965.420 1635.410 ;
        RECT 1965.220 1620.790 1965.480 1621.110 ;
        RECT 1966.140 1545.650 1966.400 1545.970 ;
        RECT 1966.200 1400.790 1966.340 1545.650 ;
        RECT 1966.140 1400.470 1966.400 1400.790 ;
        RECT 1966.140 1352.530 1966.400 1352.850 ;
        RECT 1966.200 1207.410 1966.340 1352.530 ;
        RECT 1965.740 1207.270 1966.340 1207.410 ;
        RECT 1965.740 1159.390 1965.880 1207.270 ;
        RECT 1965.680 1159.070 1965.940 1159.390 ;
        RECT 1966.140 1159.245 1966.400 1159.390 ;
        RECT 1966.130 1158.875 1966.410 1159.245 ;
        RECT 1967.050 1158.875 1967.330 1159.245 ;
        RECT 1966.200 1111.110 1966.340 1111.265 ;
        RECT 1967.120 1111.110 1967.260 1158.875 ;
        RECT 1966.140 1110.850 1966.400 1111.110 ;
        RECT 1965.740 1110.790 1966.400 1110.850 ;
        RECT 1967.060 1110.790 1967.320 1111.110 ;
        RECT 1965.740 1110.710 1966.340 1110.790 ;
        RECT 1965.740 1062.830 1965.880 1110.710 ;
        RECT 1965.680 1062.510 1965.940 1062.830 ;
        RECT 1966.140 1062.685 1966.400 1062.830 ;
        RECT 1966.130 1062.315 1966.410 1062.685 ;
        RECT 1967.050 1062.315 1967.330 1062.685 ;
        RECT 1966.200 1014.550 1966.340 1014.705 ;
        RECT 1967.120 1014.550 1967.260 1062.315 ;
        RECT 1966.140 1014.290 1966.400 1014.550 ;
        RECT 1965.740 1014.230 1966.400 1014.290 ;
        RECT 1967.060 1014.230 1967.320 1014.550 ;
        RECT 1965.740 1014.150 1966.340 1014.230 ;
        RECT 1965.740 966.270 1965.880 1014.150 ;
        RECT 1965.680 965.950 1965.940 966.270 ;
        RECT 1966.140 966.125 1966.400 966.270 ;
        RECT 1966.130 965.755 1966.410 966.125 ;
        RECT 1967.050 965.755 1967.330 966.125 ;
        RECT 1967.120 917.990 1967.260 965.755 ;
        RECT 1966.140 917.670 1966.400 917.990 ;
        RECT 1967.060 917.670 1967.320 917.990 ;
        RECT 1966.200 772.810 1966.340 917.670 ;
        RECT 1966.140 772.490 1966.400 772.810 ;
        RECT 1967.060 772.490 1967.320 772.810 ;
        RECT 1967.120 724.725 1967.260 772.490 ;
        RECT 1966.130 724.355 1966.410 724.725 ;
        RECT 1967.050 724.355 1967.330 724.725 ;
        RECT 1966.140 724.210 1966.400 724.355 ;
        RECT 1966.140 676.270 1966.400 676.590 ;
        RECT 1966.200 627.970 1966.340 676.270 ;
        RECT 1966.140 627.650 1966.400 627.970 ;
        RECT 1966.140 579.710 1966.400 580.030 ;
        RECT 1966.200 579.350 1966.340 579.710 ;
        RECT 1966.140 579.030 1966.400 579.350 ;
        RECT 1966.600 579.030 1966.860 579.350 ;
        RECT 1966.660 531.490 1966.800 579.030 ;
        RECT 1966.200 531.410 1966.800 531.490 ;
        RECT 1966.140 531.350 1966.800 531.410 ;
        RECT 1966.140 531.090 1966.400 531.350 ;
        RECT 1967.060 531.090 1967.320 531.410 ;
        RECT 1967.120 483.325 1967.260 531.090 ;
        RECT 1966.130 482.955 1966.410 483.325 ;
        RECT 1967.050 482.955 1967.330 483.325 ;
        RECT 1966.200 475.990 1966.340 482.955 ;
        RECT 1966.140 475.670 1966.400 475.990 ;
        RECT 1967.060 427.730 1967.320 428.050 ;
        RECT 1967.120 339.165 1967.260 427.730 ;
        RECT 1967.050 338.795 1967.330 339.165 ;
        RECT 1966.130 338.115 1966.410 338.485 ;
        RECT 1966.200 337.950 1966.340 338.115 ;
        RECT 1966.140 337.630 1966.400 337.950 ;
        RECT 1966.140 289.690 1966.400 290.010 ;
        RECT 1966.200 144.830 1966.340 289.690 ;
        RECT 1966.140 144.510 1966.400 144.830 ;
        RECT 1966.140 96.570 1966.400 96.890 ;
        RECT 1966.200 72.490 1966.340 96.570 ;
        RECT 1965.280 72.350 1966.340 72.490 ;
        RECT 1965.280 48.270 1965.420 72.350 ;
        RECT 1965.220 47.950 1965.480 48.270 ;
        RECT 1965.220 2.730 1965.480 3.050 ;
        RECT 1965.280 2.400 1965.420 2.730 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
      LAYER via2 ;
        RECT 1966.130 1158.920 1966.410 1159.200 ;
        RECT 1967.050 1158.920 1967.330 1159.200 ;
        RECT 1966.130 1062.360 1966.410 1062.640 ;
        RECT 1967.050 1062.360 1967.330 1062.640 ;
        RECT 1966.130 965.800 1966.410 966.080 ;
        RECT 1967.050 965.800 1967.330 966.080 ;
        RECT 1966.130 724.400 1966.410 724.680 ;
        RECT 1967.050 724.400 1967.330 724.680 ;
        RECT 1966.130 483.000 1966.410 483.280 ;
        RECT 1967.050 483.000 1967.330 483.280 ;
        RECT 1967.050 338.840 1967.330 339.120 ;
        RECT 1966.130 338.160 1966.410 338.440 ;
      LAYER met3 ;
        RECT 1966.105 1159.210 1966.435 1159.225 ;
        RECT 1967.025 1159.210 1967.355 1159.225 ;
        RECT 1966.105 1158.910 1967.355 1159.210 ;
        RECT 1966.105 1158.895 1966.435 1158.910 ;
        RECT 1967.025 1158.895 1967.355 1158.910 ;
        RECT 1966.105 1062.650 1966.435 1062.665 ;
        RECT 1967.025 1062.650 1967.355 1062.665 ;
        RECT 1966.105 1062.350 1967.355 1062.650 ;
        RECT 1966.105 1062.335 1966.435 1062.350 ;
        RECT 1967.025 1062.335 1967.355 1062.350 ;
        RECT 1966.105 966.090 1966.435 966.105 ;
        RECT 1967.025 966.090 1967.355 966.105 ;
        RECT 1966.105 965.790 1967.355 966.090 ;
        RECT 1966.105 965.775 1966.435 965.790 ;
        RECT 1967.025 965.775 1967.355 965.790 ;
        RECT 1966.105 724.690 1966.435 724.705 ;
        RECT 1967.025 724.690 1967.355 724.705 ;
        RECT 1966.105 724.390 1967.355 724.690 ;
        RECT 1966.105 724.375 1966.435 724.390 ;
        RECT 1967.025 724.375 1967.355 724.390 ;
        RECT 1966.105 483.290 1966.435 483.305 ;
        RECT 1967.025 483.290 1967.355 483.305 ;
        RECT 1966.105 482.990 1967.355 483.290 ;
        RECT 1966.105 482.975 1966.435 482.990 ;
        RECT 1967.025 482.975 1967.355 482.990 ;
        RECT 1967.025 339.130 1967.355 339.145 ;
        RECT 1965.430 338.830 1967.355 339.130 ;
        RECT 1965.430 338.450 1965.730 338.830 ;
        RECT 1967.025 338.815 1967.355 338.830 ;
        RECT 1966.105 338.450 1966.435 338.465 ;
        RECT 1965.430 338.150 1966.435 338.450 ;
        RECT 1966.105 338.135 1966.435 338.150 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2042.085 17.085 2042.255 18.275 ;
        RECT 2068.305 17.085 2068.475 20.655 ;
        RECT 2090.385 17.085 2090.555 18.615 ;
      LAYER mcon ;
        RECT 2068.305 20.485 2068.475 20.655 ;
        RECT 2042.085 18.105 2042.255 18.275 ;
        RECT 2090.385 18.445 2090.555 18.615 ;
      LAYER met1 ;
        RECT 2042.930 20.980 2043.250 21.040 ;
        RECT 2042.930 20.840 2063.400 20.980 ;
        RECT 2042.930 20.780 2043.250 20.840 ;
        RECT 2063.260 20.640 2063.400 20.840 ;
        RECT 2068.245 20.640 2068.535 20.685 ;
        RECT 2063.260 20.500 2068.535 20.640 ;
        RECT 2068.245 20.455 2068.535 20.500 ;
        RECT 2090.325 18.600 2090.615 18.645 ;
        RECT 2090.325 18.460 2114.920 18.600 ;
        RECT 2090.325 18.415 2090.615 18.460 ;
        RECT 2042.025 18.260 2042.315 18.305 ;
        RECT 2042.470 18.260 2042.790 18.320 ;
        RECT 2042.025 18.120 2042.790 18.260 ;
        RECT 2042.025 18.075 2042.315 18.120 ;
        RECT 2042.470 18.060 2042.790 18.120 ;
        RECT 2114.780 17.920 2114.920 18.460 ;
        RECT 2166.670 17.920 2166.990 17.980 ;
        RECT 2114.780 17.780 2166.990 17.920 ;
        RECT 2166.670 17.720 2166.990 17.780 ;
        RECT 2042.025 17.240 2042.315 17.285 ;
        RECT 2018.180 17.100 2042.315 17.240 ;
        RECT 1983.130 16.900 1983.450 16.960 ;
        RECT 2018.180 16.900 2018.320 17.100 ;
        RECT 2042.025 17.055 2042.315 17.100 ;
        RECT 2068.245 17.240 2068.535 17.285 ;
        RECT 2090.325 17.240 2090.615 17.285 ;
        RECT 2068.245 17.100 2090.615 17.240 ;
        RECT 2068.245 17.055 2068.535 17.100 ;
        RECT 2090.325 17.055 2090.615 17.100 ;
        RECT 1983.130 16.760 2018.320 16.900 ;
        RECT 1983.130 16.700 1983.450 16.760 ;
      LAYER via ;
        RECT 2042.960 20.780 2043.220 21.040 ;
        RECT 2042.500 18.060 2042.760 18.320 ;
        RECT 2166.700 17.720 2166.960 17.980 ;
        RECT 1983.160 16.700 1983.420 16.960 ;
      LAYER met2 ;
        RECT 2169.380 1700.410 2169.660 1702.400 ;
        RECT 2166.760 1700.270 2169.660 1700.410 ;
        RECT 2042.960 20.810 2043.220 21.070 ;
        RECT 2042.560 20.750 2043.220 20.810 ;
        RECT 2042.560 20.670 2043.160 20.750 ;
        RECT 2042.560 18.350 2042.700 20.670 ;
        RECT 2042.500 18.030 2042.760 18.350 ;
        RECT 2166.760 18.010 2166.900 1700.270 ;
        RECT 2169.380 1700.000 2169.660 1700.270 ;
        RECT 2166.700 17.690 2166.960 18.010 ;
        RECT 1983.160 16.670 1983.420 16.990 ;
        RECT 1983.220 2.400 1983.360 16.670 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2115.225 18.105 2115.395 19.635 ;
      LAYER mcon ;
        RECT 2115.225 19.465 2115.395 19.635 ;
      LAYER met1 ;
        RECT 2162.990 1683.920 2163.310 1683.980 ;
        RECT 2178.630 1683.920 2178.950 1683.980 ;
        RECT 2162.990 1683.780 2178.950 1683.920 ;
        RECT 2162.990 1683.720 2163.310 1683.780 ;
        RECT 2178.630 1683.720 2178.950 1683.780 ;
        RECT 2001.070 20.640 2001.390 20.700 ;
        RECT 2042.010 20.640 2042.330 20.700 ;
        RECT 2001.070 20.500 2042.330 20.640 ;
        RECT 2001.070 20.440 2001.390 20.500 ;
        RECT 2042.010 20.440 2042.330 20.500 ;
        RECT 2042.930 19.620 2043.250 19.680 ;
        RECT 2115.165 19.620 2115.455 19.665 ;
        RECT 2042.930 19.480 2115.455 19.620 ;
        RECT 2042.930 19.420 2043.250 19.480 ;
        RECT 2115.165 19.435 2115.455 19.480 ;
        RECT 2115.165 18.260 2115.455 18.305 ;
        RECT 2162.990 18.260 2163.310 18.320 ;
        RECT 2115.165 18.120 2163.310 18.260 ;
        RECT 2115.165 18.075 2115.455 18.120 ;
        RECT 2162.990 18.060 2163.310 18.120 ;
      LAYER via ;
        RECT 2163.020 1683.720 2163.280 1683.980 ;
        RECT 2178.660 1683.720 2178.920 1683.980 ;
        RECT 2001.100 20.440 2001.360 20.700 ;
        RECT 2042.040 20.440 2042.300 20.700 ;
        RECT 2042.960 19.420 2043.220 19.680 ;
        RECT 2163.020 18.060 2163.280 18.320 ;
      LAYER met2 ;
        RECT 2178.580 1700.000 2178.860 1702.400 ;
        RECT 2178.720 1684.010 2178.860 1700.000 ;
        RECT 2163.020 1683.690 2163.280 1684.010 ;
        RECT 2178.660 1683.690 2178.920 1684.010 ;
        RECT 2001.100 20.410 2001.360 20.730 ;
        RECT 2042.040 20.410 2042.300 20.730 ;
        RECT 2001.160 2.400 2001.300 20.410 ;
        RECT 2042.100 19.565 2042.240 20.410 ;
        RECT 2042.960 19.565 2043.220 19.710 ;
        RECT 2042.030 19.195 2042.310 19.565 ;
        RECT 2042.950 19.195 2043.230 19.565 ;
        RECT 2163.080 18.350 2163.220 1683.690 ;
        RECT 2163.020 18.030 2163.280 18.350 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
      LAYER via2 ;
        RECT 2042.030 19.240 2042.310 19.520 ;
        RECT 2042.950 19.240 2043.230 19.520 ;
      LAYER met3 ;
        RECT 2042.005 19.530 2042.335 19.545 ;
        RECT 2042.925 19.530 2043.255 19.545 ;
        RECT 2042.005 19.230 2043.255 19.530 ;
        RECT 2042.005 19.215 2042.335 19.230 ;
        RECT 2042.925 19.215 2043.255 19.230 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2018.550 19.280 2018.870 19.340 ;
        RECT 2188.290 19.280 2188.610 19.340 ;
        RECT 2018.550 19.140 2188.610 19.280 ;
        RECT 2018.550 19.080 2018.870 19.140 ;
        RECT 2188.290 19.080 2188.610 19.140 ;
      LAYER via ;
        RECT 2018.580 19.080 2018.840 19.340 ;
        RECT 2188.320 19.080 2188.580 19.340 ;
      LAYER met2 ;
        RECT 2187.780 1700.410 2188.060 1702.400 ;
        RECT 2187.780 1700.270 2188.520 1700.410 ;
        RECT 2187.780 1700.000 2188.060 1700.270 ;
        RECT 2188.380 19.370 2188.520 1700.270 ;
        RECT 2018.580 19.050 2018.840 19.370 ;
        RECT 2188.320 19.050 2188.580 19.370 ;
        RECT 2018.640 2.400 2018.780 19.050 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2066.925 16.745 2067.095 20.315 ;
      LAYER mcon ;
        RECT 2066.925 20.145 2067.095 20.315 ;
      LAYER met1 ;
        RECT 2066.865 20.300 2067.155 20.345 ;
        RECT 2194.730 20.300 2195.050 20.360 ;
        RECT 2066.865 20.160 2195.050 20.300 ;
        RECT 2066.865 20.115 2067.155 20.160 ;
        RECT 2194.730 20.100 2195.050 20.160 ;
        RECT 2066.865 16.900 2067.155 16.945 ;
        RECT 2048.080 16.760 2067.155 16.900 ;
        RECT 2036.490 16.560 2036.810 16.620 ;
        RECT 2048.080 16.560 2048.220 16.760 ;
        RECT 2066.865 16.715 2067.155 16.760 ;
        RECT 2036.490 16.420 2048.220 16.560 ;
        RECT 2036.490 16.360 2036.810 16.420 ;
      LAYER via ;
        RECT 2194.760 20.100 2195.020 20.360 ;
        RECT 2036.520 16.360 2036.780 16.620 ;
      LAYER met2 ;
        RECT 2196.980 1700.410 2197.260 1702.400 ;
        RECT 2194.820 1700.270 2197.260 1700.410 ;
        RECT 2194.820 20.390 2194.960 1700.270 ;
        RECT 2196.980 1700.000 2197.260 1700.270 ;
        RECT 2194.760 20.070 2195.020 20.390 ;
        RECT 2036.520 16.330 2036.780 16.650 ;
        RECT 2036.580 2.400 2036.720 16.330 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2114.765 1684.105 2114.935 1689.375 ;
      LAYER mcon ;
        RECT 2114.765 1689.205 2114.935 1689.375 ;
      LAYER met1 ;
        RECT 2114.705 1689.360 2114.995 1689.405 ;
        RECT 2206.230 1689.360 2206.550 1689.420 ;
        RECT 2114.705 1689.220 2206.550 1689.360 ;
        RECT 2114.705 1689.175 2114.995 1689.220 ;
        RECT 2206.230 1689.160 2206.550 1689.220 ;
        RECT 2066.390 1684.260 2066.710 1684.320 ;
        RECT 2114.705 1684.260 2114.995 1684.305 ;
        RECT 2066.390 1684.120 2114.995 1684.260 ;
        RECT 2066.390 1684.060 2066.710 1684.120 ;
        RECT 2114.705 1684.075 2114.995 1684.120 ;
        RECT 2054.430 20.300 2054.750 20.360 ;
        RECT 2066.390 20.300 2066.710 20.360 ;
        RECT 2054.430 20.160 2066.710 20.300 ;
        RECT 2054.430 20.100 2054.750 20.160 ;
        RECT 2066.390 20.100 2066.710 20.160 ;
      LAYER via ;
        RECT 2206.260 1689.160 2206.520 1689.420 ;
        RECT 2066.420 1684.060 2066.680 1684.320 ;
        RECT 2054.460 20.100 2054.720 20.360 ;
        RECT 2066.420 20.100 2066.680 20.360 ;
      LAYER met2 ;
        RECT 2206.180 1700.000 2206.460 1702.400 ;
        RECT 2206.320 1689.450 2206.460 1700.000 ;
        RECT 2206.260 1689.130 2206.520 1689.450 ;
        RECT 2066.420 1684.030 2066.680 1684.350 ;
        RECT 2066.480 20.390 2066.620 1684.030 ;
        RECT 2054.460 20.070 2054.720 20.390 ;
        RECT 2066.420 20.070 2066.680 20.390 ;
        RECT 2054.520 2.400 2054.660 20.070 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1540.225 386.325 1540.395 434.775 ;
        RECT 1540.225 289.765 1540.395 337.875 ;
        RECT 1540.685 193.205 1540.855 241.315 ;
        RECT 1540.225 96.645 1540.395 144.755 ;
      LAYER mcon ;
        RECT 1540.225 434.605 1540.395 434.775 ;
        RECT 1540.225 337.705 1540.395 337.875 ;
        RECT 1540.685 241.145 1540.855 241.315 ;
        RECT 1540.225 144.585 1540.395 144.755 ;
      LAYER met1 ;
        RECT 1540.610 869.620 1540.930 869.680 ;
        RECT 1541.530 869.620 1541.850 869.680 ;
        RECT 1540.610 869.480 1541.850 869.620 ;
        RECT 1540.610 869.420 1540.930 869.480 ;
        RECT 1541.530 869.420 1541.850 869.480 ;
        RECT 1540.610 821.000 1540.930 821.060 ;
        RECT 1541.530 821.000 1541.850 821.060 ;
        RECT 1540.610 820.860 1541.850 821.000 ;
        RECT 1540.610 820.800 1540.930 820.860 ;
        RECT 1541.530 820.800 1541.850 820.860 ;
        RECT 1540.610 724.440 1540.930 724.500 ;
        RECT 1541.530 724.440 1541.850 724.500 ;
        RECT 1540.610 724.300 1541.850 724.440 ;
        RECT 1540.610 724.240 1540.930 724.300 ;
        RECT 1541.530 724.240 1541.850 724.300 ;
        RECT 1540.610 627.880 1540.930 627.940 ;
        RECT 1541.530 627.880 1541.850 627.940 ;
        RECT 1540.610 627.740 1541.850 627.880 ;
        RECT 1540.610 627.680 1540.930 627.740 ;
        RECT 1541.530 627.680 1541.850 627.740 ;
        RECT 1540.150 531.320 1540.470 531.380 ;
        RECT 1541.070 531.320 1541.390 531.380 ;
        RECT 1540.150 531.180 1541.390 531.320 ;
        RECT 1540.150 531.120 1540.470 531.180 ;
        RECT 1541.070 531.120 1541.390 531.180 ;
        RECT 1540.150 434.760 1540.470 434.820 ;
        RECT 1539.955 434.620 1540.470 434.760 ;
        RECT 1540.150 434.560 1540.470 434.620 ;
        RECT 1540.150 386.480 1540.470 386.540 ;
        RECT 1539.955 386.340 1540.470 386.480 ;
        RECT 1540.150 386.280 1540.470 386.340 ;
        RECT 1540.150 337.860 1540.470 337.920 ;
        RECT 1539.955 337.720 1540.470 337.860 ;
        RECT 1540.150 337.660 1540.470 337.720 ;
        RECT 1540.150 289.920 1540.470 289.980 ;
        RECT 1539.955 289.780 1540.470 289.920 ;
        RECT 1540.150 289.720 1540.470 289.780 ;
        RECT 1540.610 241.300 1540.930 241.360 ;
        RECT 1540.415 241.160 1540.930 241.300 ;
        RECT 1540.610 241.100 1540.930 241.160 ;
        RECT 1540.610 193.360 1540.930 193.420 ;
        RECT 1540.415 193.220 1540.930 193.360 ;
        RECT 1540.610 193.160 1540.930 193.220 ;
        RECT 1540.165 144.740 1540.455 144.785 ;
        RECT 1540.610 144.740 1540.930 144.800 ;
        RECT 1540.165 144.600 1540.930 144.740 ;
        RECT 1540.165 144.555 1540.455 144.600 ;
        RECT 1540.610 144.540 1540.930 144.600 ;
        RECT 1540.150 96.800 1540.470 96.860 ;
        RECT 1539.955 96.660 1540.470 96.800 ;
        RECT 1540.150 96.600 1540.470 96.660 ;
        RECT 772.410 50.560 772.730 50.620 ;
        RECT 1539.230 50.560 1539.550 50.620 ;
        RECT 772.410 50.420 1539.550 50.560 ;
        RECT 772.410 50.360 772.730 50.420 ;
        RECT 1539.230 50.360 1539.550 50.420 ;
      LAYER via ;
        RECT 1540.640 869.420 1540.900 869.680 ;
        RECT 1541.560 869.420 1541.820 869.680 ;
        RECT 1540.640 820.800 1540.900 821.060 ;
        RECT 1541.560 820.800 1541.820 821.060 ;
        RECT 1540.640 724.240 1540.900 724.500 ;
        RECT 1541.560 724.240 1541.820 724.500 ;
        RECT 1540.640 627.680 1540.900 627.940 ;
        RECT 1541.560 627.680 1541.820 627.940 ;
        RECT 1540.180 531.120 1540.440 531.380 ;
        RECT 1541.100 531.120 1541.360 531.380 ;
        RECT 1540.180 434.560 1540.440 434.820 ;
        RECT 1540.180 386.280 1540.440 386.540 ;
        RECT 1540.180 337.660 1540.440 337.920 ;
        RECT 1540.180 289.720 1540.440 289.980 ;
        RECT 1540.640 241.100 1540.900 241.360 ;
        RECT 1540.640 193.160 1540.900 193.420 ;
        RECT 1540.640 144.540 1540.900 144.800 ;
        RECT 1540.180 96.600 1540.440 96.860 ;
        RECT 772.440 50.360 772.700 50.620 ;
        RECT 1539.260 50.360 1539.520 50.620 ;
      LAYER met2 ;
        RECT 1544.700 1700.410 1544.980 1702.400 ;
        RECT 1542.540 1700.270 1544.980 1700.410 ;
        RECT 1542.540 1656.210 1542.680 1700.270 ;
        RECT 1544.700 1700.000 1544.980 1700.270 ;
        RECT 1540.240 1656.070 1542.680 1656.210 ;
        RECT 1540.240 917.845 1540.380 1656.070 ;
        RECT 1540.170 917.475 1540.450 917.845 ;
        RECT 1541.550 917.475 1541.830 917.845 ;
        RECT 1541.620 869.710 1541.760 917.475 ;
        RECT 1540.640 869.390 1540.900 869.710 ;
        RECT 1541.560 869.390 1541.820 869.710 ;
        RECT 1540.700 821.090 1540.840 869.390 ;
        RECT 1540.640 820.770 1540.900 821.090 ;
        RECT 1541.560 820.770 1541.820 821.090 ;
        RECT 1541.620 773.005 1541.760 820.770 ;
        RECT 1540.170 772.635 1540.450 773.005 ;
        RECT 1541.550 772.635 1541.830 773.005 ;
        RECT 1540.240 738.210 1540.380 772.635 ;
        RECT 1540.240 738.070 1540.840 738.210 ;
        RECT 1540.700 724.530 1540.840 738.070 ;
        RECT 1540.640 724.210 1540.900 724.530 ;
        RECT 1541.560 724.210 1541.820 724.530 ;
        RECT 1541.620 676.445 1541.760 724.210 ;
        RECT 1540.630 676.075 1540.910 676.445 ;
        RECT 1541.550 676.075 1541.830 676.445 ;
        RECT 1540.700 627.970 1540.840 676.075 ;
        RECT 1540.640 627.650 1540.900 627.970 ;
        RECT 1541.560 627.650 1541.820 627.970 ;
        RECT 1541.620 579.885 1541.760 627.650 ;
        RECT 1540.170 579.515 1540.450 579.885 ;
        RECT 1541.550 579.515 1541.830 579.885 ;
        RECT 1540.240 531.410 1540.380 579.515 ;
        RECT 1540.180 531.090 1540.440 531.410 ;
        RECT 1541.100 531.090 1541.360 531.410 ;
        RECT 1541.160 483.325 1541.300 531.090 ;
        RECT 1540.170 482.955 1540.450 483.325 ;
        RECT 1541.090 482.955 1541.370 483.325 ;
        RECT 1540.240 434.850 1540.380 482.955 ;
        RECT 1540.180 434.530 1540.440 434.850 ;
        RECT 1540.180 386.250 1540.440 386.570 ;
        RECT 1540.240 337.950 1540.380 386.250 ;
        RECT 1540.180 337.630 1540.440 337.950 ;
        RECT 1540.180 289.690 1540.440 290.010 ;
        RECT 1540.240 254.730 1540.380 289.690 ;
        RECT 1540.240 254.590 1540.840 254.730 ;
        RECT 1540.700 241.390 1540.840 254.590 ;
        RECT 1540.640 241.070 1540.900 241.390 ;
        RECT 1540.640 193.130 1540.900 193.450 ;
        RECT 1540.700 144.830 1540.840 193.130 ;
        RECT 1540.640 144.510 1540.900 144.830 ;
        RECT 1540.180 96.570 1540.440 96.890 ;
        RECT 1540.240 62.970 1540.380 96.570 ;
        RECT 1539.320 62.830 1540.380 62.970 ;
        RECT 1539.320 50.650 1539.460 62.830 ;
        RECT 772.440 50.330 772.700 50.650 ;
        RECT 1539.260 50.330 1539.520 50.650 ;
        RECT 772.500 16.730 772.640 50.330 ;
        RECT 769.740 16.590 772.640 16.730 ;
        RECT 769.740 2.400 769.880 16.590 ;
        RECT 769.530 -4.800 770.090 2.400 ;
      LAYER via2 ;
        RECT 1540.170 917.520 1540.450 917.800 ;
        RECT 1541.550 917.520 1541.830 917.800 ;
        RECT 1540.170 772.680 1540.450 772.960 ;
        RECT 1541.550 772.680 1541.830 772.960 ;
        RECT 1540.630 676.120 1540.910 676.400 ;
        RECT 1541.550 676.120 1541.830 676.400 ;
        RECT 1540.170 579.560 1540.450 579.840 ;
        RECT 1541.550 579.560 1541.830 579.840 ;
        RECT 1540.170 483.000 1540.450 483.280 ;
        RECT 1541.090 483.000 1541.370 483.280 ;
      LAYER met3 ;
        RECT 1540.145 917.810 1540.475 917.825 ;
        RECT 1541.525 917.810 1541.855 917.825 ;
        RECT 1540.145 917.510 1541.855 917.810 ;
        RECT 1540.145 917.495 1540.475 917.510 ;
        RECT 1541.525 917.495 1541.855 917.510 ;
        RECT 1540.145 772.970 1540.475 772.985 ;
        RECT 1541.525 772.970 1541.855 772.985 ;
        RECT 1540.145 772.670 1541.855 772.970 ;
        RECT 1540.145 772.655 1540.475 772.670 ;
        RECT 1541.525 772.655 1541.855 772.670 ;
        RECT 1540.605 676.410 1540.935 676.425 ;
        RECT 1541.525 676.410 1541.855 676.425 ;
        RECT 1540.605 676.110 1541.855 676.410 ;
        RECT 1540.605 676.095 1540.935 676.110 ;
        RECT 1541.525 676.095 1541.855 676.110 ;
        RECT 1540.145 579.850 1540.475 579.865 ;
        RECT 1541.525 579.850 1541.855 579.865 ;
        RECT 1540.145 579.550 1541.855 579.850 ;
        RECT 1540.145 579.535 1540.475 579.550 ;
        RECT 1541.525 579.535 1541.855 579.550 ;
        RECT 1540.145 483.290 1540.475 483.305 ;
        RECT 1541.065 483.290 1541.395 483.305 ;
        RECT 1540.145 482.990 1541.395 483.290 ;
        RECT 1540.145 482.975 1540.475 482.990 ;
        RECT 1541.065 482.975 1541.395 482.990 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2080.190 1689.700 2080.510 1689.760 ;
        RECT 2214.970 1689.700 2215.290 1689.760 ;
        RECT 2080.190 1689.560 2215.290 1689.700 ;
        RECT 2080.190 1689.500 2080.510 1689.560 ;
        RECT 2214.970 1689.500 2215.290 1689.560 ;
        RECT 2072.370 20.640 2072.690 20.700 ;
        RECT 2080.190 20.640 2080.510 20.700 ;
        RECT 2072.370 20.500 2080.510 20.640 ;
        RECT 2072.370 20.440 2072.690 20.500 ;
        RECT 2080.190 20.440 2080.510 20.500 ;
      LAYER via ;
        RECT 2080.220 1689.500 2080.480 1689.760 ;
        RECT 2215.000 1689.500 2215.260 1689.760 ;
        RECT 2072.400 20.440 2072.660 20.700 ;
        RECT 2080.220 20.440 2080.480 20.700 ;
      LAYER met2 ;
        RECT 2214.920 1700.000 2215.200 1702.400 ;
        RECT 2215.060 1689.790 2215.200 1700.000 ;
        RECT 2080.220 1689.470 2080.480 1689.790 ;
        RECT 2215.000 1689.470 2215.260 1689.790 ;
        RECT 2080.280 20.730 2080.420 1689.470 ;
        RECT 2072.400 20.410 2072.660 20.730 ;
        RECT 2080.220 20.410 2080.480 20.730 ;
        RECT 2072.460 2.400 2072.600 20.410 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2090.845 14.025 2091.015 16.915 ;
        RECT 2138.685 14.025 2138.855 17.255 ;
      LAYER mcon ;
        RECT 2138.685 17.085 2138.855 17.255 ;
        RECT 2090.845 16.745 2091.015 16.915 ;
      LAYER met1 ;
        RECT 2138.625 17.240 2138.915 17.285 ;
        RECT 2138.625 17.100 2215.660 17.240 ;
        RECT 2138.625 17.055 2138.915 17.100 ;
        RECT 2089.850 16.900 2090.170 16.960 ;
        RECT 2090.785 16.900 2091.075 16.945 ;
        RECT 2089.850 16.760 2091.075 16.900 ;
        RECT 2215.520 16.900 2215.660 17.100 ;
        RECT 2222.790 16.900 2223.110 16.960 ;
        RECT 2215.520 16.760 2223.110 16.900 ;
        RECT 2089.850 16.700 2090.170 16.760 ;
        RECT 2090.785 16.715 2091.075 16.760 ;
        RECT 2222.790 16.700 2223.110 16.760 ;
        RECT 2090.785 14.180 2091.075 14.225 ;
        RECT 2138.625 14.180 2138.915 14.225 ;
        RECT 2090.785 14.040 2138.915 14.180 ;
        RECT 2090.785 13.995 2091.075 14.040 ;
        RECT 2138.625 13.995 2138.915 14.040 ;
      LAYER via ;
        RECT 2089.880 16.700 2090.140 16.960 ;
        RECT 2222.820 16.700 2223.080 16.960 ;
      LAYER met2 ;
        RECT 2224.120 1700.410 2224.400 1702.400 ;
        RECT 2222.880 1700.270 2224.400 1700.410 ;
        RECT 2222.880 16.990 2223.020 1700.270 ;
        RECT 2224.120 1700.000 2224.400 1700.270 ;
        RECT 2089.880 16.670 2090.140 16.990 ;
        RECT 2222.820 16.670 2223.080 16.990 ;
        RECT 2089.940 2.400 2090.080 16.670 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2115.225 1686.145 2115.395 1687.335 ;
      LAYER mcon ;
        RECT 2115.225 1687.165 2115.395 1687.335 ;
      LAYER met1 ;
        RECT 2233.370 1687.660 2233.690 1687.720 ;
        RECT 2220.580 1687.520 2233.690 1687.660 ;
        RECT 2115.165 1687.320 2115.455 1687.365 ;
        RECT 2220.580 1687.320 2220.720 1687.520 ;
        RECT 2233.370 1687.460 2233.690 1687.520 ;
        RECT 2115.165 1687.180 2220.720 1687.320 ;
        RECT 2115.165 1687.135 2115.455 1687.180 ;
        RECT 2111.010 1686.300 2111.330 1686.360 ;
        RECT 2115.165 1686.300 2115.455 1686.345 ;
        RECT 2111.010 1686.160 2115.455 1686.300 ;
        RECT 2111.010 1686.100 2111.330 1686.160 ;
        RECT 2115.165 1686.115 2115.455 1686.160 ;
        RECT 2107.790 14.520 2108.110 14.580 ;
        RECT 2111.010 14.520 2111.330 14.580 ;
        RECT 2107.790 14.380 2111.330 14.520 ;
        RECT 2107.790 14.320 2108.110 14.380 ;
        RECT 2111.010 14.320 2111.330 14.380 ;
      LAYER via ;
        RECT 2233.400 1687.460 2233.660 1687.720 ;
        RECT 2111.040 1686.100 2111.300 1686.360 ;
        RECT 2107.820 14.320 2108.080 14.580 ;
        RECT 2111.040 14.320 2111.300 14.580 ;
      LAYER met2 ;
        RECT 2233.320 1700.000 2233.600 1702.400 ;
        RECT 2233.460 1687.750 2233.600 1700.000 ;
        RECT 2233.400 1687.430 2233.660 1687.750 ;
        RECT 2111.040 1686.070 2111.300 1686.390 ;
        RECT 2111.100 14.610 2111.240 1686.070 ;
        RECT 2107.820 14.290 2108.080 14.610 ;
        RECT 2111.040 14.290 2111.300 14.610 ;
        RECT 2107.880 2.400 2108.020 14.290 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2242.570 19.960 2242.890 20.020 ;
        RECT 2163.540 19.820 2242.890 19.960 ;
        RECT 2125.730 19.620 2126.050 19.680 ;
        RECT 2163.540 19.620 2163.680 19.820 ;
        RECT 2242.570 19.760 2242.890 19.820 ;
        RECT 2125.730 19.480 2163.680 19.620 ;
        RECT 2125.730 19.420 2126.050 19.480 ;
      LAYER via ;
        RECT 2125.760 19.420 2126.020 19.680 ;
        RECT 2242.600 19.760 2242.860 20.020 ;
      LAYER met2 ;
        RECT 2242.520 1700.000 2242.800 1702.400 ;
        RECT 2242.660 20.050 2242.800 1700.000 ;
        RECT 2242.600 19.730 2242.860 20.050 ;
        RECT 2125.760 19.390 2126.020 19.710 ;
        RECT 2125.820 2.400 2125.960 19.390 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2167.205 1686.485 2167.375 1687.675 ;
        RECT 2210.905 1686.485 2211.075 1689.375 ;
      LAYER mcon ;
        RECT 2210.905 1689.205 2211.075 1689.375 ;
        RECT 2167.205 1687.505 2167.375 1687.675 ;
      LAYER met1 ;
        RECT 2251.770 1690.040 2252.090 1690.100 ;
        RECT 2218.740 1689.900 2252.090 1690.040 ;
        RECT 2210.845 1689.360 2211.135 1689.405 ;
        RECT 2218.740 1689.360 2218.880 1689.900 ;
        RECT 2251.770 1689.840 2252.090 1689.900 ;
        RECT 2210.845 1689.220 2218.880 1689.360 ;
        RECT 2210.845 1689.175 2211.135 1689.220 ;
        RECT 2145.510 1687.660 2145.830 1687.720 ;
        RECT 2167.145 1687.660 2167.435 1687.705 ;
        RECT 2145.510 1687.520 2167.435 1687.660 ;
        RECT 2145.510 1687.460 2145.830 1687.520 ;
        RECT 2167.145 1687.475 2167.435 1687.520 ;
        RECT 2167.145 1686.640 2167.435 1686.685 ;
        RECT 2210.845 1686.640 2211.135 1686.685 ;
        RECT 2167.145 1686.500 2211.135 1686.640 ;
        RECT 2167.145 1686.455 2167.435 1686.500 ;
        RECT 2210.845 1686.455 2211.135 1686.500 ;
      LAYER via ;
        RECT 2251.800 1689.840 2252.060 1690.100 ;
        RECT 2145.540 1687.460 2145.800 1687.720 ;
      LAYER met2 ;
        RECT 2251.720 1700.000 2252.000 1702.400 ;
        RECT 2251.860 1690.130 2252.000 1700.000 ;
        RECT 2251.800 1689.810 2252.060 1690.130 ;
        RECT 2145.540 1687.430 2145.800 1687.750 ;
        RECT 2145.600 3.130 2145.740 1687.430 ;
        RECT 2143.760 2.990 2145.740 3.130 ;
        RECT 2143.760 2.400 2143.900 2.990 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2257.365 1652.485 2257.535 1690.395 ;
        RECT 2257.825 1510.365 2257.995 1579.895 ;
        RECT 2257.825 1317.245 2257.995 1368.755 ;
        RECT 2257.825 1220.685 2257.995 1297.015 ;
        RECT 2258.285 869.465 2258.455 917.575 ;
        RECT 2258.285 737.885 2258.455 772.735 ;
        RECT 2257.365 572.645 2257.535 620.755 ;
        RECT 2257.825 476.085 2257.995 524.195 ;
        RECT 2257.365 338.045 2257.535 427.635 ;
        RECT 2257.365 303.365 2257.535 331.075 ;
        RECT 2258.285 234.685 2258.455 282.795 ;
        RECT 2258.745 96.645 2258.915 144.755 ;
      LAYER mcon ;
        RECT 2257.365 1690.225 2257.535 1690.395 ;
        RECT 2257.825 1579.725 2257.995 1579.895 ;
        RECT 2257.825 1368.585 2257.995 1368.755 ;
        RECT 2257.825 1296.845 2257.995 1297.015 ;
        RECT 2258.285 917.405 2258.455 917.575 ;
        RECT 2258.285 772.565 2258.455 772.735 ;
        RECT 2257.365 620.585 2257.535 620.755 ;
        RECT 2257.825 524.025 2257.995 524.195 ;
        RECT 2257.365 427.465 2257.535 427.635 ;
        RECT 2257.365 330.905 2257.535 331.075 ;
        RECT 2258.285 282.625 2258.455 282.795 ;
        RECT 2258.745 144.585 2258.915 144.755 ;
      LAYER met1 ;
        RECT 2257.305 1690.380 2257.595 1690.425 ;
        RECT 2258.670 1690.380 2258.990 1690.440 ;
        RECT 2257.305 1690.240 2258.990 1690.380 ;
        RECT 2257.305 1690.195 2257.595 1690.240 ;
        RECT 2258.670 1690.180 2258.990 1690.240 ;
        RECT 2257.305 1652.640 2257.595 1652.685 ;
        RECT 2257.750 1652.640 2258.070 1652.700 ;
        RECT 2257.305 1652.500 2258.070 1652.640 ;
        RECT 2257.305 1652.455 2257.595 1652.500 ;
        RECT 2257.750 1652.440 2258.070 1652.500 ;
        RECT 2257.750 1580.560 2258.070 1580.620 ;
        RECT 2258.670 1580.560 2258.990 1580.620 ;
        RECT 2257.750 1580.420 2258.990 1580.560 ;
        RECT 2257.750 1580.360 2258.070 1580.420 ;
        RECT 2258.670 1580.360 2258.990 1580.420 ;
        RECT 2257.750 1579.880 2258.070 1579.940 ;
        RECT 2257.555 1579.740 2258.070 1579.880 ;
        RECT 2257.750 1579.680 2258.070 1579.740 ;
        RECT 2257.750 1510.520 2258.070 1510.580 ;
        RECT 2257.555 1510.380 2258.070 1510.520 ;
        RECT 2257.750 1510.320 2258.070 1510.380 ;
        RECT 2257.750 1463.260 2258.070 1463.320 ;
        RECT 2257.380 1463.120 2258.070 1463.260 ;
        RECT 2257.380 1462.640 2257.520 1463.120 ;
        RECT 2257.750 1463.060 2258.070 1463.120 ;
        RECT 2257.290 1462.380 2257.610 1462.640 ;
        RECT 2256.370 1393.900 2256.690 1393.960 ;
        RECT 2257.750 1393.900 2258.070 1393.960 ;
        RECT 2256.370 1393.760 2258.070 1393.900 ;
        RECT 2256.370 1393.700 2256.690 1393.760 ;
        RECT 2257.750 1393.700 2258.070 1393.760 ;
        RECT 2257.750 1368.740 2258.070 1368.800 ;
        RECT 2257.555 1368.600 2258.070 1368.740 ;
        RECT 2257.750 1368.540 2258.070 1368.600 ;
        RECT 2257.750 1317.400 2258.070 1317.460 ;
        RECT 2257.555 1317.260 2258.070 1317.400 ;
        RECT 2257.750 1317.200 2258.070 1317.260 ;
        RECT 2257.750 1297.000 2258.070 1297.060 ;
        RECT 2257.555 1296.860 2258.070 1297.000 ;
        RECT 2257.750 1296.800 2258.070 1296.860 ;
        RECT 2257.750 1220.840 2258.070 1220.900 ;
        RECT 2257.555 1220.700 2258.070 1220.840 ;
        RECT 2257.750 1220.640 2258.070 1220.700 ;
        RECT 2257.750 1173.580 2258.070 1173.640 ;
        RECT 2257.380 1173.440 2258.070 1173.580 ;
        RECT 2257.380 1172.960 2257.520 1173.440 ;
        RECT 2257.750 1173.380 2258.070 1173.440 ;
        RECT 2257.290 1172.700 2257.610 1172.960 ;
        RECT 2256.370 1111.020 2256.690 1111.080 ;
        RECT 2257.750 1111.020 2258.070 1111.080 ;
        RECT 2256.370 1110.880 2258.070 1111.020 ;
        RECT 2256.370 1110.820 2256.690 1110.880 ;
        RECT 2257.750 1110.820 2258.070 1110.880 ;
        RECT 2257.750 1077.020 2258.070 1077.080 ;
        RECT 2257.380 1076.880 2258.070 1077.020 ;
        RECT 2257.380 1076.400 2257.520 1076.880 ;
        RECT 2257.750 1076.820 2258.070 1076.880 ;
        RECT 2257.290 1076.140 2257.610 1076.400 ;
        RECT 2256.370 1014.460 2256.690 1014.520 ;
        RECT 2257.750 1014.460 2258.070 1014.520 ;
        RECT 2256.370 1014.320 2258.070 1014.460 ;
        RECT 2256.370 1014.260 2256.690 1014.320 ;
        RECT 2257.750 1014.260 2258.070 1014.320 ;
        RECT 2257.750 980.460 2258.070 980.520 ;
        RECT 2257.380 980.320 2258.070 980.460 ;
        RECT 2257.380 979.840 2257.520 980.320 ;
        RECT 2257.750 980.260 2258.070 980.320 ;
        RECT 2257.290 979.580 2257.610 979.840 ;
        RECT 2257.290 931.500 2257.610 931.560 ;
        RECT 2258.210 931.500 2258.530 931.560 ;
        RECT 2257.290 931.360 2258.530 931.500 ;
        RECT 2257.290 931.300 2257.610 931.360 ;
        RECT 2258.210 931.300 2258.530 931.360 ;
        RECT 2258.210 917.560 2258.530 917.620 ;
        RECT 2258.015 917.420 2258.530 917.560 ;
        RECT 2258.210 917.360 2258.530 917.420 ;
        RECT 2258.225 869.620 2258.515 869.665 ;
        RECT 2258.670 869.620 2258.990 869.680 ;
        RECT 2258.225 869.480 2258.990 869.620 ;
        RECT 2258.225 869.435 2258.515 869.480 ;
        RECT 2258.670 869.420 2258.990 869.480 ;
        RECT 2258.210 786.460 2258.530 786.720 ;
        RECT 2258.300 786.040 2258.440 786.460 ;
        RECT 2258.210 785.780 2258.530 786.040 ;
        RECT 2258.210 772.720 2258.530 772.780 ;
        RECT 2258.015 772.580 2258.530 772.720 ;
        RECT 2258.210 772.520 2258.530 772.580 ;
        RECT 2258.210 738.040 2258.530 738.100 ;
        RECT 2258.015 737.900 2258.530 738.040 ;
        RECT 2258.210 737.840 2258.530 737.900 ;
        RECT 2258.210 676.500 2258.530 676.560 ;
        RECT 2258.670 676.500 2258.990 676.560 ;
        RECT 2258.210 676.360 2258.990 676.500 ;
        RECT 2258.210 676.300 2258.530 676.360 ;
        RECT 2258.670 676.300 2258.990 676.360 ;
        RECT 2257.290 620.740 2257.610 620.800 ;
        RECT 2257.095 620.600 2257.610 620.740 ;
        RECT 2257.290 620.540 2257.610 620.600 ;
        RECT 2257.305 572.800 2257.595 572.845 ;
        RECT 2257.750 572.800 2258.070 572.860 ;
        RECT 2257.305 572.660 2258.070 572.800 ;
        RECT 2257.305 572.615 2257.595 572.660 ;
        RECT 2257.750 572.600 2258.070 572.660 ;
        RECT 2257.750 524.180 2258.070 524.240 ;
        RECT 2257.555 524.040 2258.070 524.180 ;
        RECT 2257.750 523.980 2258.070 524.040 ;
        RECT 2257.750 476.240 2258.070 476.300 ;
        RECT 2257.555 476.100 2258.070 476.240 ;
        RECT 2257.750 476.040 2258.070 476.100 ;
        RECT 2257.305 427.620 2257.595 427.665 ;
        RECT 2257.750 427.620 2258.070 427.680 ;
        RECT 2257.305 427.480 2258.070 427.620 ;
        RECT 2257.305 427.435 2257.595 427.480 ;
        RECT 2257.750 427.420 2258.070 427.480 ;
        RECT 2257.290 338.200 2257.610 338.260 ;
        RECT 2257.095 338.060 2257.610 338.200 ;
        RECT 2257.290 338.000 2257.610 338.060 ;
        RECT 2257.290 331.060 2257.610 331.120 ;
        RECT 2257.095 330.920 2257.610 331.060 ;
        RECT 2257.290 330.860 2257.610 330.920 ;
        RECT 2257.305 303.520 2257.595 303.565 ;
        RECT 2258.210 303.520 2258.530 303.580 ;
        RECT 2257.305 303.380 2258.530 303.520 ;
        RECT 2257.305 303.335 2257.595 303.380 ;
        RECT 2258.210 303.320 2258.530 303.380 ;
        RECT 2258.210 282.780 2258.530 282.840 ;
        RECT 2258.015 282.640 2258.530 282.780 ;
        RECT 2258.210 282.580 2258.530 282.640 ;
        RECT 2258.225 234.840 2258.515 234.885 ;
        RECT 2259.130 234.840 2259.450 234.900 ;
        RECT 2258.225 234.700 2259.450 234.840 ;
        RECT 2258.225 234.655 2258.515 234.700 ;
        RECT 2259.130 234.640 2259.450 234.700 ;
        RECT 2258.210 158.680 2258.530 158.740 ;
        RECT 2259.130 158.680 2259.450 158.740 ;
        RECT 2258.210 158.540 2259.450 158.680 ;
        RECT 2258.210 158.480 2258.530 158.540 ;
        RECT 2259.130 158.480 2259.450 158.540 ;
        RECT 2258.685 144.740 2258.975 144.785 ;
        RECT 2259.130 144.740 2259.450 144.800 ;
        RECT 2258.685 144.600 2259.450 144.740 ;
        RECT 2258.685 144.555 2258.975 144.600 ;
        RECT 2259.130 144.540 2259.450 144.600 ;
        RECT 2258.670 96.800 2258.990 96.860 ;
        RECT 2258.475 96.660 2258.990 96.800 ;
        RECT 2258.670 96.600 2258.990 96.660 ;
        RECT 2161.610 17.580 2161.930 17.640 ;
        RECT 2257.750 17.580 2258.070 17.640 ;
        RECT 2161.610 17.440 2258.070 17.580 ;
        RECT 2161.610 17.380 2161.930 17.440 ;
        RECT 2257.750 17.380 2258.070 17.440 ;
      LAYER via ;
        RECT 2258.700 1690.180 2258.960 1690.440 ;
        RECT 2257.780 1652.440 2258.040 1652.700 ;
        RECT 2257.780 1580.360 2258.040 1580.620 ;
        RECT 2258.700 1580.360 2258.960 1580.620 ;
        RECT 2257.780 1579.680 2258.040 1579.940 ;
        RECT 2257.780 1510.320 2258.040 1510.580 ;
        RECT 2257.780 1463.060 2258.040 1463.320 ;
        RECT 2257.320 1462.380 2257.580 1462.640 ;
        RECT 2256.400 1393.700 2256.660 1393.960 ;
        RECT 2257.780 1393.700 2258.040 1393.960 ;
        RECT 2257.780 1368.540 2258.040 1368.800 ;
        RECT 2257.780 1317.200 2258.040 1317.460 ;
        RECT 2257.780 1296.800 2258.040 1297.060 ;
        RECT 2257.780 1220.640 2258.040 1220.900 ;
        RECT 2257.780 1173.380 2258.040 1173.640 ;
        RECT 2257.320 1172.700 2257.580 1172.960 ;
        RECT 2256.400 1110.820 2256.660 1111.080 ;
        RECT 2257.780 1110.820 2258.040 1111.080 ;
        RECT 2257.780 1076.820 2258.040 1077.080 ;
        RECT 2257.320 1076.140 2257.580 1076.400 ;
        RECT 2256.400 1014.260 2256.660 1014.520 ;
        RECT 2257.780 1014.260 2258.040 1014.520 ;
        RECT 2257.780 980.260 2258.040 980.520 ;
        RECT 2257.320 979.580 2257.580 979.840 ;
        RECT 2257.320 931.300 2257.580 931.560 ;
        RECT 2258.240 931.300 2258.500 931.560 ;
        RECT 2258.240 917.360 2258.500 917.620 ;
        RECT 2258.700 869.420 2258.960 869.680 ;
        RECT 2258.240 786.460 2258.500 786.720 ;
        RECT 2258.240 785.780 2258.500 786.040 ;
        RECT 2258.240 772.520 2258.500 772.780 ;
        RECT 2258.240 737.840 2258.500 738.100 ;
        RECT 2258.240 676.300 2258.500 676.560 ;
        RECT 2258.700 676.300 2258.960 676.560 ;
        RECT 2257.320 620.540 2257.580 620.800 ;
        RECT 2257.780 572.600 2258.040 572.860 ;
        RECT 2257.780 523.980 2258.040 524.240 ;
        RECT 2257.780 476.040 2258.040 476.300 ;
        RECT 2257.780 427.420 2258.040 427.680 ;
        RECT 2257.320 338.000 2257.580 338.260 ;
        RECT 2257.320 330.860 2257.580 331.120 ;
        RECT 2258.240 303.320 2258.500 303.580 ;
        RECT 2258.240 282.580 2258.500 282.840 ;
        RECT 2259.160 234.640 2259.420 234.900 ;
        RECT 2258.240 158.480 2258.500 158.740 ;
        RECT 2259.160 158.480 2259.420 158.740 ;
        RECT 2259.160 144.540 2259.420 144.800 ;
        RECT 2258.700 96.600 2258.960 96.860 ;
        RECT 2161.640 17.380 2161.900 17.640 ;
        RECT 2257.780 17.380 2258.040 17.640 ;
      LAYER met2 ;
        RECT 2260.920 1701.090 2261.200 1702.400 ;
        RECT 2258.760 1700.950 2261.200 1701.090 ;
        RECT 2258.760 1690.470 2258.900 1700.950 ;
        RECT 2260.920 1700.000 2261.200 1700.950 ;
        RECT 2258.700 1690.150 2258.960 1690.470 ;
        RECT 2257.780 1652.410 2258.040 1652.730 ;
        RECT 2257.840 1628.445 2257.980 1652.410 ;
        RECT 2257.770 1628.075 2258.050 1628.445 ;
        RECT 2258.690 1628.075 2258.970 1628.445 ;
        RECT 2258.760 1580.650 2258.900 1628.075 ;
        RECT 2257.780 1580.330 2258.040 1580.650 ;
        RECT 2258.700 1580.330 2258.960 1580.650 ;
        RECT 2257.840 1579.970 2257.980 1580.330 ;
        RECT 2257.780 1579.650 2258.040 1579.970 ;
        RECT 2257.780 1510.290 2258.040 1510.610 ;
        RECT 2257.840 1463.350 2257.980 1510.290 ;
        RECT 2257.780 1463.030 2258.040 1463.350 ;
        RECT 2257.320 1462.350 2257.580 1462.670 ;
        RECT 2257.380 1442.125 2257.520 1462.350 ;
        RECT 2256.390 1441.755 2256.670 1442.125 ;
        RECT 2257.310 1441.755 2257.590 1442.125 ;
        RECT 2256.460 1393.990 2256.600 1441.755 ;
        RECT 2256.400 1393.670 2256.660 1393.990 ;
        RECT 2257.780 1393.670 2258.040 1393.990 ;
        RECT 2257.840 1368.830 2257.980 1393.670 ;
        RECT 2257.780 1368.510 2258.040 1368.830 ;
        RECT 2257.780 1317.170 2258.040 1317.490 ;
        RECT 2257.840 1297.090 2257.980 1317.170 ;
        RECT 2257.780 1296.770 2258.040 1297.090 ;
        RECT 2257.780 1220.610 2258.040 1220.930 ;
        RECT 2257.840 1173.670 2257.980 1220.610 ;
        RECT 2257.780 1173.350 2258.040 1173.670 ;
        RECT 2257.320 1172.670 2257.580 1172.990 ;
        RECT 2257.380 1159.245 2257.520 1172.670 ;
        RECT 2256.390 1158.875 2256.670 1159.245 ;
        RECT 2257.310 1158.875 2257.590 1159.245 ;
        RECT 2256.460 1111.110 2256.600 1158.875 ;
        RECT 2256.400 1110.790 2256.660 1111.110 ;
        RECT 2257.780 1110.790 2258.040 1111.110 ;
        RECT 2257.840 1077.110 2257.980 1110.790 ;
        RECT 2257.780 1076.790 2258.040 1077.110 ;
        RECT 2257.320 1076.110 2257.580 1076.430 ;
        RECT 2257.380 1062.685 2257.520 1076.110 ;
        RECT 2256.390 1062.315 2256.670 1062.685 ;
        RECT 2257.310 1062.315 2257.590 1062.685 ;
        RECT 2256.460 1014.550 2256.600 1062.315 ;
        RECT 2256.400 1014.230 2256.660 1014.550 ;
        RECT 2257.780 1014.230 2258.040 1014.550 ;
        RECT 2257.840 980.550 2257.980 1014.230 ;
        RECT 2257.780 980.230 2258.040 980.550 ;
        RECT 2257.320 979.550 2257.580 979.870 ;
        RECT 2257.380 931.590 2257.520 979.550 ;
        RECT 2257.320 931.270 2257.580 931.590 ;
        RECT 2258.240 931.270 2258.500 931.590 ;
        RECT 2258.300 917.650 2258.440 931.270 ;
        RECT 2258.240 917.330 2258.500 917.650 ;
        RECT 2258.700 869.390 2258.960 869.710 ;
        RECT 2258.760 834.770 2258.900 869.390 ;
        RECT 2258.300 834.630 2258.900 834.770 ;
        RECT 2258.300 786.750 2258.440 834.630 ;
        RECT 2258.240 786.430 2258.500 786.750 ;
        RECT 2258.240 785.750 2258.500 786.070 ;
        RECT 2258.300 772.810 2258.440 785.750 ;
        RECT 2258.240 772.490 2258.500 772.810 ;
        RECT 2258.240 737.810 2258.500 738.130 ;
        RECT 2258.300 724.610 2258.440 737.810 ;
        RECT 2258.300 724.470 2258.900 724.610 ;
        RECT 2258.760 676.590 2258.900 724.470 ;
        RECT 2258.240 676.330 2258.500 676.590 ;
        RECT 2257.840 676.270 2258.500 676.330 ;
        RECT 2258.700 676.270 2258.960 676.590 ;
        RECT 2257.840 676.190 2258.440 676.270 ;
        RECT 2257.840 642.330 2257.980 676.190 ;
        RECT 2257.840 642.190 2258.440 642.330 ;
        RECT 2258.300 640.970 2258.440 642.190 ;
        RECT 2257.380 640.830 2258.440 640.970 ;
        RECT 2257.380 620.830 2257.520 640.830 ;
        RECT 2257.320 620.510 2257.580 620.830 ;
        RECT 2257.780 572.570 2258.040 572.890 ;
        RECT 2257.840 524.270 2257.980 572.570 ;
        RECT 2257.780 523.950 2258.040 524.270 ;
        RECT 2257.780 476.010 2258.040 476.330 ;
        RECT 2257.840 427.710 2257.980 476.010 ;
        RECT 2257.780 427.390 2258.040 427.710 ;
        RECT 2257.320 337.970 2257.580 338.290 ;
        RECT 2257.380 331.150 2257.520 337.970 ;
        RECT 2257.320 330.830 2257.580 331.150 ;
        RECT 2258.240 303.290 2258.500 303.610 ;
        RECT 2258.300 282.870 2258.440 303.290 ;
        RECT 2258.240 282.550 2258.500 282.870 ;
        RECT 2259.160 234.610 2259.420 234.930 ;
        RECT 2259.220 234.330 2259.360 234.610 ;
        RECT 2258.300 234.190 2259.360 234.330 ;
        RECT 2258.300 158.770 2258.440 234.190 ;
        RECT 2258.240 158.450 2258.500 158.770 ;
        RECT 2259.160 158.450 2259.420 158.770 ;
        RECT 2259.220 144.830 2259.360 158.450 ;
        RECT 2259.160 144.510 2259.420 144.830 ;
        RECT 2258.700 96.570 2258.960 96.890 ;
        RECT 2258.760 62.290 2258.900 96.570 ;
        RECT 2257.840 62.150 2258.900 62.290 ;
        RECT 2257.840 17.670 2257.980 62.150 ;
        RECT 2161.640 17.350 2161.900 17.670 ;
        RECT 2257.780 17.350 2258.040 17.670 ;
        RECT 2161.700 2.400 2161.840 17.350 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
      LAYER via2 ;
        RECT 2257.770 1628.120 2258.050 1628.400 ;
        RECT 2258.690 1628.120 2258.970 1628.400 ;
        RECT 2256.390 1441.800 2256.670 1442.080 ;
        RECT 2257.310 1441.800 2257.590 1442.080 ;
        RECT 2256.390 1158.920 2256.670 1159.200 ;
        RECT 2257.310 1158.920 2257.590 1159.200 ;
        RECT 2256.390 1062.360 2256.670 1062.640 ;
        RECT 2257.310 1062.360 2257.590 1062.640 ;
      LAYER met3 ;
        RECT 2257.745 1628.410 2258.075 1628.425 ;
        RECT 2258.665 1628.410 2258.995 1628.425 ;
        RECT 2257.745 1628.110 2258.995 1628.410 ;
        RECT 2257.745 1628.095 2258.075 1628.110 ;
        RECT 2258.665 1628.095 2258.995 1628.110 ;
        RECT 2256.365 1442.090 2256.695 1442.105 ;
        RECT 2257.285 1442.090 2257.615 1442.105 ;
        RECT 2256.365 1441.790 2257.615 1442.090 ;
        RECT 2256.365 1441.775 2256.695 1441.790 ;
        RECT 2257.285 1441.775 2257.615 1441.790 ;
        RECT 2256.365 1159.210 2256.695 1159.225 ;
        RECT 2257.285 1159.210 2257.615 1159.225 ;
        RECT 2256.365 1158.910 2257.615 1159.210 ;
        RECT 2256.365 1158.895 2256.695 1158.910 ;
        RECT 2257.285 1158.895 2257.615 1158.910 ;
        RECT 2256.365 1062.650 2256.695 1062.665 ;
        RECT 2257.285 1062.650 2257.615 1062.665 ;
        RECT 2256.365 1062.350 2257.615 1062.650 ;
        RECT 2256.365 1062.335 2256.695 1062.350 ;
        RECT 2257.285 1062.335 2257.615 1062.350 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.010 1685.280 2180.330 1685.340 ;
        RECT 2270.170 1685.280 2270.490 1685.340 ;
        RECT 2180.010 1685.140 2270.490 1685.280 ;
        RECT 2180.010 1685.080 2180.330 1685.140 ;
        RECT 2270.170 1685.080 2270.490 1685.140 ;
        RECT 2179.090 2.960 2179.410 3.020 ;
        RECT 2180.010 2.960 2180.330 3.020 ;
        RECT 2179.090 2.820 2180.330 2.960 ;
        RECT 2179.090 2.760 2179.410 2.820 ;
        RECT 2180.010 2.760 2180.330 2.820 ;
      LAYER via ;
        RECT 2180.040 1685.080 2180.300 1685.340 ;
        RECT 2270.200 1685.080 2270.460 1685.340 ;
        RECT 2179.120 2.760 2179.380 3.020 ;
        RECT 2180.040 2.760 2180.300 3.020 ;
      LAYER met2 ;
        RECT 2270.120 1700.000 2270.400 1702.400 ;
        RECT 2270.260 1685.370 2270.400 1700.000 ;
        RECT 2180.040 1685.050 2180.300 1685.370 ;
        RECT 2270.200 1685.050 2270.460 1685.370 ;
        RECT 2180.100 3.050 2180.240 1685.050 ;
        RECT 2179.120 2.730 2179.380 3.050 ;
        RECT 2180.040 2.730 2180.300 3.050 ;
        RECT 2179.180 2.400 2179.320 2.730 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2238.505 17.765 2238.675 18.615 ;
      LAYER mcon ;
        RECT 2238.505 18.445 2238.675 18.615 ;
      LAYER met1 ;
        RECT 2277.990 18.940 2278.310 19.000 ;
        RECT 2239.440 18.800 2278.310 18.940 ;
        RECT 2238.445 18.600 2238.735 18.645 ;
        RECT 2239.440 18.600 2239.580 18.800 ;
        RECT 2277.990 18.740 2278.310 18.800 ;
        RECT 2238.445 18.460 2239.580 18.600 ;
        RECT 2238.445 18.415 2238.735 18.460 ;
        RECT 2197.030 17.920 2197.350 17.980 ;
        RECT 2238.445 17.920 2238.735 17.965 ;
        RECT 2197.030 17.780 2238.735 17.920 ;
        RECT 2197.030 17.720 2197.350 17.780 ;
        RECT 2238.445 17.735 2238.735 17.780 ;
      LAYER via ;
        RECT 2278.020 18.740 2278.280 19.000 ;
        RECT 2197.060 17.720 2197.320 17.980 ;
      LAYER met2 ;
        RECT 2279.320 1700.410 2279.600 1702.400 ;
        RECT 2278.080 1700.270 2279.600 1700.410 ;
        RECT 2278.080 19.030 2278.220 1700.270 ;
        RECT 2279.320 1700.000 2279.600 1700.270 ;
        RECT 2278.020 18.710 2278.280 19.030 ;
        RECT 2197.060 17.690 2197.320 18.010 ;
        RECT 2197.120 2.400 2197.260 17.690 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2214.970 18.260 2215.290 18.320 ;
        RECT 2284.430 18.260 2284.750 18.320 ;
        RECT 2214.970 18.120 2284.750 18.260 ;
        RECT 2214.970 18.060 2215.290 18.120 ;
        RECT 2284.430 18.060 2284.750 18.120 ;
      LAYER via ;
        RECT 2215.000 18.060 2215.260 18.320 ;
        RECT 2284.460 18.060 2284.720 18.320 ;
      LAYER met2 ;
        RECT 2288.520 1701.090 2288.800 1702.400 ;
        RECT 2286.360 1700.950 2288.800 1701.090 ;
        RECT 2286.360 1656.210 2286.500 1700.950 ;
        RECT 2288.520 1700.000 2288.800 1700.950 ;
        RECT 2284.520 1656.070 2286.500 1656.210 ;
        RECT 2284.520 18.350 2284.660 1656.070 ;
        RECT 2215.000 18.030 2215.260 18.350 ;
        RECT 2284.460 18.030 2284.720 18.350 ;
        RECT 2215.060 2.400 2215.200 18.030 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2298.690 17.580 2299.010 17.640 ;
        RECT 2259.680 17.440 2299.010 17.580 ;
        RECT 2232.910 17.240 2233.230 17.300 ;
        RECT 2259.680 17.240 2259.820 17.440 ;
        RECT 2298.690 17.380 2299.010 17.440 ;
        RECT 2232.910 17.100 2259.820 17.240 ;
        RECT 2232.910 17.040 2233.230 17.100 ;
      LAYER via ;
        RECT 2232.940 17.040 2233.200 17.300 ;
        RECT 2298.720 17.380 2298.980 17.640 ;
      LAYER met2 ;
        RECT 2297.720 1700.410 2298.000 1702.400 ;
        RECT 2297.720 1700.270 2298.920 1700.410 ;
        RECT 2297.720 1700.000 2298.000 1700.270 ;
        RECT 2298.780 17.670 2298.920 1700.270 ;
        RECT 2298.720 17.350 2298.980 17.670 ;
        RECT 2232.940 17.010 2233.200 17.330 ;
        RECT 2233.000 2.400 2233.140 17.010 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 50.220 793.430 50.280 ;
        RECT 1552.570 50.220 1552.890 50.280 ;
        RECT 793.110 50.080 1552.890 50.220 ;
        RECT 793.110 50.020 793.430 50.080 ;
        RECT 1552.570 50.020 1552.890 50.080 ;
      LAYER via ;
        RECT 793.140 50.020 793.400 50.280 ;
        RECT 1552.600 50.020 1552.860 50.280 ;
      LAYER met2 ;
        RECT 1553.900 1700.410 1554.180 1702.400 ;
        RECT 1552.660 1700.270 1554.180 1700.410 ;
        RECT 1552.660 50.310 1552.800 1700.270 ;
        RECT 1553.900 1700.000 1554.180 1700.270 ;
        RECT 793.140 49.990 793.400 50.310 ;
        RECT 1552.600 49.990 1552.860 50.310 ;
        RECT 793.200 16.730 793.340 49.990 ;
        RECT 787.680 16.590 793.340 16.730 ;
        RECT 787.680 2.400 787.820 16.590 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2255.910 1687.660 2256.230 1687.720 ;
        RECT 2306.970 1687.660 2307.290 1687.720 ;
        RECT 2255.910 1687.520 2307.290 1687.660 ;
        RECT 2255.910 1687.460 2256.230 1687.520 ;
        RECT 2306.970 1687.460 2307.290 1687.520 ;
        RECT 2250.850 18.600 2251.170 18.660 ;
        RECT 2255.910 18.600 2256.230 18.660 ;
        RECT 2250.850 18.460 2256.230 18.600 ;
        RECT 2250.850 18.400 2251.170 18.460 ;
        RECT 2255.910 18.400 2256.230 18.460 ;
      LAYER via ;
        RECT 2255.940 1687.460 2256.200 1687.720 ;
        RECT 2307.000 1687.460 2307.260 1687.720 ;
        RECT 2250.880 18.400 2251.140 18.660 ;
        RECT 2255.940 18.400 2256.200 18.660 ;
      LAYER met2 ;
        RECT 2306.920 1700.000 2307.200 1702.400 ;
        RECT 2307.060 1687.750 2307.200 1700.000 ;
        RECT 2255.940 1687.430 2256.200 1687.750 ;
        RECT 2307.000 1687.430 2307.260 1687.750 ;
        RECT 2256.000 18.690 2256.140 1687.430 ;
        RECT 2250.880 18.370 2251.140 18.690 ;
        RECT 2255.940 18.370 2256.200 18.690 ;
        RECT 2250.940 2.400 2251.080 18.370 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.710 1688.000 2270.030 1688.060 ;
        RECT 2316.170 1688.000 2316.490 1688.060 ;
        RECT 2269.710 1687.860 2316.490 1688.000 ;
        RECT 2269.710 1687.800 2270.030 1687.860 ;
        RECT 2316.170 1687.800 2316.490 1687.860 ;
        RECT 2268.330 2.960 2268.650 3.020 ;
        RECT 2269.710 2.960 2270.030 3.020 ;
        RECT 2268.330 2.820 2270.030 2.960 ;
        RECT 2268.330 2.760 2268.650 2.820 ;
        RECT 2269.710 2.760 2270.030 2.820 ;
      LAYER via ;
        RECT 2269.740 1687.800 2270.000 1688.060 ;
        RECT 2316.200 1687.800 2316.460 1688.060 ;
        RECT 2268.360 2.760 2268.620 3.020 ;
        RECT 2269.740 2.760 2270.000 3.020 ;
      LAYER met2 ;
        RECT 2316.120 1700.000 2316.400 1702.400 ;
        RECT 2316.260 1688.090 2316.400 1700.000 ;
        RECT 2269.740 1687.770 2270.000 1688.090 ;
        RECT 2316.200 1687.770 2316.460 1688.090 ;
        RECT 2269.800 3.050 2269.940 1687.770 ;
        RECT 2268.360 2.730 2268.620 3.050 ;
        RECT 2269.740 2.730 2270.000 3.050 ;
        RECT 2268.420 2.400 2268.560 2.730 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2286.270 18.600 2286.590 18.660 ;
        RECT 2326.750 18.600 2327.070 18.660 ;
        RECT 2286.270 18.460 2327.070 18.600 ;
        RECT 2286.270 18.400 2286.590 18.460 ;
        RECT 2326.750 18.400 2327.070 18.460 ;
      LAYER via ;
        RECT 2286.300 18.400 2286.560 18.660 ;
        RECT 2326.780 18.400 2327.040 18.660 ;
      LAYER met2 ;
        RECT 2325.320 1700.410 2325.600 1702.400 ;
        RECT 2325.320 1700.270 2326.980 1700.410 ;
        RECT 2325.320 1700.000 2325.600 1700.270 ;
        RECT 2326.840 18.690 2326.980 1700.270 ;
        RECT 2286.300 18.370 2286.560 18.690 ;
        RECT 2326.780 18.370 2327.040 18.690 ;
        RECT 2286.360 2.400 2286.500 18.370 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2304.210 1686.980 2304.530 1687.040 ;
        RECT 2334.570 1686.980 2334.890 1687.040 ;
        RECT 2304.210 1686.840 2334.890 1686.980 ;
        RECT 2304.210 1686.780 2304.530 1686.840 ;
        RECT 2334.570 1686.780 2334.890 1686.840 ;
      LAYER via ;
        RECT 2304.240 1686.780 2304.500 1687.040 ;
        RECT 2334.600 1686.780 2334.860 1687.040 ;
      LAYER met2 ;
        RECT 2334.520 1700.000 2334.800 1702.400 ;
        RECT 2334.660 1687.070 2334.800 1700.000 ;
        RECT 2304.240 1686.750 2304.500 1687.070 ;
        RECT 2334.600 1686.750 2334.860 1687.070 ;
        RECT 2304.300 2.400 2304.440 1686.750 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2324.910 1689.020 2325.230 1689.080 ;
        RECT 2343.770 1689.020 2344.090 1689.080 ;
        RECT 2324.910 1688.880 2344.090 1689.020 ;
        RECT 2324.910 1688.820 2325.230 1688.880 ;
        RECT 2343.770 1688.820 2344.090 1688.880 ;
        RECT 2322.150 16.560 2322.470 16.620 ;
        RECT 2324.910 16.560 2325.230 16.620 ;
        RECT 2322.150 16.420 2325.230 16.560 ;
        RECT 2322.150 16.360 2322.470 16.420 ;
        RECT 2324.910 16.360 2325.230 16.420 ;
      LAYER via ;
        RECT 2324.940 1688.820 2325.200 1689.080 ;
        RECT 2343.800 1688.820 2344.060 1689.080 ;
        RECT 2322.180 16.360 2322.440 16.620 ;
        RECT 2324.940 16.360 2325.200 16.620 ;
      LAYER met2 ;
        RECT 2343.720 1700.000 2344.000 1702.400 ;
        RECT 2343.860 1689.110 2344.000 1700.000 ;
        RECT 2324.940 1688.790 2325.200 1689.110 ;
        RECT 2343.800 1688.790 2344.060 1689.110 ;
        RECT 2325.000 16.650 2325.140 1688.790 ;
        RECT 2322.180 16.330 2322.440 16.650 ;
        RECT 2324.940 16.330 2325.200 16.650 ;
        RECT 2322.240 2.400 2322.380 16.330 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2339.630 17.920 2339.950 17.980 ;
        RECT 2353.890 17.920 2354.210 17.980 ;
        RECT 2339.630 17.780 2354.210 17.920 ;
        RECT 2339.630 17.720 2339.950 17.780 ;
        RECT 2353.890 17.720 2354.210 17.780 ;
      LAYER via ;
        RECT 2339.660 17.720 2339.920 17.980 ;
        RECT 2353.920 17.720 2354.180 17.980 ;
      LAYER met2 ;
        RECT 2352.920 1700.410 2353.200 1702.400 ;
        RECT 2352.920 1700.270 2354.120 1700.410 ;
        RECT 2352.920 1700.000 2353.200 1700.270 ;
        RECT 2353.980 18.010 2354.120 1700.270 ;
        RECT 2339.660 17.690 2339.920 18.010 ;
        RECT 2353.920 17.690 2354.180 18.010 ;
        RECT 2339.720 2.400 2339.860 17.690 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2357.570 14.180 2357.890 14.240 ;
        RECT 2359.410 14.180 2359.730 14.240 ;
        RECT 2357.570 14.040 2359.730 14.180 ;
        RECT 2357.570 13.980 2357.890 14.040 ;
        RECT 2359.410 13.980 2359.730 14.040 ;
      LAYER via ;
        RECT 2357.600 13.980 2357.860 14.240 ;
        RECT 2359.440 13.980 2359.700 14.240 ;
      LAYER met2 ;
        RECT 2362.120 1700.410 2362.400 1702.400 ;
        RECT 2359.960 1700.270 2362.400 1700.410 ;
        RECT 2359.960 1684.090 2360.100 1700.270 ;
        RECT 2362.120 1700.000 2362.400 1700.270 ;
        RECT 2359.500 1683.950 2360.100 1684.090 ;
        RECT 2359.500 14.270 2359.640 1683.950 ;
        RECT 2357.600 13.950 2357.860 14.270 ;
        RECT 2359.440 13.950 2359.700 14.270 ;
        RECT 2357.660 2.400 2357.800 13.950 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2373.210 20.640 2373.530 20.700 ;
        RECT 2375.510 20.640 2375.830 20.700 ;
        RECT 2373.210 20.500 2375.830 20.640 ;
        RECT 2373.210 20.440 2373.530 20.500 ;
        RECT 2375.510 20.440 2375.830 20.500 ;
      LAYER via ;
        RECT 2373.240 20.440 2373.500 20.700 ;
        RECT 2375.540 20.440 2375.800 20.700 ;
      LAYER met2 ;
        RECT 2371.320 1700.410 2371.600 1702.400 ;
        RECT 2371.320 1700.270 2373.440 1700.410 ;
        RECT 2371.320 1700.000 2371.600 1700.270 ;
        RECT 2373.300 20.730 2373.440 1700.270 ;
        RECT 2373.240 20.410 2373.500 20.730 ;
        RECT 2375.540 20.410 2375.800 20.730 ;
        RECT 2375.600 2.400 2375.740 20.410 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2380.570 1684.600 2380.890 1684.660 ;
        RECT 2388.850 1684.600 2389.170 1684.660 ;
        RECT 2380.570 1684.460 2389.170 1684.600 ;
        RECT 2380.570 1684.400 2380.890 1684.460 ;
        RECT 2388.850 1684.400 2389.170 1684.460 ;
        RECT 2388.850 2.960 2389.170 3.020 ;
        RECT 2393.450 2.960 2393.770 3.020 ;
        RECT 2388.850 2.820 2393.770 2.960 ;
        RECT 2388.850 2.760 2389.170 2.820 ;
        RECT 2393.450 2.760 2393.770 2.820 ;
      LAYER via ;
        RECT 2380.600 1684.400 2380.860 1684.660 ;
        RECT 2388.880 1684.400 2389.140 1684.660 ;
        RECT 2388.880 2.760 2389.140 3.020 ;
        RECT 2393.480 2.760 2393.740 3.020 ;
      LAYER met2 ;
        RECT 2380.520 1700.000 2380.800 1702.400 ;
        RECT 2380.660 1684.690 2380.800 1700.000 ;
        RECT 2380.600 1684.370 2380.860 1684.690 ;
        RECT 2388.880 1684.370 2389.140 1684.690 ;
        RECT 2388.940 3.050 2389.080 1684.370 ;
        RECT 2388.880 2.730 2389.140 3.050 ;
        RECT 2393.480 2.730 2393.740 3.050 ;
        RECT 2393.540 2.400 2393.680 2.730 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2389.770 1688.680 2390.090 1688.740 ;
        RECT 2393.910 1688.680 2394.230 1688.740 ;
        RECT 2389.770 1688.540 2394.230 1688.680 ;
        RECT 2389.770 1688.480 2390.090 1688.540 ;
        RECT 2393.910 1688.480 2394.230 1688.540 ;
        RECT 2393.910 18.260 2394.230 18.320 ;
        RECT 2411.390 18.260 2411.710 18.320 ;
        RECT 2393.910 18.120 2411.710 18.260 ;
        RECT 2393.910 18.060 2394.230 18.120 ;
        RECT 2411.390 18.060 2411.710 18.120 ;
      LAYER via ;
        RECT 2389.800 1688.480 2390.060 1688.740 ;
        RECT 2393.940 1688.480 2394.200 1688.740 ;
        RECT 2393.940 18.060 2394.200 18.320 ;
        RECT 2411.420 18.060 2411.680 18.320 ;
      LAYER met2 ;
        RECT 2389.720 1700.000 2390.000 1702.400 ;
        RECT 2389.860 1688.770 2390.000 1700.000 ;
        RECT 2389.800 1688.450 2390.060 1688.770 ;
        RECT 2393.940 1688.450 2394.200 1688.770 ;
        RECT 2394.000 18.350 2394.140 1688.450 ;
        RECT 2393.940 18.030 2394.200 18.350 ;
        RECT 2411.420 18.030 2411.680 18.350 ;
        RECT 2411.480 2.400 2411.620 18.030 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.470 1689.360 1559.790 1689.420 ;
        RECT 1561.310 1689.360 1561.630 1689.420 ;
        RECT 1559.470 1689.220 1561.630 1689.360 ;
        RECT 1559.470 1689.160 1559.790 1689.220 ;
        RECT 1561.310 1689.160 1561.630 1689.220 ;
        RECT 806.910 49.880 807.230 49.940 ;
        RECT 1559.470 49.880 1559.790 49.940 ;
        RECT 806.910 49.740 1559.790 49.880 ;
        RECT 806.910 49.680 807.230 49.740 ;
        RECT 1559.470 49.680 1559.790 49.740 ;
      LAYER via ;
        RECT 1559.500 1689.160 1559.760 1689.420 ;
        RECT 1561.340 1689.160 1561.600 1689.420 ;
        RECT 806.940 49.680 807.200 49.940 ;
        RECT 1559.500 49.680 1559.760 49.940 ;
      LAYER met2 ;
        RECT 1563.100 1700.410 1563.380 1702.400 ;
        RECT 1561.400 1700.270 1563.380 1700.410 ;
        RECT 1561.400 1689.450 1561.540 1700.270 ;
        RECT 1563.100 1700.000 1563.380 1700.270 ;
        RECT 1559.500 1689.130 1559.760 1689.450 ;
        RECT 1561.340 1689.130 1561.600 1689.450 ;
        RECT 1559.560 49.970 1559.700 1689.130 ;
        RECT 806.940 49.650 807.200 49.970 ;
        RECT 1559.500 49.650 1559.760 49.970 ;
        RECT 807.000 16.730 807.140 49.650 ;
        RECT 805.620 16.590 807.140 16.730 ;
        RECT 805.620 2.400 805.760 16.590 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.470 1678.140 1145.790 1678.200 ;
        RECT 1149.150 1678.140 1149.470 1678.200 ;
        RECT 1145.470 1678.000 1149.470 1678.140 ;
        RECT 1145.470 1677.940 1145.790 1678.000 ;
        RECT 1149.150 1677.940 1149.470 1678.000 ;
        RECT 2.830 24.380 3.150 24.440 ;
        RECT 1145.470 24.380 1145.790 24.440 ;
        RECT 2.830 24.240 1145.790 24.380 ;
        RECT 2.830 24.180 3.150 24.240 ;
        RECT 1145.470 24.180 1145.790 24.240 ;
      LAYER via ;
        RECT 1145.500 1677.940 1145.760 1678.200 ;
        RECT 1149.180 1677.940 1149.440 1678.200 ;
        RECT 2.860 24.180 3.120 24.440 ;
        RECT 1145.500 24.180 1145.760 24.440 ;
      LAYER met2 ;
        RECT 1150.020 1700.410 1150.300 1702.400 ;
        RECT 1149.240 1700.270 1150.300 1700.410 ;
        RECT 1149.240 1678.230 1149.380 1700.270 ;
        RECT 1150.020 1700.000 1150.300 1700.270 ;
        RECT 1145.500 1677.910 1145.760 1678.230 ;
        RECT 1149.180 1677.910 1149.440 1678.230 ;
        RECT 1145.560 24.470 1145.700 1677.910 ;
        RECT 2.860 24.150 3.120 24.470 ;
        RECT 1145.500 24.150 1145.760 24.470 ;
        RECT 2.920 2.400 3.060 24.150 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 24.040 8.670 24.100 ;
        RECT 1152.830 24.040 1153.150 24.100 ;
        RECT 8.350 23.900 1153.150 24.040 ;
        RECT 8.350 23.840 8.670 23.900 ;
        RECT 1152.830 23.840 1153.150 23.900 ;
      LAYER via ;
        RECT 8.380 23.840 8.640 24.100 ;
        RECT 1152.860 23.840 1153.120 24.100 ;
      LAYER met2 ;
        RECT 1152.780 1700.000 1153.060 1702.400 ;
        RECT 1152.920 24.130 1153.060 1700.000 ;
        RECT 8.380 23.810 8.640 24.130 ;
        RECT 1152.860 23.810 1153.120 24.130 ;
        RECT 8.440 2.400 8.580 23.810 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1152.370 1678.140 1152.690 1678.200 ;
        RECT 1154.670 1678.140 1154.990 1678.200 ;
        RECT 1152.370 1678.000 1154.990 1678.140 ;
        RECT 1152.370 1677.940 1152.690 1678.000 ;
        RECT 1154.670 1677.940 1154.990 1678.000 ;
        RECT 14.330 24.720 14.650 24.780 ;
        RECT 1152.370 24.720 1152.690 24.780 ;
        RECT 14.330 24.580 1152.690 24.720 ;
        RECT 14.330 24.520 14.650 24.580 ;
        RECT 1152.370 24.520 1152.690 24.580 ;
      LAYER via ;
        RECT 1152.400 1677.940 1152.660 1678.200 ;
        RECT 1154.700 1677.940 1154.960 1678.200 ;
        RECT 14.360 24.520 14.620 24.780 ;
        RECT 1152.400 24.520 1152.660 24.780 ;
      LAYER met2 ;
        RECT 1156.000 1700.410 1156.280 1702.400 ;
        RECT 1154.760 1700.270 1156.280 1700.410 ;
        RECT 1154.760 1678.230 1154.900 1700.270 ;
        RECT 1156.000 1700.000 1156.280 1700.270 ;
        RECT 1152.400 1677.910 1152.660 1678.230 ;
        RECT 1154.700 1677.910 1154.960 1678.230 ;
        RECT 1152.460 24.810 1152.600 1677.910 ;
        RECT 14.360 24.490 14.620 24.810 ;
        RECT 1152.400 24.490 1152.660 24.810 ;
        RECT 14.420 2.400 14.560 24.490 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 1166.170 25.060 1166.490 25.120 ;
        RECT 38.250 24.920 1166.490 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 1166.170 24.860 1166.490 24.920 ;
      LAYER via ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 1166.200 24.860 1166.460 25.120 ;
      LAYER met2 ;
        RECT 1167.960 1700.410 1168.240 1702.400 ;
        RECT 1166.260 1700.270 1168.240 1700.410 ;
        RECT 1166.260 25.150 1166.400 1700.270 ;
        RECT 1167.960 1700.000 1168.240 1700.270 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 1166.200 24.830 1166.460 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1272.380 1700.410 1272.660 1702.400 ;
        RECT 1269.760 1700.270 1272.660 1700.410 ;
        RECT 1269.760 31.125 1269.900 1700.270 ;
        RECT 1272.380 1700.000 1272.660 1700.270 ;
        RECT 240.670 30.755 240.950 31.125 ;
        RECT 1269.690 30.755 1269.970 31.125 ;
        RECT 240.740 2.400 240.880 30.755 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 240.670 30.800 240.950 31.080 ;
        RECT 1269.690 30.800 1269.970 31.080 ;
      LAYER met3 ;
        RECT 240.645 31.090 240.975 31.105 ;
        RECT 1269.665 31.090 1269.995 31.105 ;
        RECT 240.645 30.790 1269.995 31.090 ;
        RECT 240.645 30.775 240.975 30.790 ;
        RECT 1269.665 30.775 1269.995 30.790 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1277.565 1442.025 1277.735 1490.475 ;
        RECT 1277.105 234.685 1277.275 282.795 ;
        RECT 1277.565 137.785 1277.735 224.315 ;
      LAYER mcon ;
        RECT 1277.565 1490.305 1277.735 1490.475 ;
        RECT 1277.105 282.625 1277.275 282.795 ;
        RECT 1277.565 224.145 1277.735 224.315 ;
      LAYER met1 ;
        RECT 1277.030 1587.020 1277.350 1587.080 ;
        RECT 1277.950 1587.020 1278.270 1587.080 ;
        RECT 1277.030 1586.880 1278.270 1587.020 ;
        RECT 1277.030 1586.820 1277.350 1586.880 ;
        RECT 1277.950 1586.820 1278.270 1586.880 ;
        RECT 1277.490 1490.460 1277.810 1490.520 ;
        RECT 1277.295 1490.320 1277.810 1490.460 ;
        RECT 1277.490 1490.260 1277.810 1490.320 ;
        RECT 1277.490 1442.180 1277.810 1442.240 ;
        RECT 1277.295 1442.040 1277.810 1442.180 ;
        RECT 1277.490 1441.980 1277.810 1442.040 ;
        RECT 1277.490 1303.940 1277.810 1304.200 ;
        RECT 1277.580 1303.800 1277.720 1303.940 ;
        RECT 1277.950 1303.800 1278.270 1303.860 ;
        RECT 1277.580 1303.660 1278.270 1303.800 ;
        RECT 1277.950 1303.600 1278.270 1303.660 ;
        RECT 1277.490 821.000 1277.810 821.060 ;
        RECT 1277.950 821.000 1278.270 821.060 ;
        RECT 1277.490 820.860 1278.270 821.000 ;
        RECT 1277.490 820.800 1277.810 820.860 ;
        RECT 1277.950 820.800 1278.270 820.860 ;
        RECT 1277.490 627.880 1277.810 627.940 ;
        RECT 1277.950 627.880 1278.270 627.940 ;
        RECT 1277.490 627.740 1278.270 627.880 ;
        RECT 1277.490 627.680 1277.810 627.740 ;
        RECT 1277.950 627.680 1278.270 627.740 ;
        RECT 1277.045 282.780 1277.335 282.825 ;
        RECT 1277.490 282.780 1277.810 282.840 ;
        RECT 1277.045 282.640 1277.810 282.780 ;
        RECT 1277.045 282.595 1277.335 282.640 ;
        RECT 1277.490 282.580 1277.810 282.640 ;
        RECT 1277.030 234.840 1277.350 234.900 ;
        RECT 1276.835 234.700 1277.350 234.840 ;
        RECT 1277.030 234.640 1277.350 234.700 ;
        RECT 1277.030 224.300 1277.350 224.360 ;
        RECT 1277.505 224.300 1277.795 224.345 ;
        RECT 1277.030 224.160 1277.795 224.300 ;
        RECT 1277.030 224.100 1277.350 224.160 ;
        RECT 1277.505 224.115 1277.795 224.160 ;
        RECT 1276.570 137.940 1276.890 138.000 ;
        RECT 1277.505 137.940 1277.795 137.985 ;
        RECT 1276.570 137.800 1277.795 137.940 ;
        RECT 1276.570 137.740 1276.890 137.800 ;
        RECT 1277.505 137.755 1277.795 137.800 ;
        RECT 258.130 30.840 258.450 30.900 ;
        RECT 1276.570 30.840 1276.890 30.900 ;
        RECT 258.130 30.700 1276.890 30.840 ;
        RECT 258.130 30.640 258.450 30.700 ;
        RECT 1276.570 30.640 1276.890 30.700 ;
      LAYER via ;
        RECT 1277.060 1586.820 1277.320 1587.080 ;
        RECT 1277.980 1586.820 1278.240 1587.080 ;
        RECT 1277.520 1490.260 1277.780 1490.520 ;
        RECT 1277.520 1441.980 1277.780 1442.240 ;
        RECT 1277.520 1303.940 1277.780 1304.200 ;
        RECT 1277.980 1303.600 1278.240 1303.860 ;
        RECT 1277.520 820.800 1277.780 821.060 ;
        RECT 1277.980 820.800 1278.240 821.060 ;
        RECT 1277.520 627.680 1277.780 627.940 ;
        RECT 1277.980 627.680 1278.240 627.940 ;
        RECT 1277.520 282.580 1277.780 282.840 ;
        RECT 1277.060 234.640 1277.320 234.900 ;
        RECT 1277.060 224.100 1277.320 224.360 ;
        RECT 1276.600 137.740 1276.860 138.000 ;
        RECT 258.160 30.640 258.420 30.900 ;
        RECT 1276.600 30.640 1276.860 30.900 ;
      LAYER met2 ;
        RECT 1281.580 1700.410 1281.860 1702.400 ;
        RECT 1279.420 1700.270 1281.860 1700.410 ;
        RECT 1279.420 1656.210 1279.560 1700.270 ;
        RECT 1281.580 1700.000 1281.860 1700.270 ;
        RECT 1277.580 1656.070 1279.560 1656.210 ;
        RECT 1277.580 1587.530 1277.720 1656.070 ;
        RECT 1277.120 1587.390 1277.720 1587.530 ;
        RECT 1277.120 1587.110 1277.260 1587.390 ;
        RECT 1277.060 1586.790 1277.320 1587.110 ;
        RECT 1277.980 1586.790 1278.240 1587.110 ;
        RECT 1278.040 1580.165 1278.180 1586.790 ;
        RECT 1277.970 1579.795 1278.250 1580.165 ;
        RECT 1278.890 1579.795 1279.170 1580.165 ;
        RECT 1278.960 1537.210 1279.100 1579.795 ;
        RECT 1278.040 1537.070 1279.100 1537.210 ;
        RECT 1278.040 1490.970 1278.180 1537.070 ;
        RECT 1277.580 1490.830 1278.180 1490.970 ;
        RECT 1277.580 1490.550 1277.720 1490.830 ;
        RECT 1277.520 1490.230 1277.780 1490.550 ;
        RECT 1277.520 1441.950 1277.780 1442.270 ;
        RECT 1277.580 1366.530 1277.720 1441.950 ;
        RECT 1277.120 1366.390 1277.720 1366.530 ;
        RECT 1277.120 1365.850 1277.260 1366.390 ;
        RECT 1277.120 1365.710 1277.720 1365.850 ;
        RECT 1277.580 1304.230 1277.720 1365.710 ;
        RECT 1277.520 1303.910 1277.780 1304.230 ;
        RECT 1277.980 1303.570 1278.240 1303.890 ;
        RECT 1278.040 1269.290 1278.180 1303.570 ;
        RECT 1277.580 1269.150 1278.180 1269.290 ;
        RECT 1277.580 883.730 1277.720 1269.150 ;
        RECT 1277.120 883.590 1277.720 883.730 ;
        RECT 1277.120 883.050 1277.260 883.590 ;
        RECT 1277.120 882.910 1277.720 883.050 ;
        RECT 1277.580 821.090 1277.720 882.910 ;
        RECT 1277.520 820.770 1277.780 821.090 ;
        RECT 1277.980 820.770 1278.240 821.090 ;
        RECT 1278.040 786.660 1278.180 820.770 ;
        RECT 1277.580 786.520 1278.180 786.660 ;
        RECT 1277.580 690.610 1277.720 786.520 ;
        RECT 1277.120 690.470 1277.720 690.610 ;
        RECT 1277.120 688.570 1277.260 690.470 ;
        RECT 1277.120 688.430 1277.720 688.570 ;
        RECT 1277.580 627.970 1277.720 688.430 ;
        RECT 1277.520 627.650 1277.780 627.970 ;
        RECT 1277.980 627.650 1278.240 627.970 ;
        RECT 1278.040 593.370 1278.180 627.650 ;
        RECT 1277.580 593.230 1278.180 593.370 ;
        RECT 1277.580 303.690 1277.720 593.230 ;
        RECT 1277.120 303.550 1277.720 303.690 ;
        RECT 1277.120 303.010 1277.260 303.550 ;
        RECT 1277.120 302.870 1277.720 303.010 ;
        RECT 1277.580 282.870 1277.720 302.870 ;
        RECT 1277.520 282.550 1277.780 282.870 ;
        RECT 1277.060 234.610 1277.320 234.930 ;
        RECT 1277.120 224.390 1277.260 234.610 ;
        RECT 1277.060 224.070 1277.320 224.390 ;
        RECT 1276.600 137.710 1276.860 138.030 ;
        RECT 1276.660 96.970 1276.800 137.710 ;
        RECT 1276.660 96.830 1277.260 96.970 ;
        RECT 1277.120 62.290 1277.260 96.830 ;
        RECT 1277.120 62.150 1277.720 62.290 ;
        RECT 1277.580 48.520 1277.720 62.150 ;
        RECT 1276.660 48.380 1277.720 48.520 ;
        RECT 1276.660 30.930 1276.800 48.380 ;
        RECT 258.160 30.610 258.420 30.930 ;
        RECT 1276.600 30.610 1276.860 30.930 ;
        RECT 258.220 2.400 258.360 30.610 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 1277.970 1579.840 1278.250 1580.120 ;
        RECT 1278.890 1579.840 1279.170 1580.120 ;
      LAYER met3 ;
        RECT 1277.945 1580.130 1278.275 1580.145 ;
        RECT 1278.865 1580.130 1279.195 1580.145 ;
        RECT 1277.945 1579.830 1279.195 1580.130 ;
        RECT 1277.945 1579.815 1278.275 1579.830 ;
        RECT 1278.865 1579.815 1279.195 1579.830 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 31.180 276.390 31.240 ;
        RECT 1291.290 31.180 1291.610 31.240 ;
        RECT 276.070 31.040 1291.610 31.180 ;
        RECT 276.070 30.980 276.390 31.040 ;
        RECT 1291.290 30.980 1291.610 31.040 ;
      LAYER via ;
        RECT 276.100 30.980 276.360 31.240 ;
        RECT 1291.320 30.980 1291.580 31.240 ;
      LAYER met2 ;
        RECT 1290.780 1700.410 1291.060 1702.400 ;
        RECT 1290.780 1700.270 1291.520 1700.410 ;
        RECT 1290.780 1700.000 1291.060 1700.270 ;
        RECT 1291.380 31.270 1291.520 1700.270 ;
        RECT 276.100 30.950 276.360 31.270 ;
        RECT 1291.320 30.950 1291.580 31.270 ;
        RECT 276.160 2.400 276.300 30.950 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 31.520 294.330 31.580 ;
        RECT 1297.270 31.520 1297.590 31.580 ;
        RECT 294.010 31.380 1297.590 31.520 ;
        RECT 294.010 31.320 294.330 31.380 ;
        RECT 1297.270 31.320 1297.590 31.380 ;
      LAYER via ;
        RECT 294.040 31.320 294.300 31.580 ;
        RECT 1297.300 31.320 1297.560 31.580 ;
      LAYER met2 ;
        RECT 1299.980 1700.410 1300.260 1702.400 ;
        RECT 1297.360 1700.270 1300.260 1700.410 ;
        RECT 1297.360 31.610 1297.500 1700.270 ;
        RECT 1299.980 1700.000 1300.260 1700.270 ;
        RECT 294.040 31.290 294.300 31.610 ;
        RECT 1297.300 31.290 1297.560 31.610 ;
        RECT 294.100 2.400 294.240 31.290 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1304.245 276.165 1304.415 324.275 ;
        RECT 1304.705 58.565 1304.875 62.815 ;
      LAYER mcon ;
        RECT 1304.245 324.105 1304.415 324.275 ;
        RECT 1304.705 62.645 1304.875 62.815 ;
      LAYER met1 ;
        RECT 1305.090 1608.240 1305.410 1608.500 ;
        RECT 1305.180 1607.820 1305.320 1608.240 ;
        RECT 1305.090 1607.560 1305.410 1607.820 ;
        RECT 1305.090 1539.080 1305.410 1539.140 ;
        RECT 1305.550 1539.080 1305.870 1539.140 ;
        RECT 1305.090 1538.940 1305.870 1539.080 ;
        RECT 1305.090 1538.880 1305.410 1538.940 ;
        RECT 1305.550 1538.880 1305.870 1538.940 ;
        RECT 1305.090 1490.800 1305.410 1490.860 ;
        RECT 1306.010 1490.800 1306.330 1490.860 ;
        RECT 1305.090 1490.660 1306.330 1490.800 ;
        RECT 1305.090 1490.600 1305.410 1490.660 ;
        RECT 1306.010 1490.600 1306.330 1490.660 ;
        RECT 1305.090 1490.120 1305.410 1490.180 ;
        RECT 1305.550 1490.120 1305.870 1490.180 ;
        RECT 1305.090 1489.980 1305.870 1490.120 ;
        RECT 1305.090 1489.920 1305.410 1489.980 ;
        RECT 1305.550 1489.920 1305.870 1489.980 ;
        RECT 1305.550 1173.240 1305.870 1173.300 ;
        RECT 1305.180 1173.100 1305.870 1173.240 ;
        RECT 1305.180 1172.960 1305.320 1173.100 ;
        RECT 1305.550 1173.040 1305.870 1173.100 ;
        RECT 1305.090 1172.700 1305.410 1172.960 ;
        RECT 1305.550 980.120 1305.870 980.180 ;
        RECT 1305.180 979.980 1305.870 980.120 ;
        RECT 1305.180 979.840 1305.320 979.980 ;
        RECT 1305.550 979.920 1305.870 979.980 ;
        RECT 1305.090 979.580 1305.410 979.840 ;
        RECT 1305.090 593.680 1305.410 593.940 ;
        RECT 1305.180 593.260 1305.320 593.680 ;
        RECT 1305.090 593.000 1305.410 593.260 ;
        RECT 1304.170 500.380 1304.490 500.440 ;
        RECT 1305.090 500.380 1305.410 500.440 ;
        RECT 1304.170 500.240 1305.410 500.380 ;
        RECT 1304.170 500.180 1304.490 500.240 ;
        RECT 1305.090 500.180 1305.410 500.240 ;
        RECT 1303.710 428.300 1304.030 428.360 ;
        RECT 1303.710 428.160 1305.320 428.300 ;
        RECT 1303.710 428.100 1304.030 428.160 ;
        RECT 1305.180 428.020 1305.320 428.160 ;
        RECT 1305.090 427.760 1305.410 428.020 ;
        RECT 1305.090 380.020 1305.410 380.080 ;
        RECT 1304.260 379.880 1305.410 380.020 ;
        RECT 1304.260 379.400 1304.400 379.880 ;
        RECT 1305.090 379.820 1305.410 379.880 ;
        RECT 1304.170 379.140 1304.490 379.400 ;
        RECT 1304.170 331.740 1304.490 331.800 ;
        RECT 1305.090 331.740 1305.410 331.800 ;
        RECT 1304.170 331.600 1305.410 331.740 ;
        RECT 1304.170 331.540 1304.490 331.600 ;
        RECT 1305.090 331.540 1305.410 331.600 ;
        RECT 1304.185 324.260 1304.475 324.305 ;
        RECT 1305.090 324.260 1305.410 324.320 ;
        RECT 1304.185 324.120 1305.410 324.260 ;
        RECT 1304.185 324.075 1304.475 324.120 ;
        RECT 1305.090 324.060 1305.410 324.120 ;
        RECT 1304.170 276.320 1304.490 276.380 ;
        RECT 1303.975 276.180 1304.490 276.320 ;
        RECT 1304.170 276.120 1304.490 276.180 ;
        RECT 1304.630 96.800 1304.950 96.860 ;
        RECT 1305.090 96.800 1305.410 96.860 ;
        RECT 1304.630 96.660 1305.410 96.800 ;
        RECT 1304.630 96.600 1304.950 96.660 ;
        RECT 1305.090 96.600 1305.410 96.660 ;
        RECT 1304.645 62.800 1304.935 62.845 ;
        RECT 1305.090 62.800 1305.410 62.860 ;
        RECT 1304.645 62.660 1305.410 62.800 ;
        RECT 1304.645 62.615 1304.935 62.660 ;
        RECT 1305.090 62.600 1305.410 62.660 ;
        RECT 1304.630 58.720 1304.950 58.780 ;
        RECT 1304.435 58.580 1304.950 58.720 ;
        RECT 1304.630 58.520 1304.950 58.580 ;
        RECT 311.950 32.200 312.270 32.260 ;
        RECT 1304.630 32.200 1304.950 32.260 ;
        RECT 311.950 32.060 1304.950 32.200 ;
        RECT 311.950 32.000 312.270 32.060 ;
        RECT 1304.630 32.000 1304.950 32.060 ;
      LAYER via ;
        RECT 1305.120 1608.240 1305.380 1608.500 ;
        RECT 1305.120 1607.560 1305.380 1607.820 ;
        RECT 1305.120 1538.880 1305.380 1539.140 ;
        RECT 1305.580 1538.880 1305.840 1539.140 ;
        RECT 1305.120 1490.600 1305.380 1490.860 ;
        RECT 1306.040 1490.600 1306.300 1490.860 ;
        RECT 1305.120 1489.920 1305.380 1490.180 ;
        RECT 1305.580 1489.920 1305.840 1490.180 ;
        RECT 1305.580 1173.040 1305.840 1173.300 ;
        RECT 1305.120 1172.700 1305.380 1172.960 ;
        RECT 1305.580 979.920 1305.840 980.180 ;
        RECT 1305.120 979.580 1305.380 979.840 ;
        RECT 1305.120 593.680 1305.380 593.940 ;
        RECT 1305.120 593.000 1305.380 593.260 ;
        RECT 1304.200 500.180 1304.460 500.440 ;
        RECT 1305.120 500.180 1305.380 500.440 ;
        RECT 1303.740 428.100 1304.000 428.360 ;
        RECT 1305.120 427.760 1305.380 428.020 ;
        RECT 1305.120 379.820 1305.380 380.080 ;
        RECT 1304.200 379.140 1304.460 379.400 ;
        RECT 1304.200 331.540 1304.460 331.800 ;
        RECT 1305.120 331.540 1305.380 331.800 ;
        RECT 1305.120 324.060 1305.380 324.320 ;
        RECT 1304.200 276.120 1304.460 276.380 ;
        RECT 1304.660 96.600 1304.920 96.860 ;
        RECT 1305.120 96.600 1305.380 96.860 ;
        RECT 1305.120 62.600 1305.380 62.860 ;
        RECT 1304.660 58.520 1304.920 58.780 ;
        RECT 311.980 32.000 312.240 32.260 ;
        RECT 1304.660 32.000 1304.920 32.260 ;
      LAYER met2 ;
        RECT 1309.180 1701.090 1309.460 1702.400 ;
        RECT 1306.560 1700.950 1309.460 1701.090 ;
        RECT 1306.560 1677.970 1306.700 1700.950 ;
        RECT 1309.180 1700.000 1309.460 1700.950 ;
        RECT 1305.180 1677.830 1306.700 1677.970 ;
        RECT 1305.180 1608.530 1305.320 1677.830 ;
        RECT 1305.120 1608.210 1305.380 1608.530 ;
        RECT 1305.120 1607.530 1305.380 1607.850 ;
        RECT 1305.180 1595.125 1305.320 1607.530 ;
        RECT 1305.110 1594.755 1305.390 1595.125 ;
        RECT 1305.110 1594.075 1305.390 1594.445 ;
        RECT 1305.180 1559.650 1305.320 1594.075 ;
        RECT 1305.180 1559.510 1305.780 1559.650 ;
        RECT 1305.640 1539.170 1305.780 1559.510 ;
        RECT 1305.120 1538.850 1305.380 1539.170 ;
        RECT 1305.580 1538.850 1305.840 1539.170 ;
        RECT 1305.180 1538.685 1305.320 1538.850 ;
        RECT 1305.110 1538.315 1305.390 1538.685 ;
        RECT 1306.030 1538.315 1306.310 1538.685 ;
        RECT 1306.100 1490.890 1306.240 1538.315 ;
        RECT 1305.120 1490.570 1305.380 1490.890 ;
        RECT 1306.040 1490.570 1306.300 1490.890 ;
        RECT 1305.180 1490.210 1305.320 1490.570 ;
        RECT 1305.120 1489.890 1305.380 1490.210 ;
        RECT 1305.580 1489.890 1305.840 1490.210 ;
        RECT 1305.640 1462.410 1305.780 1489.890 ;
        RECT 1305.180 1462.270 1305.780 1462.410 ;
        RECT 1305.180 1400.700 1305.320 1462.270 ;
        RECT 1304.260 1400.560 1305.320 1400.700 ;
        RECT 1304.260 1364.490 1304.400 1400.560 ;
        RECT 1304.260 1364.350 1305.320 1364.490 ;
        RECT 1305.180 1269.970 1305.320 1364.350 ;
        RECT 1304.720 1269.830 1305.320 1269.970 ;
        RECT 1304.720 1269.290 1304.860 1269.830 ;
        RECT 1304.720 1269.150 1305.320 1269.290 ;
        RECT 1305.180 1207.410 1305.320 1269.150 ;
        RECT 1305.180 1207.270 1305.780 1207.410 ;
        RECT 1305.640 1173.330 1305.780 1207.270 ;
        RECT 1305.580 1173.010 1305.840 1173.330 ;
        RECT 1305.120 1172.670 1305.380 1172.990 ;
        RECT 1305.180 1076.850 1305.320 1172.670 ;
        RECT 1304.720 1076.710 1305.320 1076.850 ;
        RECT 1304.720 1076.170 1304.860 1076.710 ;
        RECT 1304.720 1076.030 1305.320 1076.170 ;
        RECT 1305.180 1014.290 1305.320 1076.030 ;
        RECT 1305.180 1014.150 1305.780 1014.290 ;
        RECT 1305.640 980.210 1305.780 1014.150 ;
        RECT 1305.580 979.890 1305.840 980.210 ;
        RECT 1305.120 979.550 1305.380 979.870 ;
        RECT 1305.180 917.730 1305.320 979.550 ;
        RECT 1304.260 917.590 1305.320 917.730 ;
        RECT 1304.260 881.690 1304.400 917.590 ;
        RECT 1304.260 881.550 1305.320 881.690 ;
        RECT 1305.180 787.170 1305.320 881.550 ;
        RECT 1304.720 787.030 1305.320 787.170 ;
        RECT 1304.720 786.490 1304.860 787.030 ;
        RECT 1304.720 786.350 1305.320 786.490 ;
        RECT 1305.180 593.970 1305.320 786.350 ;
        RECT 1305.120 593.650 1305.380 593.970 ;
        RECT 1305.120 592.970 1305.380 593.290 ;
        RECT 1305.180 500.470 1305.320 592.970 ;
        RECT 1304.200 500.150 1304.460 500.470 ;
        RECT 1305.120 500.150 1305.380 500.470 ;
        RECT 1304.260 452.610 1304.400 500.150 ;
        RECT 1303.800 452.470 1304.400 452.610 ;
        RECT 1303.800 428.390 1303.940 452.470 ;
        RECT 1303.740 428.070 1304.000 428.390 ;
        RECT 1305.120 427.730 1305.380 428.050 ;
        RECT 1305.180 380.110 1305.320 427.730 ;
        RECT 1305.120 379.790 1305.380 380.110 ;
        RECT 1304.200 379.110 1304.460 379.430 ;
        RECT 1304.260 331.830 1304.400 379.110 ;
        RECT 1304.200 331.510 1304.460 331.830 ;
        RECT 1305.120 331.510 1305.380 331.830 ;
        RECT 1305.180 324.350 1305.320 331.510 ;
        RECT 1305.120 324.030 1305.380 324.350 ;
        RECT 1304.200 276.090 1304.460 276.410 ;
        RECT 1304.260 258.130 1304.400 276.090 ;
        RECT 1304.260 257.990 1305.780 258.130 ;
        RECT 1305.640 234.330 1305.780 257.990 ;
        RECT 1304.720 234.190 1305.780 234.330 ;
        RECT 1304.720 203.050 1304.860 234.190 ;
        RECT 1304.720 202.910 1305.320 203.050 ;
        RECT 1305.180 169.050 1305.320 202.910 ;
        RECT 1304.720 168.910 1305.320 169.050 ;
        RECT 1304.720 96.890 1304.860 168.910 ;
        RECT 1304.660 96.570 1304.920 96.890 ;
        RECT 1305.120 96.570 1305.380 96.890 ;
        RECT 1305.180 62.890 1305.320 96.570 ;
        RECT 1305.120 62.570 1305.380 62.890 ;
        RECT 1304.660 58.490 1304.920 58.810 ;
        RECT 1304.720 32.290 1304.860 58.490 ;
        RECT 311.980 31.970 312.240 32.290 ;
        RECT 1304.660 31.970 1304.920 32.290 ;
        RECT 312.040 2.400 312.180 31.970 ;
        RECT 311.830 -4.800 312.390 2.400 ;
      LAYER via2 ;
        RECT 1305.110 1594.800 1305.390 1595.080 ;
        RECT 1305.110 1594.120 1305.390 1594.400 ;
        RECT 1305.110 1538.360 1305.390 1538.640 ;
        RECT 1306.030 1538.360 1306.310 1538.640 ;
      LAYER met3 ;
        RECT 1305.085 1595.090 1305.415 1595.105 ;
        RECT 1304.870 1594.775 1305.415 1595.090 ;
        RECT 1304.870 1594.425 1305.170 1594.775 ;
        RECT 1304.870 1594.110 1305.415 1594.425 ;
        RECT 1305.085 1594.095 1305.415 1594.110 ;
        RECT 1305.085 1538.650 1305.415 1538.665 ;
        RECT 1306.005 1538.650 1306.335 1538.665 ;
        RECT 1305.085 1538.350 1306.335 1538.650 ;
        RECT 1305.085 1538.335 1305.415 1538.350 ;
        RECT 1306.005 1538.335 1306.335 1538.350 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 31.860 330.210 31.920 ;
        RECT 1318.430 31.860 1318.750 31.920 ;
        RECT 329.890 31.720 1318.750 31.860 ;
        RECT 329.890 31.660 330.210 31.720 ;
        RECT 1318.430 31.660 1318.750 31.720 ;
      LAYER via ;
        RECT 329.920 31.660 330.180 31.920 ;
        RECT 1318.460 31.660 1318.720 31.920 ;
      LAYER met2 ;
        RECT 1318.380 1700.000 1318.660 1702.400 ;
        RECT 1318.520 31.950 1318.660 1700.000 ;
        RECT 329.920 31.630 330.180 31.950 ;
        RECT 1318.460 31.630 1318.720 31.950 ;
        RECT 329.980 2.400 330.120 31.630 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 32.540 347.690 32.600 ;
        RECT 1324.870 32.540 1325.190 32.600 ;
        RECT 347.370 32.400 1325.190 32.540 ;
        RECT 347.370 32.340 347.690 32.400 ;
        RECT 1324.870 32.340 1325.190 32.400 ;
      LAYER via ;
        RECT 347.400 32.340 347.660 32.600 ;
        RECT 1324.900 32.340 1325.160 32.600 ;
      LAYER met2 ;
        RECT 1327.120 1700.410 1327.400 1702.400 ;
        RECT 1324.960 1700.270 1327.400 1700.410 ;
        RECT 1324.960 32.630 1325.100 1700.270 ;
        RECT 1327.120 1700.000 1327.400 1700.270 ;
        RECT 347.400 32.310 347.660 32.630 ;
        RECT 1324.900 32.310 1325.160 32.630 ;
        RECT 347.460 2.400 347.600 32.310 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1332.305 916.725 1332.475 959.055 ;
        RECT 1332.305 662.405 1332.475 710.515 ;
      LAYER mcon ;
        RECT 1332.305 958.885 1332.475 959.055 ;
        RECT 1332.305 710.345 1332.475 710.515 ;
      LAYER met1 ;
        RECT 1331.770 966.180 1332.090 966.240 ;
        RECT 1332.690 966.180 1333.010 966.240 ;
        RECT 1331.770 966.040 1333.010 966.180 ;
        RECT 1331.770 965.980 1332.090 966.040 ;
        RECT 1332.690 965.980 1333.010 966.040 ;
        RECT 1332.245 959.040 1332.535 959.085 ;
        RECT 1332.690 959.040 1333.010 959.100 ;
        RECT 1332.245 958.900 1333.010 959.040 ;
        RECT 1332.245 958.855 1332.535 958.900 ;
        RECT 1332.690 958.840 1333.010 958.900 ;
        RECT 1332.230 916.880 1332.550 916.940 ;
        RECT 1332.035 916.740 1332.550 916.880 ;
        RECT 1332.230 916.680 1332.550 916.740 ;
        RECT 1332.230 710.500 1332.550 710.560 ;
        RECT 1332.035 710.360 1332.550 710.500 ;
        RECT 1332.230 710.300 1332.550 710.360 ;
        RECT 1332.245 662.560 1332.535 662.605 ;
        RECT 1332.690 662.560 1333.010 662.620 ;
        RECT 1332.245 662.420 1333.010 662.560 ;
        RECT 1332.245 662.375 1332.535 662.420 ;
        RECT 1332.690 662.360 1333.010 662.420 ;
        RECT 1332.690 627.880 1333.010 627.940 ;
        RECT 1333.610 627.880 1333.930 627.940 ;
        RECT 1332.690 627.740 1333.930 627.880 ;
        RECT 1332.690 627.680 1333.010 627.740 ;
        RECT 1333.610 627.680 1333.930 627.740 ;
        RECT 1332.690 352.480 1333.010 352.540 ;
        RECT 1332.320 352.340 1333.010 352.480 ;
        RECT 1332.320 351.860 1332.460 352.340 ;
        RECT 1332.690 352.280 1333.010 352.340 ;
        RECT 1332.230 351.600 1332.550 351.860 ;
        RECT 1332.230 289.920 1332.550 289.980 ;
        RECT 1332.690 289.920 1333.010 289.980 ;
        RECT 1332.230 289.780 1333.010 289.920 ;
        RECT 1332.230 289.720 1332.550 289.780 ;
        RECT 1332.690 289.720 1333.010 289.780 ;
        RECT 1331.770 144.740 1332.090 144.800 ;
        RECT 1332.690 144.740 1333.010 144.800 ;
        RECT 1331.770 144.600 1333.010 144.740 ;
        RECT 1331.770 144.540 1332.090 144.600 ;
        RECT 1332.690 144.540 1333.010 144.600 ;
        RECT 365.310 32.880 365.630 32.940 ;
        RECT 1331.770 32.880 1332.090 32.940 ;
        RECT 365.310 32.740 1332.090 32.880 ;
        RECT 365.310 32.680 365.630 32.740 ;
        RECT 1331.770 32.680 1332.090 32.740 ;
      LAYER via ;
        RECT 1331.800 965.980 1332.060 966.240 ;
        RECT 1332.720 965.980 1332.980 966.240 ;
        RECT 1332.720 958.840 1332.980 959.100 ;
        RECT 1332.260 916.680 1332.520 916.940 ;
        RECT 1332.260 710.300 1332.520 710.560 ;
        RECT 1332.720 662.360 1332.980 662.620 ;
        RECT 1332.720 627.680 1332.980 627.940 ;
        RECT 1333.640 627.680 1333.900 627.940 ;
        RECT 1332.720 352.280 1332.980 352.540 ;
        RECT 1332.260 351.600 1332.520 351.860 ;
        RECT 1332.260 289.720 1332.520 289.980 ;
        RECT 1332.720 289.720 1332.980 289.980 ;
        RECT 1331.800 144.540 1332.060 144.800 ;
        RECT 1332.720 144.540 1332.980 144.800 ;
        RECT 365.340 32.680 365.600 32.940 ;
        RECT 1331.800 32.680 1332.060 32.940 ;
      LAYER met2 ;
        RECT 1336.320 1701.090 1336.600 1702.400 ;
        RECT 1334.160 1700.950 1336.600 1701.090 ;
        RECT 1334.160 1656.210 1334.300 1700.950 ;
        RECT 1336.320 1700.000 1336.600 1700.950 ;
        RECT 1332.780 1656.070 1334.300 1656.210 ;
        RECT 1332.780 1607.930 1332.920 1656.070 ;
        RECT 1332.320 1607.790 1332.920 1607.930 ;
        RECT 1332.320 1607.250 1332.460 1607.790 ;
        RECT 1332.320 1607.110 1332.920 1607.250 ;
        RECT 1332.780 1463.090 1332.920 1607.110 ;
        RECT 1332.320 1462.950 1332.920 1463.090 ;
        RECT 1332.320 1462.410 1332.460 1462.950 ;
        RECT 1332.320 1462.270 1332.920 1462.410 ;
        RECT 1332.780 1400.700 1332.920 1462.270 ;
        RECT 1331.860 1400.560 1332.920 1400.700 ;
        RECT 1331.860 1363.810 1332.000 1400.560 ;
        RECT 1331.860 1363.670 1332.920 1363.810 ;
        RECT 1332.780 1269.970 1332.920 1363.670 ;
        RECT 1332.320 1269.830 1332.920 1269.970 ;
        RECT 1332.320 1269.290 1332.460 1269.830 ;
        RECT 1332.320 1269.150 1332.920 1269.290 ;
        RECT 1332.780 1076.850 1332.920 1269.150 ;
        RECT 1332.320 1076.710 1332.920 1076.850 ;
        RECT 1332.320 1076.170 1332.460 1076.710 ;
        RECT 1332.320 1076.030 1332.920 1076.170 ;
        RECT 1332.780 1014.405 1332.920 1076.030 ;
        RECT 1331.790 1014.035 1332.070 1014.405 ;
        RECT 1332.710 1014.035 1332.990 1014.405 ;
        RECT 1331.860 966.270 1332.000 1014.035 ;
        RECT 1331.800 965.950 1332.060 966.270 ;
        RECT 1332.720 965.950 1332.980 966.270 ;
        RECT 1332.780 959.130 1332.920 965.950 ;
        RECT 1332.720 958.810 1332.980 959.130 ;
        RECT 1332.260 916.650 1332.520 916.970 ;
        RECT 1332.320 855.170 1332.460 916.650 ;
        RECT 1332.320 855.030 1332.920 855.170 ;
        RECT 1332.780 787.170 1332.920 855.030 ;
        RECT 1332.320 787.030 1332.920 787.170 ;
        RECT 1332.320 786.490 1332.460 787.030 ;
        RECT 1332.320 786.350 1332.920 786.490 ;
        RECT 1332.780 717.810 1332.920 786.350 ;
        RECT 1332.320 717.670 1332.920 717.810 ;
        RECT 1332.320 710.590 1332.460 717.670 ;
        RECT 1332.260 710.270 1332.520 710.590 ;
        RECT 1332.720 662.330 1332.980 662.650 ;
        RECT 1332.780 627.970 1332.920 662.330 ;
        RECT 1332.720 627.650 1332.980 627.970 ;
        RECT 1333.640 627.650 1333.900 627.970 ;
        RECT 1333.700 579.885 1333.840 627.650 ;
        RECT 1333.630 579.515 1333.910 579.885 ;
        RECT 1332.710 578.835 1332.990 579.205 ;
        RECT 1332.780 497.490 1332.920 578.835 ;
        RECT 1332.780 497.350 1333.380 497.490 ;
        RECT 1333.240 486.610 1333.380 497.350 ;
        RECT 1332.780 486.470 1333.380 486.610 ;
        RECT 1332.780 352.570 1332.920 486.470 ;
        RECT 1332.720 352.250 1332.980 352.570 ;
        RECT 1332.260 351.570 1332.520 351.890 ;
        RECT 1332.320 290.010 1332.460 351.570 ;
        RECT 1332.260 289.690 1332.520 290.010 ;
        RECT 1332.720 289.690 1332.980 290.010 ;
        RECT 1332.780 241.810 1332.920 289.690 ;
        RECT 1332.320 241.670 1332.920 241.810 ;
        RECT 1332.320 210.530 1332.460 241.670 ;
        RECT 1332.320 210.390 1332.920 210.530 ;
        RECT 1332.780 144.830 1332.920 210.390 ;
        RECT 1331.800 144.510 1332.060 144.830 ;
        RECT 1332.720 144.510 1332.980 144.830 ;
        RECT 1331.860 96.970 1332.000 144.510 ;
        RECT 1331.860 96.830 1332.460 96.970 ;
        RECT 1332.320 72.490 1332.460 96.830 ;
        RECT 1331.400 72.350 1332.460 72.490 ;
        RECT 1331.400 61.610 1331.540 72.350 ;
        RECT 1331.400 61.470 1332.000 61.610 ;
        RECT 1331.860 32.970 1332.000 61.470 ;
        RECT 365.340 32.650 365.600 32.970 ;
        RECT 1331.800 32.650 1332.060 32.970 ;
        RECT 365.400 2.400 365.540 32.650 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 1331.790 1014.080 1332.070 1014.360 ;
        RECT 1332.710 1014.080 1332.990 1014.360 ;
        RECT 1333.630 579.560 1333.910 579.840 ;
        RECT 1332.710 578.880 1332.990 579.160 ;
      LAYER met3 ;
        RECT 1331.765 1014.370 1332.095 1014.385 ;
        RECT 1332.685 1014.370 1333.015 1014.385 ;
        RECT 1331.765 1014.070 1333.015 1014.370 ;
        RECT 1331.765 1014.055 1332.095 1014.070 ;
        RECT 1332.685 1014.055 1333.015 1014.070 ;
        RECT 1333.605 579.850 1333.935 579.865 ;
        RECT 1332.470 579.550 1333.935 579.850 ;
        RECT 1332.470 579.185 1332.770 579.550 ;
        RECT 1333.605 579.535 1333.935 579.550 ;
        RECT 1332.470 578.870 1333.015 579.185 ;
        RECT 1332.685 578.855 1333.015 578.870 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 33.220 383.570 33.280 ;
        RECT 1345.570 33.220 1345.890 33.280 ;
        RECT 383.250 33.080 1345.890 33.220 ;
        RECT 383.250 33.020 383.570 33.080 ;
        RECT 1345.570 33.020 1345.890 33.080 ;
      LAYER via ;
        RECT 383.280 33.020 383.540 33.280 ;
        RECT 1345.600 33.020 1345.860 33.280 ;
      LAYER met2 ;
        RECT 1345.520 1700.000 1345.800 1702.400 ;
        RECT 1345.660 33.310 1345.800 1700.000 ;
        RECT 383.280 32.990 383.540 33.310 ;
        RECT 1345.600 32.990 1345.860 33.310 ;
        RECT 383.340 2.400 383.480 32.990 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 33.560 401.510 33.620 ;
        RECT 1352.930 33.560 1353.250 33.620 ;
        RECT 401.190 33.420 1353.250 33.560 ;
        RECT 401.190 33.360 401.510 33.420 ;
        RECT 1352.930 33.360 1353.250 33.420 ;
      LAYER via ;
        RECT 401.220 33.360 401.480 33.620 ;
        RECT 1352.960 33.360 1353.220 33.620 ;
      LAYER met2 ;
        RECT 1354.720 1700.410 1355.000 1702.400 ;
        RECT 1352.560 1700.270 1355.000 1700.410 ;
        RECT 1352.560 48.010 1352.700 1700.270 ;
        RECT 1354.720 1700.000 1355.000 1700.270 ;
        RECT 1352.560 47.870 1353.160 48.010 ;
        RECT 1353.020 33.650 1353.160 47.870 ;
        RECT 401.220 33.330 401.480 33.650 ;
        RECT 1352.960 33.330 1353.220 33.650 ;
        RECT 401.280 2.400 401.420 33.330 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 25.400 62.490 25.460 ;
        RECT 1180.430 25.400 1180.750 25.460 ;
        RECT 62.170 25.260 1180.750 25.400 ;
        RECT 62.170 25.200 62.490 25.260 ;
        RECT 1180.430 25.200 1180.750 25.260 ;
      LAYER via ;
        RECT 62.200 25.200 62.460 25.460 ;
        RECT 1180.460 25.200 1180.720 25.460 ;
      LAYER met2 ;
        RECT 1180.380 1700.000 1180.660 1702.400 ;
        RECT 1180.520 25.490 1180.660 1700.000 ;
        RECT 62.200 25.170 62.460 25.490 ;
        RECT 1180.460 25.170 1180.720 25.490 ;
        RECT 62.260 2.400 62.400 25.170 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1359.905 317.645 1360.075 365.755 ;
        RECT 1359.905 227.885 1360.075 292.995 ;
        RECT 1360.365 186.065 1360.535 193.715 ;
        RECT 1359.905 89.845 1360.075 137.955 ;
      LAYER mcon ;
        RECT 1359.905 365.585 1360.075 365.755 ;
        RECT 1359.905 292.825 1360.075 292.995 ;
        RECT 1360.365 193.545 1360.535 193.715 ;
        RECT 1359.905 137.785 1360.075 137.955 ;
      LAYER met1 ;
        RECT 1360.290 1365.820 1360.610 1366.080 ;
        RECT 1360.380 1365.400 1360.520 1365.820 ;
        RECT 1360.290 1365.140 1360.610 1365.400 ;
        RECT 1360.290 1269.260 1360.610 1269.520 ;
        RECT 1360.380 1268.840 1360.520 1269.260 ;
        RECT 1360.290 1268.580 1360.610 1268.840 ;
        RECT 1360.290 1172.700 1360.610 1172.960 ;
        RECT 1360.380 1172.280 1360.520 1172.700 ;
        RECT 1360.290 1172.020 1360.610 1172.280 ;
        RECT 1360.290 1076.140 1360.610 1076.400 ;
        RECT 1360.380 1075.720 1360.520 1076.140 ;
        RECT 1360.290 1075.460 1360.610 1075.720 ;
        RECT 1360.290 821.000 1360.610 821.060 ;
        RECT 1361.210 821.000 1361.530 821.060 ;
        RECT 1360.290 820.860 1361.530 821.000 ;
        RECT 1360.290 820.800 1360.610 820.860 ;
        RECT 1361.210 820.800 1361.530 820.860 ;
        RECT 1358.910 772.720 1359.230 772.780 ;
        RECT 1360.290 772.720 1360.610 772.780 ;
        RECT 1358.910 772.580 1360.610 772.720 ;
        RECT 1358.910 772.520 1359.230 772.580 ;
        RECT 1360.290 772.520 1360.610 772.580 ;
        RECT 1359.830 724.440 1360.150 724.500 ;
        RECT 1360.290 724.440 1360.610 724.500 ;
        RECT 1359.830 724.300 1360.610 724.440 ;
        RECT 1359.830 724.240 1360.150 724.300 ;
        RECT 1360.290 724.240 1360.610 724.300 ;
        RECT 1359.830 652.020 1360.150 652.080 ;
        RECT 1360.750 652.020 1361.070 652.080 ;
        RECT 1359.830 651.880 1361.070 652.020 ;
        RECT 1359.830 651.820 1360.150 651.880 ;
        RECT 1360.750 651.820 1361.070 651.880 ;
        RECT 1360.290 579.940 1360.610 580.000 ;
        RECT 1360.750 579.940 1361.070 580.000 ;
        RECT 1360.290 579.800 1361.070 579.940 ;
        RECT 1360.290 579.740 1360.610 579.800 ;
        RECT 1360.750 579.740 1361.070 579.800 ;
        RECT 1359.830 434.760 1360.150 434.820 ;
        RECT 1360.290 434.760 1360.610 434.820 ;
        RECT 1359.830 434.620 1360.610 434.760 ;
        RECT 1359.830 434.560 1360.150 434.620 ;
        RECT 1360.290 434.560 1360.610 434.620 ;
        RECT 1359.845 365.740 1360.135 365.785 ;
        RECT 1360.290 365.740 1360.610 365.800 ;
        RECT 1359.845 365.600 1360.610 365.740 ;
        RECT 1359.845 365.555 1360.135 365.600 ;
        RECT 1360.290 365.540 1360.610 365.600 ;
        RECT 1359.830 317.800 1360.150 317.860 ;
        RECT 1359.635 317.660 1360.150 317.800 ;
        RECT 1359.830 317.600 1360.150 317.660 ;
        RECT 1359.830 292.980 1360.150 293.040 ;
        RECT 1359.635 292.840 1360.150 292.980 ;
        RECT 1359.830 292.780 1360.150 292.840 ;
        RECT 1359.845 228.040 1360.135 228.085 ;
        RECT 1360.290 228.040 1360.610 228.100 ;
        RECT 1359.845 227.900 1360.610 228.040 ;
        RECT 1359.845 227.855 1360.135 227.900 ;
        RECT 1360.290 227.840 1360.610 227.900 ;
        RECT 1360.290 193.700 1360.610 193.760 ;
        RECT 1360.095 193.560 1360.610 193.700 ;
        RECT 1360.290 193.500 1360.610 193.560 ;
        RECT 1360.290 186.220 1360.610 186.280 ;
        RECT 1360.095 186.080 1360.610 186.220 ;
        RECT 1360.290 186.020 1360.610 186.080 ;
        RECT 1359.845 137.940 1360.135 137.985 ;
        RECT 1360.290 137.940 1360.610 138.000 ;
        RECT 1359.845 137.800 1360.610 137.940 ;
        RECT 1359.845 137.755 1360.135 137.800 ;
        RECT 1360.290 137.740 1360.610 137.800 ;
        RECT 1359.830 90.000 1360.150 90.060 ;
        RECT 1359.635 89.860 1360.150 90.000 ;
        RECT 1359.830 89.800 1360.150 89.860 ;
        RECT 419.130 33.900 419.450 33.960 ;
        RECT 1359.370 33.900 1359.690 33.960 ;
        RECT 419.130 33.760 1359.690 33.900 ;
        RECT 419.130 33.700 419.450 33.760 ;
        RECT 1359.370 33.700 1359.690 33.760 ;
      LAYER via ;
        RECT 1360.320 1365.820 1360.580 1366.080 ;
        RECT 1360.320 1365.140 1360.580 1365.400 ;
        RECT 1360.320 1269.260 1360.580 1269.520 ;
        RECT 1360.320 1268.580 1360.580 1268.840 ;
        RECT 1360.320 1172.700 1360.580 1172.960 ;
        RECT 1360.320 1172.020 1360.580 1172.280 ;
        RECT 1360.320 1076.140 1360.580 1076.400 ;
        RECT 1360.320 1075.460 1360.580 1075.720 ;
        RECT 1360.320 820.800 1360.580 821.060 ;
        RECT 1361.240 820.800 1361.500 821.060 ;
        RECT 1358.940 772.520 1359.200 772.780 ;
        RECT 1360.320 772.520 1360.580 772.780 ;
        RECT 1359.860 724.240 1360.120 724.500 ;
        RECT 1360.320 724.240 1360.580 724.500 ;
        RECT 1359.860 651.820 1360.120 652.080 ;
        RECT 1360.780 651.820 1361.040 652.080 ;
        RECT 1360.320 579.740 1360.580 580.000 ;
        RECT 1360.780 579.740 1361.040 580.000 ;
        RECT 1359.860 434.560 1360.120 434.820 ;
        RECT 1360.320 434.560 1360.580 434.820 ;
        RECT 1360.320 365.540 1360.580 365.800 ;
        RECT 1359.860 317.600 1360.120 317.860 ;
        RECT 1359.860 292.780 1360.120 293.040 ;
        RECT 1360.320 227.840 1360.580 228.100 ;
        RECT 1360.320 193.500 1360.580 193.760 ;
        RECT 1360.320 186.020 1360.580 186.280 ;
        RECT 1360.320 137.740 1360.580 138.000 ;
        RECT 1359.860 89.800 1360.120 90.060 ;
        RECT 419.160 33.700 419.420 33.960 ;
        RECT 1359.400 33.700 1359.660 33.960 ;
      LAYER met2 ;
        RECT 1363.920 1701.090 1364.200 1702.400 ;
        RECT 1361.760 1700.950 1364.200 1701.090 ;
        RECT 1361.760 1677.970 1361.900 1700.950 ;
        RECT 1363.920 1700.000 1364.200 1700.950 ;
        RECT 1360.380 1677.830 1361.900 1677.970 ;
        RECT 1360.380 1607.930 1360.520 1677.830 ;
        RECT 1359.920 1607.790 1360.520 1607.930 ;
        RECT 1359.920 1607.250 1360.060 1607.790 ;
        RECT 1359.920 1607.110 1360.520 1607.250 ;
        RECT 1360.380 1463.090 1360.520 1607.110 ;
        RECT 1359.920 1462.950 1360.520 1463.090 ;
        RECT 1359.920 1462.410 1360.060 1462.950 ;
        RECT 1359.920 1462.270 1360.520 1462.410 ;
        RECT 1360.380 1366.110 1360.520 1462.270 ;
        RECT 1360.320 1365.790 1360.580 1366.110 ;
        RECT 1360.320 1365.110 1360.580 1365.430 ;
        RECT 1360.380 1269.550 1360.520 1365.110 ;
        RECT 1360.320 1269.230 1360.580 1269.550 ;
        RECT 1360.320 1268.550 1360.580 1268.870 ;
        RECT 1360.380 1172.990 1360.520 1268.550 ;
        RECT 1360.320 1172.670 1360.580 1172.990 ;
        RECT 1360.320 1171.990 1360.580 1172.310 ;
        RECT 1360.380 1076.430 1360.520 1171.990 ;
        RECT 1360.320 1076.110 1360.580 1076.430 ;
        RECT 1360.320 1075.430 1360.580 1075.750 ;
        RECT 1360.380 980.290 1360.520 1075.430 ;
        RECT 1359.920 980.150 1360.520 980.290 ;
        RECT 1359.920 979.610 1360.060 980.150 ;
        RECT 1359.920 979.470 1360.520 979.610 ;
        RECT 1360.380 942.210 1360.520 979.470 ;
        RECT 1359.920 942.070 1360.520 942.210 ;
        RECT 1359.920 917.845 1360.060 942.070 ;
        RECT 1359.850 917.475 1360.130 917.845 ;
        RECT 1361.230 916.795 1361.510 917.165 ;
        RECT 1361.300 821.285 1361.440 916.795 ;
        RECT 1360.310 820.915 1360.590 821.285 ;
        RECT 1361.230 820.915 1361.510 821.285 ;
        RECT 1360.320 820.770 1360.580 820.915 ;
        RECT 1361.240 820.770 1361.500 820.915 ;
        RECT 1361.300 773.005 1361.440 820.770 ;
        RECT 1358.940 772.490 1359.200 772.810 ;
        RECT 1360.310 772.635 1360.590 773.005 ;
        RECT 1361.230 772.635 1361.510 773.005 ;
        RECT 1360.320 772.490 1360.580 772.635 ;
        RECT 1359.000 724.725 1359.140 772.490 ;
        RECT 1358.930 724.355 1359.210 724.725 ;
        RECT 1359.850 724.355 1360.130 724.725 ;
        RECT 1359.860 724.210 1360.120 724.355 ;
        RECT 1360.320 724.210 1360.580 724.530 ;
        RECT 1360.380 699.450 1360.520 724.210 ;
        RECT 1359.920 699.310 1360.520 699.450 ;
        RECT 1359.920 652.110 1360.060 699.310 ;
        RECT 1359.860 651.790 1360.120 652.110 ;
        RECT 1360.780 651.790 1361.040 652.110 ;
        RECT 1360.840 580.030 1360.980 651.790 ;
        RECT 1360.320 579.710 1360.580 580.030 ;
        RECT 1360.780 579.710 1361.040 580.030 ;
        RECT 1360.380 483.890 1360.520 579.710 ;
        RECT 1359.920 483.750 1360.520 483.890 ;
        RECT 1359.920 483.210 1360.060 483.750 ;
        RECT 1359.920 483.070 1360.520 483.210 ;
        RECT 1360.380 434.850 1360.520 483.070 ;
        RECT 1359.860 434.530 1360.120 434.850 ;
        RECT 1360.320 434.530 1360.580 434.850 ;
        RECT 1359.920 366.250 1360.060 434.530 ;
        RECT 1359.920 366.110 1360.520 366.250 ;
        RECT 1360.380 365.830 1360.520 366.110 ;
        RECT 1360.320 365.510 1360.580 365.830 ;
        RECT 1359.860 317.570 1360.120 317.890 ;
        RECT 1359.920 293.070 1360.060 317.570 ;
        RECT 1359.860 292.750 1360.120 293.070 ;
        RECT 1360.320 227.810 1360.580 228.130 ;
        RECT 1360.380 193.790 1360.520 227.810 ;
        RECT 1360.320 193.470 1360.580 193.790 ;
        RECT 1360.320 185.990 1360.580 186.310 ;
        RECT 1360.380 138.030 1360.520 185.990 ;
        RECT 1360.320 137.710 1360.580 138.030 ;
        RECT 1359.860 89.770 1360.120 90.090 ;
        RECT 1359.920 72.490 1360.060 89.770 ;
        RECT 1359.000 72.350 1360.060 72.490 ;
        RECT 1359.000 61.610 1359.140 72.350 ;
        RECT 1359.000 61.470 1359.600 61.610 ;
        RECT 1359.460 33.990 1359.600 61.470 ;
        RECT 419.160 33.670 419.420 33.990 ;
        RECT 1359.400 33.670 1359.660 33.990 ;
        RECT 419.220 2.400 419.360 33.670 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 1359.850 917.520 1360.130 917.800 ;
        RECT 1361.230 916.840 1361.510 917.120 ;
        RECT 1360.310 820.960 1360.590 821.240 ;
        RECT 1361.230 820.960 1361.510 821.240 ;
        RECT 1360.310 772.680 1360.590 772.960 ;
        RECT 1361.230 772.680 1361.510 772.960 ;
        RECT 1358.930 724.400 1359.210 724.680 ;
        RECT 1359.850 724.400 1360.130 724.680 ;
      LAYER met3 ;
        RECT 1359.825 917.810 1360.155 917.825 ;
        RECT 1359.150 917.510 1360.155 917.810 ;
        RECT 1359.150 917.130 1359.450 917.510 ;
        RECT 1359.825 917.495 1360.155 917.510 ;
        RECT 1361.205 917.130 1361.535 917.145 ;
        RECT 1359.150 916.830 1361.535 917.130 ;
        RECT 1361.205 916.815 1361.535 916.830 ;
        RECT 1360.285 821.250 1360.615 821.265 ;
        RECT 1361.205 821.250 1361.535 821.265 ;
        RECT 1360.285 820.950 1361.535 821.250 ;
        RECT 1360.285 820.935 1360.615 820.950 ;
        RECT 1361.205 820.935 1361.535 820.950 ;
        RECT 1360.285 772.970 1360.615 772.985 ;
        RECT 1361.205 772.970 1361.535 772.985 ;
        RECT 1360.285 772.670 1361.535 772.970 ;
        RECT 1360.285 772.655 1360.615 772.670 ;
        RECT 1361.205 772.655 1361.535 772.670 ;
        RECT 1358.905 724.690 1359.235 724.705 ;
        RECT 1359.825 724.690 1360.155 724.705 ;
        RECT 1358.905 724.390 1360.155 724.690 ;
        RECT 1358.905 724.375 1359.235 724.390 ;
        RECT 1359.825 724.375 1360.155 724.390 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 37.640 436.930 37.700 ;
        RECT 1373.170 37.640 1373.490 37.700 ;
        RECT 436.610 37.500 1373.490 37.640 ;
        RECT 436.610 37.440 436.930 37.500 ;
        RECT 1373.170 37.440 1373.490 37.500 ;
      LAYER via ;
        RECT 436.640 37.440 436.900 37.700 ;
        RECT 1373.200 37.440 1373.460 37.700 ;
      LAYER met2 ;
        RECT 1373.120 1700.000 1373.400 1702.400 ;
        RECT 1373.260 37.730 1373.400 1700.000 ;
        RECT 436.640 37.410 436.900 37.730 ;
        RECT 1373.200 37.410 1373.460 37.730 ;
        RECT 436.700 2.400 436.840 37.410 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 37.300 454.870 37.360 ;
        RECT 1380.070 37.300 1380.390 37.360 ;
        RECT 454.550 37.160 1380.390 37.300 ;
        RECT 454.550 37.100 454.870 37.160 ;
        RECT 1380.070 37.100 1380.390 37.160 ;
      LAYER via ;
        RECT 454.580 37.100 454.840 37.360 ;
        RECT 1380.100 37.100 1380.360 37.360 ;
      LAYER met2 ;
        RECT 1382.320 1700.410 1382.600 1702.400 ;
        RECT 1380.160 1700.270 1382.600 1700.410 ;
        RECT 1380.160 37.390 1380.300 1700.270 ;
        RECT 1382.320 1700.000 1382.600 1700.270 ;
        RECT 454.580 37.070 454.840 37.390 ;
        RECT 1380.100 37.070 1380.360 37.390 ;
        RECT 454.640 2.400 454.780 37.070 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1387.965 1531.785 1388.135 1559.495 ;
        RECT 1387.965 1400.885 1388.135 1490.475 ;
        RECT 1388.425 1345.465 1388.595 1375.555 ;
        RECT 1387.045 351.645 1387.215 386.155 ;
        RECT 1387.965 179.605 1388.135 227.715 ;
        RECT 1387.505 83.045 1387.675 131.155 ;
      LAYER mcon ;
        RECT 1387.965 1559.325 1388.135 1559.495 ;
        RECT 1387.965 1490.305 1388.135 1490.475 ;
        RECT 1388.425 1375.385 1388.595 1375.555 ;
        RECT 1387.045 385.985 1387.215 386.155 ;
        RECT 1387.965 227.545 1388.135 227.715 ;
        RECT 1387.505 130.985 1387.675 131.155 ;
      LAYER met1 ;
        RECT 1388.350 1580.220 1388.670 1580.280 ;
        RECT 1389.270 1580.220 1389.590 1580.280 ;
        RECT 1388.350 1580.080 1389.590 1580.220 ;
        RECT 1388.350 1580.020 1388.670 1580.080 ;
        RECT 1389.270 1580.020 1389.590 1580.080 ;
        RECT 1387.890 1559.480 1388.210 1559.540 ;
        RECT 1387.695 1559.340 1388.210 1559.480 ;
        RECT 1387.890 1559.280 1388.210 1559.340 ;
        RECT 1387.890 1531.940 1388.210 1532.000 ;
        RECT 1387.695 1531.800 1388.210 1531.940 ;
        RECT 1387.890 1531.740 1388.210 1531.800 ;
        RECT 1387.890 1497.740 1388.210 1498.000 ;
        RECT 1387.980 1497.320 1388.120 1497.740 ;
        RECT 1387.890 1497.060 1388.210 1497.320 ;
        RECT 1387.890 1490.460 1388.210 1490.520 ;
        RECT 1387.695 1490.320 1388.210 1490.460 ;
        RECT 1387.890 1490.260 1388.210 1490.320 ;
        RECT 1387.905 1401.040 1388.195 1401.085 ;
        RECT 1388.350 1401.040 1388.670 1401.100 ;
        RECT 1387.905 1400.900 1388.670 1401.040 ;
        RECT 1387.905 1400.855 1388.195 1400.900 ;
        RECT 1388.350 1400.840 1388.670 1400.900 ;
        RECT 1388.350 1375.540 1388.670 1375.600 ;
        RECT 1388.155 1375.400 1388.670 1375.540 ;
        RECT 1388.350 1375.340 1388.670 1375.400 ;
        RECT 1388.365 1345.620 1388.655 1345.665 ;
        RECT 1388.810 1345.620 1389.130 1345.680 ;
        RECT 1388.365 1345.480 1389.130 1345.620 ;
        RECT 1388.365 1345.435 1388.655 1345.480 ;
        RECT 1388.810 1345.420 1389.130 1345.480 ;
        RECT 1387.890 1304.140 1388.210 1304.200 ;
        RECT 1388.350 1304.140 1388.670 1304.200 ;
        RECT 1387.890 1304.000 1388.670 1304.140 ;
        RECT 1387.890 1303.940 1388.210 1304.000 ;
        RECT 1388.350 1303.940 1388.670 1304.000 ;
        RECT 1387.890 1159.300 1388.210 1159.360 ;
        RECT 1388.350 1159.300 1388.670 1159.360 ;
        RECT 1387.890 1159.160 1388.670 1159.300 ;
        RECT 1387.890 1159.100 1388.210 1159.160 ;
        RECT 1388.350 1159.100 1388.670 1159.160 ;
        RECT 1387.890 1062.740 1388.210 1062.800 ;
        RECT 1388.350 1062.740 1388.670 1062.800 ;
        RECT 1387.890 1062.600 1388.670 1062.740 ;
        RECT 1387.890 1062.540 1388.210 1062.600 ;
        RECT 1388.350 1062.540 1388.670 1062.600 ;
        RECT 1387.430 979.780 1387.750 979.840 ;
        RECT 1388.350 979.780 1388.670 979.840 ;
        RECT 1387.430 979.640 1388.670 979.780 ;
        RECT 1387.430 979.580 1387.750 979.640 ;
        RECT 1388.350 979.580 1388.670 979.640 ;
        RECT 1387.890 917.900 1388.210 917.960 ;
        RECT 1388.350 917.900 1388.670 917.960 ;
        RECT 1387.890 917.760 1388.670 917.900 ;
        RECT 1387.890 917.700 1388.210 917.760 ;
        RECT 1388.350 917.700 1388.670 917.760 ;
        RECT 1387.890 883.020 1388.210 883.280 ;
        RECT 1387.980 882.600 1388.120 883.020 ;
        RECT 1387.890 882.340 1388.210 882.600 ;
        RECT 1387.890 690.240 1388.210 690.500 ;
        RECT 1387.980 689.820 1388.120 690.240 ;
        RECT 1387.890 689.560 1388.210 689.820 ;
        RECT 1387.890 496.780 1388.210 497.040 ;
        RECT 1387.980 496.640 1388.120 496.780 ;
        RECT 1388.350 496.640 1388.670 496.700 ;
        RECT 1387.980 496.500 1388.670 496.640 ;
        RECT 1388.350 496.440 1388.670 496.500 ;
        RECT 1387.430 400.760 1387.750 400.820 ;
        RECT 1387.060 400.620 1387.750 400.760 ;
        RECT 1387.060 400.140 1387.200 400.620 ;
        RECT 1387.430 400.560 1387.750 400.620 ;
        RECT 1386.970 399.880 1387.290 400.140 ;
        RECT 1386.970 386.140 1387.290 386.200 ;
        RECT 1386.775 386.000 1387.290 386.140 ;
        RECT 1386.970 385.940 1387.290 386.000 ;
        RECT 1386.985 351.800 1387.275 351.845 ;
        RECT 1387.430 351.800 1387.750 351.860 ;
        RECT 1386.985 351.660 1387.750 351.800 ;
        RECT 1386.985 351.615 1387.275 351.660 ;
        RECT 1387.430 351.600 1387.750 351.660 ;
        RECT 1387.890 289.380 1388.210 289.640 ;
        RECT 1387.980 289.240 1388.120 289.380 ;
        RECT 1388.350 289.240 1388.670 289.300 ;
        RECT 1387.980 289.100 1388.670 289.240 ;
        RECT 1388.350 289.040 1388.670 289.100 ;
        RECT 1387.430 282.780 1387.750 282.840 ;
        RECT 1388.350 282.780 1388.670 282.840 ;
        RECT 1387.430 282.640 1388.670 282.780 ;
        RECT 1387.430 282.580 1387.750 282.640 ;
        RECT 1388.350 282.580 1388.670 282.640 ;
        RECT 1387.890 227.700 1388.210 227.760 ;
        RECT 1387.695 227.560 1388.210 227.700 ;
        RECT 1387.890 227.500 1388.210 227.560 ;
        RECT 1387.890 179.760 1388.210 179.820 ;
        RECT 1387.695 179.620 1388.210 179.760 ;
        RECT 1387.890 179.560 1388.210 179.620 ;
        RECT 1387.890 138.620 1388.210 138.680 ;
        RECT 1388.350 138.620 1388.670 138.680 ;
        RECT 1387.890 138.480 1388.670 138.620 ;
        RECT 1387.890 138.420 1388.210 138.480 ;
        RECT 1388.350 138.420 1388.670 138.480 ;
        RECT 1387.445 131.140 1387.735 131.185 ;
        RECT 1387.890 131.140 1388.210 131.200 ;
        RECT 1387.445 131.000 1388.210 131.140 ;
        RECT 1387.445 130.955 1387.735 131.000 ;
        RECT 1387.890 130.940 1388.210 131.000 ;
        RECT 1387.430 83.200 1387.750 83.260 ;
        RECT 1387.235 83.060 1387.750 83.200 ;
        RECT 1387.430 83.000 1387.750 83.060 ;
        RECT 472.490 36.960 472.810 37.020 ;
        RECT 1387.890 36.960 1388.210 37.020 ;
        RECT 472.490 36.820 1388.210 36.960 ;
        RECT 472.490 36.760 472.810 36.820 ;
        RECT 1387.890 36.760 1388.210 36.820 ;
      LAYER via ;
        RECT 1388.380 1580.020 1388.640 1580.280 ;
        RECT 1389.300 1580.020 1389.560 1580.280 ;
        RECT 1387.920 1559.280 1388.180 1559.540 ;
        RECT 1387.920 1531.740 1388.180 1532.000 ;
        RECT 1387.920 1497.740 1388.180 1498.000 ;
        RECT 1387.920 1497.060 1388.180 1497.320 ;
        RECT 1387.920 1490.260 1388.180 1490.520 ;
        RECT 1388.380 1400.840 1388.640 1401.100 ;
        RECT 1388.380 1375.340 1388.640 1375.600 ;
        RECT 1388.840 1345.420 1389.100 1345.680 ;
        RECT 1387.920 1303.940 1388.180 1304.200 ;
        RECT 1388.380 1303.940 1388.640 1304.200 ;
        RECT 1387.920 1159.100 1388.180 1159.360 ;
        RECT 1388.380 1159.100 1388.640 1159.360 ;
        RECT 1387.920 1062.540 1388.180 1062.800 ;
        RECT 1388.380 1062.540 1388.640 1062.800 ;
        RECT 1387.460 979.580 1387.720 979.840 ;
        RECT 1388.380 979.580 1388.640 979.840 ;
        RECT 1387.920 917.700 1388.180 917.960 ;
        RECT 1388.380 917.700 1388.640 917.960 ;
        RECT 1387.920 883.020 1388.180 883.280 ;
        RECT 1387.920 882.340 1388.180 882.600 ;
        RECT 1387.920 690.240 1388.180 690.500 ;
        RECT 1387.920 689.560 1388.180 689.820 ;
        RECT 1387.920 496.780 1388.180 497.040 ;
        RECT 1388.380 496.440 1388.640 496.700 ;
        RECT 1387.460 400.560 1387.720 400.820 ;
        RECT 1387.000 399.880 1387.260 400.140 ;
        RECT 1387.000 385.940 1387.260 386.200 ;
        RECT 1387.460 351.600 1387.720 351.860 ;
        RECT 1387.920 289.380 1388.180 289.640 ;
        RECT 1388.380 289.040 1388.640 289.300 ;
        RECT 1387.460 282.580 1387.720 282.840 ;
        RECT 1388.380 282.580 1388.640 282.840 ;
        RECT 1387.920 227.500 1388.180 227.760 ;
        RECT 1387.920 179.560 1388.180 179.820 ;
        RECT 1387.920 138.420 1388.180 138.680 ;
        RECT 1388.380 138.420 1388.640 138.680 ;
        RECT 1387.920 130.940 1388.180 131.200 ;
        RECT 1387.460 83.000 1387.720 83.260 ;
        RECT 472.520 36.760 472.780 37.020 ;
        RECT 1387.920 36.760 1388.180 37.020 ;
      LAYER met2 ;
        RECT 1391.520 1700.410 1391.800 1702.400 ;
        RECT 1389.820 1700.270 1391.800 1700.410 ;
        RECT 1389.820 1676.725 1389.960 1700.270 ;
        RECT 1391.520 1700.000 1391.800 1700.270 ;
        RECT 1388.370 1676.355 1388.650 1676.725 ;
        RECT 1389.750 1676.355 1390.030 1676.725 ;
        RECT 1388.440 1628.445 1388.580 1676.355 ;
        RECT 1388.370 1628.075 1388.650 1628.445 ;
        RECT 1389.290 1628.075 1389.570 1628.445 ;
        RECT 1388.440 1580.310 1388.580 1580.465 ;
        RECT 1389.360 1580.310 1389.500 1628.075 ;
        RECT 1388.380 1580.050 1388.640 1580.310 ;
        RECT 1387.980 1579.990 1388.640 1580.050 ;
        RECT 1389.300 1579.990 1389.560 1580.310 ;
        RECT 1387.980 1579.910 1388.580 1579.990 ;
        RECT 1387.980 1559.570 1388.120 1579.910 ;
        RECT 1387.920 1559.250 1388.180 1559.570 ;
        RECT 1387.920 1531.710 1388.180 1532.030 ;
        RECT 1387.980 1498.030 1388.120 1531.710 ;
        RECT 1387.920 1497.710 1388.180 1498.030 ;
        RECT 1387.920 1497.030 1388.180 1497.350 ;
        RECT 1387.980 1490.550 1388.120 1497.030 ;
        RECT 1387.920 1490.230 1388.180 1490.550 ;
        RECT 1388.380 1400.810 1388.640 1401.130 ;
        RECT 1388.440 1375.630 1388.580 1400.810 ;
        RECT 1388.380 1375.310 1388.640 1375.630 ;
        RECT 1388.840 1345.390 1389.100 1345.710 ;
        RECT 1388.900 1327.770 1389.040 1345.390 ;
        RECT 1387.980 1327.630 1389.040 1327.770 ;
        RECT 1387.980 1304.230 1388.120 1327.630 ;
        RECT 1387.920 1303.910 1388.180 1304.230 ;
        RECT 1388.380 1303.910 1388.640 1304.230 ;
        RECT 1388.440 1221.010 1388.580 1303.910 ;
        RECT 1387.980 1220.870 1388.580 1221.010 ;
        RECT 1387.980 1159.390 1388.120 1220.870 ;
        RECT 1387.920 1159.070 1388.180 1159.390 ;
        RECT 1388.380 1159.070 1388.640 1159.390 ;
        RECT 1388.440 1124.450 1388.580 1159.070 ;
        RECT 1387.980 1124.310 1388.580 1124.450 ;
        RECT 1387.980 1062.830 1388.120 1124.310 ;
        RECT 1387.920 1062.510 1388.180 1062.830 ;
        RECT 1388.380 1062.510 1388.640 1062.830 ;
        RECT 1388.440 1027.890 1388.580 1062.510 ;
        RECT 1387.980 1027.750 1388.580 1027.890 ;
        RECT 1387.980 980.290 1388.120 1027.750 ;
        RECT 1387.520 980.150 1388.120 980.290 ;
        RECT 1387.520 979.870 1387.660 980.150 ;
        RECT 1387.460 979.550 1387.720 979.870 ;
        RECT 1388.380 979.550 1388.640 979.870 ;
        RECT 1388.440 917.990 1388.580 979.550 ;
        RECT 1387.920 917.670 1388.180 917.990 ;
        RECT 1388.380 917.670 1388.640 917.990 ;
        RECT 1387.980 883.310 1388.120 917.670 ;
        RECT 1387.920 882.990 1388.180 883.310 ;
        RECT 1387.920 882.310 1388.180 882.630 ;
        RECT 1387.980 834.770 1388.120 882.310 ;
        RECT 1387.060 834.630 1388.120 834.770 ;
        RECT 1387.060 773.005 1387.200 834.630 ;
        RECT 1386.990 772.635 1387.270 773.005 ;
        RECT 1388.370 772.635 1388.650 773.005 ;
        RECT 1388.440 738.210 1388.580 772.635 ;
        RECT 1387.980 738.070 1388.580 738.210 ;
        RECT 1387.980 690.530 1388.120 738.070 ;
        RECT 1387.920 690.210 1388.180 690.530 ;
        RECT 1387.920 689.530 1388.180 689.850 ;
        RECT 1387.980 592.690 1388.120 689.530 ;
        RECT 1387.980 592.550 1388.580 592.690 ;
        RECT 1388.440 545.090 1388.580 592.550 ;
        RECT 1387.980 544.950 1388.580 545.090 ;
        RECT 1387.980 497.070 1388.120 544.950 ;
        RECT 1387.920 496.750 1388.180 497.070 ;
        RECT 1388.380 496.410 1388.640 496.730 ;
        RECT 1388.440 448.530 1388.580 496.410 ;
        RECT 1387.520 448.390 1388.580 448.530 ;
        RECT 1387.520 400.850 1387.660 448.390 ;
        RECT 1387.460 400.530 1387.720 400.850 ;
        RECT 1387.000 399.850 1387.260 400.170 ;
        RECT 1387.060 386.230 1387.200 399.850 ;
        RECT 1387.000 385.910 1387.260 386.230 ;
        RECT 1387.460 351.570 1387.720 351.890 ;
        RECT 1387.520 303.010 1387.660 351.570 ;
        RECT 1387.520 302.870 1388.120 303.010 ;
        RECT 1387.980 289.670 1388.120 302.870 ;
        RECT 1387.920 289.350 1388.180 289.670 ;
        RECT 1388.380 289.010 1388.640 289.330 ;
        RECT 1388.440 282.870 1388.580 289.010 ;
        RECT 1387.460 282.550 1387.720 282.870 ;
        RECT 1388.380 282.550 1388.640 282.870 ;
        RECT 1387.520 235.010 1387.660 282.550 ;
        RECT 1387.520 234.870 1388.120 235.010 ;
        RECT 1387.980 227.790 1388.120 234.870 ;
        RECT 1387.920 227.470 1388.180 227.790 ;
        RECT 1387.920 179.530 1388.180 179.850 ;
        RECT 1387.980 144.570 1388.120 179.530 ;
        RECT 1387.980 144.430 1388.580 144.570 ;
        RECT 1388.440 138.710 1388.580 144.430 ;
        RECT 1387.920 138.390 1388.180 138.710 ;
        RECT 1388.380 138.390 1388.640 138.710 ;
        RECT 1387.980 131.230 1388.120 138.390 ;
        RECT 1387.920 130.910 1388.180 131.230 ;
        RECT 1387.460 82.970 1387.720 83.290 ;
        RECT 1387.520 42.685 1387.660 82.970 ;
        RECT 1387.450 42.315 1387.730 42.685 ;
        RECT 1387.910 41.635 1388.190 42.005 ;
        RECT 1387.980 37.050 1388.120 41.635 ;
        RECT 472.520 36.730 472.780 37.050 ;
        RECT 1387.920 36.730 1388.180 37.050 ;
        RECT 472.580 2.400 472.720 36.730 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 1388.370 1676.400 1388.650 1676.680 ;
        RECT 1389.750 1676.400 1390.030 1676.680 ;
        RECT 1388.370 1628.120 1388.650 1628.400 ;
        RECT 1389.290 1628.120 1389.570 1628.400 ;
        RECT 1386.990 772.680 1387.270 772.960 ;
        RECT 1388.370 772.680 1388.650 772.960 ;
        RECT 1387.450 42.360 1387.730 42.640 ;
        RECT 1387.910 41.680 1388.190 41.960 ;
      LAYER met3 ;
        RECT 1388.345 1676.690 1388.675 1676.705 ;
        RECT 1389.725 1676.690 1390.055 1676.705 ;
        RECT 1388.345 1676.390 1390.055 1676.690 ;
        RECT 1388.345 1676.375 1388.675 1676.390 ;
        RECT 1389.725 1676.375 1390.055 1676.390 ;
        RECT 1388.345 1628.410 1388.675 1628.425 ;
        RECT 1389.265 1628.410 1389.595 1628.425 ;
        RECT 1388.345 1628.110 1389.595 1628.410 ;
        RECT 1388.345 1628.095 1388.675 1628.110 ;
        RECT 1389.265 1628.095 1389.595 1628.110 ;
        RECT 1386.965 772.970 1387.295 772.985 ;
        RECT 1388.345 772.970 1388.675 772.985 ;
        RECT 1386.965 772.670 1388.675 772.970 ;
        RECT 1386.965 772.655 1387.295 772.670 ;
        RECT 1388.345 772.655 1388.675 772.670 ;
        RECT 1387.425 42.650 1387.755 42.665 ;
        RECT 1387.425 42.350 1388.890 42.650 ;
        RECT 1387.425 42.335 1387.755 42.350 ;
        RECT 1387.885 41.970 1388.215 41.985 ;
        RECT 1388.590 41.970 1388.890 42.350 ;
        RECT 1387.885 41.670 1388.890 41.970 ;
        RECT 1387.885 41.655 1388.215 41.670 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 495.950 51.920 496.270 51.980 ;
        RECT 1400.770 51.920 1401.090 51.980 ;
        RECT 495.950 51.780 1401.090 51.920 ;
        RECT 495.950 51.720 496.270 51.780 ;
        RECT 1400.770 51.720 1401.090 51.780 ;
        RECT 490.430 15.540 490.750 15.600 ;
        RECT 495.950 15.540 496.270 15.600 ;
        RECT 490.430 15.400 496.270 15.540 ;
        RECT 490.430 15.340 490.750 15.400 ;
        RECT 495.950 15.340 496.270 15.400 ;
      LAYER via ;
        RECT 495.980 51.720 496.240 51.980 ;
        RECT 1400.800 51.720 1401.060 51.980 ;
        RECT 490.460 15.340 490.720 15.600 ;
        RECT 495.980 15.340 496.240 15.600 ;
      LAYER met2 ;
        RECT 1400.720 1700.000 1401.000 1702.400 ;
        RECT 1400.860 52.010 1401.000 1700.000 ;
        RECT 495.980 51.690 496.240 52.010 ;
        RECT 1400.800 51.690 1401.060 52.010 ;
        RECT 496.040 15.630 496.180 51.690 ;
        RECT 490.460 15.310 490.720 15.630 ;
        RECT 495.980 15.310 496.240 15.630 ;
        RECT 490.520 2.400 490.660 15.310 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 52.260 508.230 52.320 ;
        RECT 1407.670 52.260 1407.990 52.320 ;
        RECT 507.910 52.120 1407.990 52.260 ;
        RECT 507.910 52.060 508.230 52.120 ;
        RECT 1407.670 52.060 1407.990 52.120 ;
      LAYER via ;
        RECT 507.940 52.060 508.200 52.320 ;
        RECT 1407.700 52.060 1407.960 52.320 ;
      LAYER met2 ;
        RECT 1409.920 1700.410 1410.200 1702.400 ;
        RECT 1407.760 1700.270 1410.200 1700.410 ;
        RECT 1407.760 52.350 1407.900 1700.270 ;
        RECT 1409.920 1700.000 1410.200 1700.270 ;
        RECT 507.940 52.030 508.200 52.350 ;
        RECT 1407.700 52.030 1407.960 52.350 ;
        RECT 508.000 2.400 508.140 52.030 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1415.565 1352.605 1415.735 1400.715 ;
        RECT 1415.565 1256.045 1415.735 1304.155 ;
        RECT 1415.565 774.605 1415.735 821.015 ;
        RECT 1415.565 579.785 1415.735 627.895 ;
        RECT 1415.565 483.225 1415.735 531.335 ;
        RECT 1414.645 235.025 1414.815 282.795 ;
        RECT 1414.645 138.125 1414.815 227.715 ;
      LAYER mcon ;
        RECT 1415.565 1400.545 1415.735 1400.715 ;
        RECT 1415.565 1303.985 1415.735 1304.155 ;
        RECT 1415.565 820.845 1415.735 821.015 ;
        RECT 1415.565 627.725 1415.735 627.895 ;
        RECT 1415.565 531.165 1415.735 531.335 ;
        RECT 1414.645 282.625 1414.815 282.795 ;
        RECT 1414.645 227.545 1414.815 227.715 ;
      LAYER met1 ;
        RECT 1415.030 1593.820 1415.350 1593.880 ;
        RECT 1415.490 1593.820 1415.810 1593.880 ;
        RECT 1415.030 1593.680 1415.810 1593.820 ;
        RECT 1415.030 1593.620 1415.350 1593.680 ;
        RECT 1415.490 1593.620 1415.810 1593.680 ;
        RECT 1415.030 1587.020 1415.350 1587.080 ;
        RECT 1416.410 1587.020 1416.730 1587.080 ;
        RECT 1415.030 1586.880 1416.730 1587.020 ;
        RECT 1415.030 1586.820 1415.350 1586.880 ;
        RECT 1416.410 1586.820 1416.730 1586.880 ;
        RECT 1415.490 1400.700 1415.810 1400.760 ;
        RECT 1415.295 1400.560 1415.810 1400.700 ;
        RECT 1415.490 1400.500 1415.810 1400.560 ;
        RECT 1415.490 1352.760 1415.810 1352.820 ;
        RECT 1415.295 1352.620 1415.810 1352.760 ;
        RECT 1415.490 1352.560 1415.810 1352.620 ;
        RECT 1415.490 1304.140 1415.810 1304.200 ;
        RECT 1415.295 1304.000 1415.810 1304.140 ;
        RECT 1415.490 1303.940 1415.810 1304.000 ;
        RECT 1415.490 1256.200 1415.810 1256.260 ;
        RECT 1415.295 1256.060 1415.810 1256.200 ;
        RECT 1415.490 1256.000 1415.810 1256.060 ;
        RECT 1414.570 1159.300 1414.890 1159.360 ;
        RECT 1415.490 1159.300 1415.810 1159.360 ;
        RECT 1414.570 1159.160 1415.810 1159.300 ;
        RECT 1414.570 1159.100 1414.890 1159.160 ;
        RECT 1415.490 1159.100 1415.810 1159.160 ;
        RECT 1414.570 869.620 1414.890 869.680 ;
        RECT 1415.490 869.620 1415.810 869.680 ;
        RECT 1414.570 869.480 1415.810 869.620 ;
        RECT 1414.570 869.420 1414.890 869.480 ;
        RECT 1415.490 869.420 1415.810 869.480 ;
        RECT 1415.490 821.000 1415.810 821.060 ;
        RECT 1415.295 820.860 1415.810 821.000 ;
        RECT 1415.490 820.800 1415.810 820.860 ;
        RECT 1415.490 774.760 1415.810 774.820 ;
        RECT 1415.295 774.620 1415.810 774.760 ;
        RECT 1415.490 774.560 1415.810 774.620 ;
        RECT 1415.490 627.880 1415.810 627.940 ;
        RECT 1415.295 627.740 1415.810 627.880 ;
        RECT 1415.490 627.680 1415.810 627.740 ;
        RECT 1415.490 579.940 1415.810 580.000 ;
        RECT 1415.295 579.800 1415.810 579.940 ;
        RECT 1415.490 579.740 1415.810 579.800 ;
        RECT 1415.490 531.320 1415.810 531.380 ;
        RECT 1415.295 531.180 1415.810 531.320 ;
        RECT 1415.490 531.120 1415.810 531.180 ;
        RECT 1415.490 483.380 1415.810 483.440 ;
        RECT 1415.295 483.240 1415.810 483.380 ;
        RECT 1415.490 483.180 1415.810 483.240 ;
        RECT 1414.585 282.780 1414.875 282.825 ;
        RECT 1415.490 282.780 1415.810 282.840 ;
        RECT 1414.585 282.640 1415.810 282.780 ;
        RECT 1414.585 282.595 1414.875 282.640 ;
        RECT 1415.490 282.580 1415.810 282.640 ;
        RECT 1414.570 235.180 1414.890 235.240 ;
        RECT 1414.375 235.040 1414.890 235.180 ;
        RECT 1414.570 234.980 1414.890 235.040 ;
        RECT 1414.570 234.500 1414.890 234.560 ;
        RECT 1415.490 234.500 1415.810 234.560 ;
        RECT 1414.570 234.360 1415.810 234.500 ;
        RECT 1414.570 234.300 1414.890 234.360 ;
        RECT 1415.490 234.300 1415.810 234.360 ;
        RECT 1414.585 227.700 1414.875 227.745 ;
        RECT 1415.490 227.700 1415.810 227.760 ;
        RECT 1414.585 227.560 1415.810 227.700 ;
        RECT 1414.585 227.515 1414.875 227.560 ;
        RECT 1415.490 227.500 1415.810 227.560 ;
        RECT 1414.570 138.280 1414.890 138.340 ;
        RECT 1414.375 138.140 1414.890 138.280 ;
        RECT 1414.570 138.080 1414.890 138.140 ;
        RECT 1414.570 96.800 1414.890 96.860 ;
        RECT 1415.950 96.800 1416.270 96.860 ;
        RECT 1414.570 96.660 1416.270 96.800 ;
        RECT 1414.570 96.600 1414.890 96.660 ;
        RECT 1415.950 96.600 1416.270 96.660 ;
        RECT 525.850 52.600 526.170 52.660 ;
        RECT 1415.950 52.600 1416.270 52.660 ;
        RECT 525.850 52.460 1416.270 52.600 ;
        RECT 525.850 52.400 526.170 52.460 ;
        RECT 1415.950 52.400 1416.270 52.460 ;
      LAYER via ;
        RECT 1415.060 1593.620 1415.320 1593.880 ;
        RECT 1415.520 1593.620 1415.780 1593.880 ;
        RECT 1415.060 1586.820 1415.320 1587.080 ;
        RECT 1416.440 1586.820 1416.700 1587.080 ;
        RECT 1415.520 1400.500 1415.780 1400.760 ;
        RECT 1415.520 1352.560 1415.780 1352.820 ;
        RECT 1415.520 1303.940 1415.780 1304.200 ;
        RECT 1415.520 1256.000 1415.780 1256.260 ;
        RECT 1414.600 1159.100 1414.860 1159.360 ;
        RECT 1415.520 1159.100 1415.780 1159.360 ;
        RECT 1414.600 869.420 1414.860 869.680 ;
        RECT 1415.520 869.420 1415.780 869.680 ;
        RECT 1415.520 820.800 1415.780 821.060 ;
        RECT 1415.520 774.560 1415.780 774.820 ;
        RECT 1415.520 627.680 1415.780 627.940 ;
        RECT 1415.520 579.740 1415.780 580.000 ;
        RECT 1415.520 531.120 1415.780 531.380 ;
        RECT 1415.520 483.180 1415.780 483.440 ;
        RECT 1415.520 282.580 1415.780 282.840 ;
        RECT 1414.600 234.980 1414.860 235.240 ;
        RECT 1414.600 234.300 1414.860 234.560 ;
        RECT 1415.520 234.300 1415.780 234.560 ;
        RECT 1415.520 227.500 1415.780 227.760 ;
        RECT 1414.600 138.080 1414.860 138.340 ;
        RECT 1414.600 96.600 1414.860 96.860 ;
        RECT 1415.980 96.600 1416.240 96.860 ;
        RECT 525.880 52.400 526.140 52.660 ;
        RECT 1415.980 52.400 1416.240 52.660 ;
      LAYER met2 ;
        RECT 1419.120 1701.090 1419.400 1702.400 ;
        RECT 1416.500 1700.950 1419.400 1701.090 ;
        RECT 1416.500 1677.970 1416.640 1700.950 ;
        RECT 1419.120 1700.000 1419.400 1700.950 ;
        RECT 1415.580 1677.830 1416.640 1677.970 ;
        RECT 1415.580 1593.910 1415.720 1677.830 ;
        RECT 1415.060 1593.590 1415.320 1593.910 ;
        RECT 1415.520 1593.590 1415.780 1593.910 ;
        RECT 1415.120 1587.110 1415.260 1593.590 ;
        RECT 1415.060 1586.790 1415.320 1587.110 ;
        RECT 1416.440 1586.790 1416.700 1587.110 ;
        RECT 1416.500 1462.920 1416.640 1586.790 ;
        RECT 1415.580 1462.780 1416.640 1462.920 ;
        RECT 1415.580 1400.790 1415.720 1462.780 ;
        RECT 1415.520 1400.470 1415.780 1400.790 ;
        RECT 1415.520 1352.530 1415.780 1352.850 ;
        RECT 1415.580 1304.230 1415.720 1352.530 ;
        RECT 1415.520 1303.910 1415.780 1304.230 ;
        RECT 1415.520 1255.970 1415.780 1256.290 ;
        RECT 1415.580 1207.525 1415.720 1255.970 ;
        RECT 1414.590 1207.155 1414.870 1207.525 ;
        RECT 1415.510 1207.155 1415.790 1207.525 ;
        RECT 1414.660 1159.390 1414.800 1207.155 ;
        RECT 1414.600 1159.070 1414.860 1159.390 ;
        RECT 1415.520 1159.070 1415.780 1159.390 ;
        RECT 1415.580 1076.850 1415.720 1159.070 ;
        RECT 1415.120 1076.710 1415.720 1076.850 ;
        RECT 1415.120 1076.170 1415.260 1076.710 ;
        RECT 1415.120 1076.030 1415.720 1076.170 ;
        RECT 1415.580 980.290 1415.720 1076.030 ;
        RECT 1415.120 980.150 1415.720 980.290 ;
        RECT 1415.120 979.610 1415.260 980.150 ;
        RECT 1415.120 979.470 1415.720 979.610 ;
        RECT 1415.580 917.845 1415.720 979.470 ;
        RECT 1414.590 917.475 1414.870 917.845 ;
        RECT 1415.510 917.475 1415.790 917.845 ;
        RECT 1414.660 869.710 1414.800 917.475 ;
        RECT 1414.600 869.390 1414.860 869.710 ;
        RECT 1415.520 869.390 1415.780 869.710 ;
        RECT 1415.580 821.090 1415.720 869.390 ;
        RECT 1415.520 820.770 1415.780 821.090 ;
        RECT 1415.520 774.530 1415.780 774.850 ;
        RECT 1415.580 690.610 1415.720 774.530 ;
        RECT 1415.120 690.470 1415.720 690.610 ;
        RECT 1415.120 689.250 1415.260 690.470 ;
        RECT 1415.120 689.110 1415.720 689.250 ;
        RECT 1415.580 627.970 1415.720 689.110 ;
        RECT 1415.520 627.650 1415.780 627.970 ;
        RECT 1415.520 579.710 1415.780 580.030 ;
        RECT 1415.580 531.410 1415.720 579.710 ;
        RECT 1415.520 531.090 1415.780 531.410 ;
        RECT 1415.520 483.150 1415.780 483.470 ;
        RECT 1415.580 303.690 1415.720 483.150 ;
        RECT 1415.120 303.550 1415.720 303.690 ;
        RECT 1415.120 303.010 1415.260 303.550 ;
        RECT 1415.120 302.870 1415.720 303.010 ;
        RECT 1415.580 282.870 1415.720 302.870 ;
        RECT 1415.520 282.550 1415.780 282.870 ;
        RECT 1414.600 234.950 1414.860 235.270 ;
        RECT 1414.660 234.590 1414.800 234.950 ;
        RECT 1414.600 234.270 1414.860 234.590 ;
        RECT 1415.520 234.270 1415.780 234.590 ;
        RECT 1415.580 227.790 1415.720 234.270 ;
        RECT 1415.520 227.470 1415.780 227.790 ;
        RECT 1414.600 138.050 1414.860 138.370 ;
        RECT 1414.660 96.890 1414.800 138.050 ;
        RECT 1414.600 96.570 1414.860 96.890 ;
        RECT 1415.980 96.570 1416.240 96.890 ;
        RECT 1416.040 52.690 1416.180 96.570 ;
        RECT 525.880 52.370 526.140 52.690 ;
        RECT 1415.980 52.370 1416.240 52.690 ;
        RECT 525.940 2.400 526.080 52.370 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 1414.590 1207.200 1414.870 1207.480 ;
        RECT 1415.510 1207.200 1415.790 1207.480 ;
        RECT 1414.590 917.520 1414.870 917.800 ;
        RECT 1415.510 917.520 1415.790 917.800 ;
      LAYER met3 ;
        RECT 1414.565 1207.490 1414.895 1207.505 ;
        RECT 1415.485 1207.490 1415.815 1207.505 ;
        RECT 1414.565 1207.190 1415.815 1207.490 ;
        RECT 1414.565 1207.175 1414.895 1207.190 ;
        RECT 1415.485 1207.175 1415.815 1207.190 ;
        RECT 1414.565 917.810 1414.895 917.825 ;
        RECT 1415.485 917.810 1415.815 917.825 ;
        RECT 1414.565 917.510 1415.815 917.810 ;
        RECT 1414.565 917.495 1414.895 917.510 ;
        RECT 1415.485 917.495 1415.815 917.510 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 52.940 544.110 53.000 ;
        RECT 1428.370 52.940 1428.690 53.000 ;
        RECT 543.790 52.800 1428.690 52.940 ;
        RECT 543.790 52.740 544.110 52.800 ;
        RECT 1428.370 52.740 1428.690 52.800 ;
      LAYER via ;
        RECT 543.820 52.740 544.080 53.000 ;
        RECT 1428.400 52.740 1428.660 53.000 ;
      LAYER met2 ;
        RECT 1428.320 1700.000 1428.600 1702.400 ;
        RECT 1428.460 53.030 1428.600 1700.000 ;
        RECT 543.820 52.710 544.080 53.030 ;
        RECT 1428.400 52.710 1428.660 53.030 ;
        RECT 543.880 2.400 544.020 52.710 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 53.280 565.730 53.340 ;
        RECT 1435.270 53.280 1435.590 53.340 ;
        RECT 565.410 53.140 1435.590 53.280 ;
        RECT 565.410 53.080 565.730 53.140 ;
        RECT 1435.270 53.080 1435.590 53.140 ;
        RECT 561.730 14.860 562.050 14.920 ;
        RECT 565.410 14.860 565.730 14.920 ;
        RECT 561.730 14.720 565.730 14.860 ;
        RECT 561.730 14.660 562.050 14.720 ;
        RECT 565.410 14.660 565.730 14.720 ;
      LAYER via ;
        RECT 565.440 53.080 565.700 53.340 ;
        RECT 1435.300 53.080 1435.560 53.340 ;
        RECT 561.760 14.660 562.020 14.920 ;
        RECT 565.440 14.660 565.700 14.920 ;
      LAYER met2 ;
        RECT 1437.520 1700.410 1437.800 1702.400 ;
        RECT 1435.360 1700.270 1437.800 1700.410 ;
        RECT 1435.360 53.370 1435.500 1700.270 ;
        RECT 1437.520 1700.000 1437.800 1700.270 ;
        RECT 565.440 53.050 565.700 53.370 ;
        RECT 1435.300 53.050 1435.560 53.370 ;
        RECT 565.500 14.950 565.640 53.050 ;
        RECT 561.760 14.630 562.020 14.950 ;
        RECT 565.440 14.630 565.700 14.950 ;
        RECT 561.820 2.400 561.960 14.630 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1443.165 1545.725 1443.335 1593.835 ;
        RECT 1443.165 774.605 1443.335 821.015 ;
        RECT 1442.705 241.485 1442.875 289.595 ;
      LAYER mcon ;
        RECT 1443.165 1593.665 1443.335 1593.835 ;
        RECT 1443.165 820.845 1443.335 821.015 ;
        RECT 1442.705 289.425 1442.875 289.595 ;
      LAYER met1 ;
        RECT 1443.090 1593.820 1443.410 1593.880 ;
        RECT 1442.895 1593.680 1443.410 1593.820 ;
        RECT 1443.090 1593.620 1443.410 1593.680 ;
        RECT 1443.090 1545.880 1443.410 1545.940 ;
        RECT 1442.895 1545.740 1443.410 1545.880 ;
        RECT 1443.090 1545.680 1443.410 1545.740 ;
        RECT 1443.090 1462.380 1443.410 1462.640 ;
        RECT 1443.180 1461.960 1443.320 1462.380 ;
        RECT 1443.090 1461.700 1443.410 1461.960 ;
        RECT 1443.090 1365.820 1443.410 1366.080 ;
        RECT 1443.180 1365.400 1443.320 1365.820 ;
        RECT 1443.090 1365.140 1443.410 1365.400 ;
        RECT 1443.090 1269.260 1443.410 1269.520 ;
        RECT 1443.180 1268.840 1443.320 1269.260 ;
        RECT 1443.090 1268.580 1443.410 1268.840 ;
        RECT 1443.090 1172.700 1443.410 1172.960 ;
        RECT 1443.180 1172.280 1443.320 1172.700 ;
        RECT 1443.090 1172.020 1443.410 1172.280 ;
        RECT 1443.090 883.020 1443.410 883.280 ;
        RECT 1443.180 882.600 1443.320 883.020 ;
        RECT 1443.090 882.340 1443.410 882.600 ;
        RECT 1443.090 821.000 1443.410 821.060 ;
        RECT 1442.895 820.860 1443.410 821.000 ;
        RECT 1443.090 820.800 1443.410 820.860 ;
        RECT 1443.090 774.760 1443.410 774.820 ;
        RECT 1442.895 774.620 1443.410 774.760 ;
        RECT 1443.090 774.560 1443.410 774.620 ;
        RECT 1442.645 289.580 1442.935 289.625 ;
        RECT 1443.090 289.580 1443.410 289.640 ;
        RECT 1442.645 289.440 1443.410 289.580 ;
        RECT 1442.645 289.395 1442.935 289.440 ;
        RECT 1443.090 289.380 1443.410 289.440 ;
        RECT 1442.630 241.640 1442.950 241.700 ;
        RECT 1442.435 241.500 1442.950 241.640 ;
        RECT 1442.630 241.440 1442.950 241.500 ;
        RECT 1442.170 96.800 1442.490 96.860 ;
        RECT 1443.090 96.800 1443.410 96.860 ;
        RECT 1442.170 96.660 1443.410 96.800 ;
        RECT 1442.170 96.600 1442.490 96.660 ;
        RECT 1443.090 96.600 1443.410 96.660 ;
        RECT 585.650 53.620 585.970 53.680 ;
        RECT 1441.710 53.620 1442.030 53.680 ;
        RECT 585.650 53.480 1442.030 53.620 ;
        RECT 585.650 53.420 585.970 53.480 ;
        RECT 1441.710 53.420 1442.030 53.480 ;
        RECT 579.670 14.860 579.990 14.920 ;
        RECT 584.730 14.860 585.050 14.920 ;
        RECT 579.670 14.720 585.050 14.860 ;
        RECT 579.670 14.660 579.990 14.720 ;
        RECT 584.730 14.660 585.050 14.720 ;
      LAYER via ;
        RECT 1443.120 1593.620 1443.380 1593.880 ;
        RECT 1443.120 1545.680 1443.380 1545.940 ;
        RECT 1443.120 1462.380 1443.380 1462.640 ;
        RECT 1443.120 1461.700 1443.380 1461.960 ;
        RECT 1443.120 1365.820 1443.380 1366.080 ;
        RECT 1443.120 1365.140 1443.380 1365.400 ;
        RECT 1443.120 1269.260 1443.380 1269.520 ;
        RECT 1443.120 1268.580 1443.380 1268.840 ;
        RECT 1443.120 1172.700 1443.380 1172.960 ;
        RECT 1443.120 1172.020 1443.380 1172.280 ;
        RECT 1443.120 883.020 1443.380 883.280 ;
        RECT 1443.120 882.340 1443.380 882.600 ;
        RECT 1443.120 820.800 1443.380 821.060 ;
        RECT 1443.120 774.560 1443.380 774.820 ;
        RECT 1443.120 289.380 1443.380 289.640 ;
        RECT 1442.660 241.440 1442.920 241.700 ;
        RECT 1442.200 96.600 1442.460 96.860 ;
        RECT 1443.120 96.600 1443.380 96.860 ;
        RECT 585.680 53.420 585.940 53.680 ;
        RECT 1441.740 53.420 1442.000 53.680 ;
        RECT 579.700 14.660 579.960 14.920 ;
        RECT 584.760 14.660 585.020 14.920 ;
      LAYER met2 ;
        RECT 1446.720 1701.090 1447.000 1702.400 ;
        RECT 1444.100 1700.950 1447.000 1701.090 ;
        RECT 1444.100 1656.210 1444.240 1700.950 ;
        RECT 1446.720 1700.000 1447.000 1700.950 ;
        RECT 1442.720 1656.070 1444.240 1656.210 ;
        RECT 1442.720 1606.570 1442.860 1656.070 ;
        RECT 1442.720 1606.430 1443.320 1606.570 ;
        RECT 1443.180 1593.910 1443.320 1606.430 ;
        RECT 1443.120 1593.590 1443.380 1593.910 ;
        RECT 1443.120 1545.650 1443.380 1545.970 ;
        RECT 1443.180 1462.670 1443.320 1545.650 ;
        RECT 1443.120 1462.350 1443.380 1462.670 ;
        RECT 1443.120 1461.670 1443.380 1461.990 ;
        RECT 1443.180 1366.110 1443.320 1461.670 ;
        RECT 1443.120 1365.790 1443.380 1366.110 ;
        RECT 1443.120 1365.110 1443.380 1365.430 ;
        RECT 1443.180 1269.550 1443.320 1365.110 ;
        RECT 1443.120 1269.230 1443.380 1269.550 ;
        RECT 1443.120 1268.550 1443.380 1268.870 ;
        RECT 1443.180 1172.990 1443.320 1268.550 ;
        RECT 1443.120 1172.670 1443.380 1172.990 ;
        RECT 1443.120 1171.990 1443.380 1172.310 ;
        RECT 1443.180 1076.850 1443.320 1171.990 ;
        RECT 1442.720 1076.710 1443.320 1076.850 ;
        RECT 1442.720 1076.170 1442.860 1076.710 ;
        RECT 1442.720 1076.030 1443.320 1076.170 ;
        RECT 1443.180 980.290 1443.320 1076.030 ;
        RECT 1442.720 980.150 1443.320 980.290 ;
        RECT 1442.720 979.610 1442.860 980.150 ;
        RECT 1442.720 979.470 1443.320 979.610 ;
        RECT 1443.180 883.310 1443.320 979.470 ;
        RECT 1443.120 882.990 1443.380 883.310 ;
        RECT 1443.120 882.310 1443.380 882.630 ;
        RECT 1443.180 821.090 1443.320 882.310 ;
        RECT 1443.120 820.770 1443.380 821.090 ;
        RECT 1443.120 774.530 1443.380 774.850 ;
        RECT 1443.180 690.610 1443.320 774.530 ;
        RECT 1442.720 690.470 1443.320 690.610 ;
        RECT 1442.720 689.250 1442.860 690.470 ;
        RECT 1442.720 689.110 1443.320 689.250 ;
        RECT 1443.180 303.690 1443.320 689.110 ;
        RECT 1442.720 303.550 1443.320 303.690 ;
        RECT 1442.720 303.010 1442.860 303.550 ;
        RECT 1442.720 302.870 1443.320 303.010 ;
        RECT 1443.180 289.670 1443.320 302.870 ;
        RECT 1443.120 289.350 1443.380 289.670 ;
        RECT 1442.660 241.410 1442.920 241.730 ;
        RECT 1442.720 241.130 1442.860 241.410 ;
        RECT 1442.720 240.990 1443.320 241.130 ;
        RECT 1443.180 96.890 1443.320 240.990 ;
        RECT 1442.200 96.570 1442.460 96.890 ;
        RECT 1443.120 96.570 1443.380 96.890 ;
        RECT 1442.260 62.970 1442.400 96.570 ;
        RECT 1441.800 62.830 1442.400 62.970 ;
        RECT 1441.800 53.710 1441.940 62.830 ;
        RECT 585.680 53.390 585.940 53.710 ;
        RECT 1441.740 53.390 1442.000 53.710 ;
        RECT 585.740 18.090 585.880 53.390 ;
        RECT 584.820 17.950 585.880 18.090 ;
        RECT 584.820 14.950 584.960 17.950 ;
        RECT 579.700 14.630 579.960 14.950 ;
        RECT 584.760 14.630 585.020 14.950 ;
        RECT 579.760 2.400 579.900 14.630 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1187.330 1668.280 1187.650 1668.340 ;
        RECT 1191.470 1668.280 1191.790 1668.340 ;
        RECT 1187.330 1668.140 1191.790 1668.280 ;
        RECT 1187.330 1668.080 1187.650 1668.140 ;
        RECT 1191.470 1668.080 1191.790 1668.140 ;
        RECT 86.550 25.740 86.870 25.800 ;
        RECT 1187.330 25.740 1187.650 25.800 ;
        RECT 86.550 25.600 1187.650 25.740 ;
        RECT 86.550 25.540 86.870 25.600 ;
        RECT 1187.330 25.540 1187.650 25.600 ;
      LAYER via ;
        RECT 1187.360 1668.080 1187.620 1668.340 ;
        RECT 1191.500 1668.080 1191.760 1668.340 ;
        RECT 86.580 25.540 86.840 25.800 ;
        RECT 1187.360 25.540 1187.620 25.800 ;
      LAYER met2 ;
        RECT 1192.800 1700.410 1193.080 1702.400 ;
        RECT 1191.560 1700.270 1193.080 1700.410 ;
        RECT 1191.560 1668.370 1191.700 1700.270 ;
        RECT 1192.800 1700.000 1193.080 1700.270 ;
        RECT 1187.360 1668.050 1187.620 1668.370 ;
        RECT 1191.500 1668.050 1191.760 1668.370 ;
        RECT 1187.420 25.830 1187.560 1668.050 ;
        RECT 86.580 25.510 86.840 25.830 ;
        RECT 1187.360 25.510 1187.620 25.830 ;
        RECT 86.640 5.170 86.780 25.510 ;
        RECT 86.180 5.030 86.780 5.170 ;
        RECT 86.180 2.400 86.320 5.030 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 53.960 600.230 54.020 ;
        RECT 1455.970 53.960 1456.290 54.020 ;
        RECT 599.910 53.820 1456.290 53.960 ;
        RECT 599.910 53.760 600.230 53.820 ;
        RECT 1455.970 53.760 1456.290 53.820 ;
        RECT 597.150 14.860 597.470 14.920 ;
        RECT 599.910 14.860 600.230 14.920 ;
        RECT 597.150 14.720 600.230 14.860 ;
        RECT 597.150 14.660 597.470 14.720 ;
        RECT 599.910 14.660 600.230 14.720 ;
      LAYER via ;
        RECT 599.940 53.760 600.200 54.020 ;
        RECT 1456.000 53.760 1456.260 54.020 ;
        RECT 597.180 14.660 597.440 14.920 ;
        RECT 599.940 14.660 600.200 14.920 ;
      LAYER met2 ;
        RECT 1455.920 1700.000 1456.200 1702.400 ;
        RECT 1456.060 54.050 1456.200 1700.000 ;
        RECT 599.940 53.730 600.200 54.050 ;
        RECT 1456.000 53.730 1456.260 54.050 ;
        RECT 600.000 14.950 600.140 53.730 ;
        RECT 597.180 14.630 597.440 14.950 ;
        RECT 599.940 14.630 600.200 14.950 ;
        RECT 597.240 2.400 597.380 14.630 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 54.300 620.930 54.360 ;
        RECT 1462.870 54.300 1463.190 54.360 ;
        RECT 620.610 54.160 1463.190 54.300 ;
        RECT 620.610 54.100 620.930 54.160 ;
        RECT 1462.870 54.100 1463.190 54.160 ;
      LAYER via ;
        RECT 620.640 54.100 620.900 54.360 ;
        RECT 1462.900 54.100 1463.160 54.360 ;
      LAYER met2 ;
        RECT 1465.120 1700.410 1465.400 1702.400 ;
        RECT 1462.960 1700.270 1465.400 1700.410 ;
        RECT 1462.960 54.390 1463.100 1700.270 ;
        RECT 1465.120 1700.000 1465.400 1700.270 ;
        RECT 620.640 54.070 620.900 54.390 ;
        RECT 1462.900 54.070 1463.160 54.390 ;
        RECT 620.700 17.410 620.840 54.070 ;
        RECT 615.180 17.270 620.840 17.410 ;
        RECT 615.180 2.400 615.320 17.270 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1200.745 662.405 1200.915 710.515 ;
      LAYER mcon ;
        RECT 1200.745 710.345 1200.915 710.515 ;
      LAYER met1 ;
        RECT 1200.670 821.000 1200.990 821.060 ;
        RECT 1201.590 821.000 1201.910 821.060 ;
        RECT 1200.670 820.860 1201.910 821.000 ;
        RECT 1200.670 820.800 1200.990 820.860 ;
        RECT 1201.590 820.800 1201.910 820.860 ;
        RECT 1200.670 765.920 1200.990 765.980 ;
        RECT 1201.130 765.920 1201.450 765.980 ;
        RECT 1200.670 765.780 1201.450 765.920 ;
        RECT 1200.670 765.720 1200.990 765.780 ;
        RECT 1201.130 765.720 1201.450 765.780 ;
        RECT 1200.670 710.500 1200.990 710.560 ;
        RECT 1200.475 710.360 1200.990 710.500 ;
        RECT 1200.670 710.300 1200.990 710.360 ;
        RECT 1200.685 662.560 1200.975 662.605 ;
        RECT 1201.590 662.560 1201.910 662.620 ;
        RECT 1200.685 662.420 1201.910 662.560 ;
        RECT 1200.685 662.375 1200.975 662.420 ;
        RECT 1201.590 662.360 1201.910 662.420 ;
        RECT 1201.130 352.280 1201.450 352.540 ;
        RECT 1201.220 351.860 1201.360 352.280 ;
        RECT 1201.130 351.600 1201.450 351.860 ;
        RECT 109.550 26.080 109.870 26.140 ;
        RECT 1201.130 26.080 1201.450 26.140 ;
        RECT 109.550 25.940 1201.450 26.080 ;
        RECT 109.550 25.880 109.870 25.940 ;
        RECT 1201.130 25.880 1201.450 25.940 ;
      LAYER via ;
        RECT 1200.700 820.800 1200.960 821.060 ;
        RECT 1201.620 820.800 1201.880 821.060 ;
        RECT 1200.700 765.720 1200.960 765.980 ;
        RECT 1201.160 765.720 1201.420 765.980 ;
        RECT 1200.700 710.300 1200.960 710.560 ;
        RECT 1201.620 662.360 1201.880 662.620 ;
        RECT 1201.160 352.280 1201.420 352.540 ;
        RECT 1201.160 351.600 1201.420 351.860 ;
        RECT 109.580 25.880 109.840 26.140 ;
        RECT 1201.160 25.880 1201.420 26.140 ;
      LAYER met2 ;
        RECT 1204.760 1700.410 1205.040 1702.400 ;
        RECT 1203.060 1700.270 1205.040 1700.410 ;
        RECT 1203.060 1656.210 1203.200 1700.270 ;
        RECT 1204.760 1700.000 1205.040 1700.270 ;
        RECT 1200.760 1656.070 1203.200 1656.210 ;
        RECT 1200.760 1655.530 1200.900 1656.070 ;
        RECT 1200.760 1655.390 1201.360 1655.530 ;
        RECT 1201.220 1511.370 1201.360 1655.390 ;
        RECT 1200.760 1511.230 1201.360 1511.370 ;
        RECT 1200.760 1510.690 1200.900 1511.230 ;
        RECT 1200.760 1510.550 1201.360 1510.690 ;
        RECT 1201.220 1414.810 1201.360 1510.550 ;
        RECT 1200.760 1414.670 1201.360 1414.810 ;
        RECT 1200.760 1414.130 1200.900 1414.670 ;
        RECT 1200.760 1413.990 1201.360 1414.130 ;
        RECT 1201.220 1318.250 1201.360 1413.990 ;
        RECT 1200.760 1318.110 1201.360 1318.250 ;
        RECT 1200.760 1317.570 1200.900 1318.110 ;
        RECT 1200.760 1317.430 1201.360 1317.570 ;
        RECT 1201.220 1221.690 1201.360 1317.430 ;
        RECT 1200.760 1221.550 1201.360 1221.690 ;
        RECT 1200.760 1221.010 1200.900 1221.550 ;
        RECT 1200.760 1220.870 1201.360 1221.010 ;
        RECT 1201.220 1125.130 1201.360 1220.870 ;
        RECT 1200.760 1124.990 1201.360 1125.130 ;
        RECT 1200.760 1124.450 1200.900 1124.990 ;
        RECT 1200.760 1124.310 1201.360 1124.450 ;
        RECT 1201.220 1028.570 1201.360 1124.310 ;
        RECT 1200.760 1028.430 1201.360 1028.570 ;
        RECT 1200.760 1027.890 1200.900 1028.430 ;
        RECT 1200.760 1027.750 1201.360 1027.890 ;
        RECT 1201.220 932.010 1201.360 1027.750 ;
        RECT 1200.760 931.870 1201.360 932.010 ;
        RECT 1200.760 931.330 1200.900 931.870 ;
        RECT 1200.760 931.190 1201.360 931.330 ;
        RECT 1201.220 835.450 1201.360 931.190 ;
        RECT 1201.220 835.310 1201.820 835.450 ;
        RECT 1201.680 821.285 1201.820 835.310 ;
        RECT 1200.690 820.915 1200.970 821.285 ;
        RECT 1201.610 820.915 1201.890 821.285 ;
        RECT 1200.700 820.770 1200.960 820.915 ;
        RECT 1201.620 820.770 1201.880 820.915 ;
        RECT 1201.680 796.010 1201.820 820.770 ;
        RECT 1201.220 795.870 1201.820 796.010 ;
        RECT 1201.220 766.010 1201.360 795.870 ;
        RECT 1200.700 765.690 1200.960 766.010 ;
        RECT 1201.160 765.690 1201.420 766.010 ;
        RECT 1200.760 718.605 1200.900 765.690 ;
        RECT 1200.690 718.235 1200.970 718.605 ;
        RECT 1200.690 717.555 1200.970 717.925 ;
        RECT 1200.760 710.590 1200.900 717.555 ;
        RECT 1200.700 710.270 1200.960 710.590 ;
        RECT 1201.620 662.330 1201.880 662.650 ;
        RECT 1201.680 640.970 1201.820 662.330 ;
        RECT 1200.760 640.830 1201.820 640.970 ;
        RECT 1200.760 596.770 1200.900 640.830 ;
        RECT 1200.760 596.630 1201.360 596.770 ;
        RECT 1201.220 449.210 1201.360 596.630 ;
        RECT 1200.760 449.070 1201.360 449.210 ;
        RECT 1200.760 448.530 1200.900 449.070 ;
        RECT 1200.760 448.390 1201.360 448.530 ;
        RECT 1201.220 352.570 1201.360 448.390 ;
        RECT 1201.160 352.250 1201.420 352.570 ;
        RECT 1201.160 351.570 1201.420 351.890 ;
        RECT 1201.220 26.170 1201.360 351.570 ;
        RECT 109.580 25.850 109.840 26.170 ;
        RECT 1201.160 25.850 1201.420 26.170 ;
        RECT 109.640 2.400 109.780 25.850 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 1200.690 820.960 1200.970 821.240 ;
        RECT 1201.610 820.960 1201.890 821.240 ;
        RECT 1200.690 718.280 1200.970 718.560 ;
        RECT 1200.690 717.600 1200.970 717.880 ;
      LAYER met3 ;
        RECT 1200.665 821.250 1200.995 821.265 ;
        RECT 1201.585 821.250 1201.915 821.265 ;
        RECT 1200.665 820.950 1201.915 821.250 ;
        RECT 1200.665 820.935 1200.995 820.950 ;
        RECT 1201.585 820.935 1201.915 820.950 ;
        RECT 1200.665 718.570 1200.995 718.585 ;
        RECT 1200.665 718.255 1201.210 718.570 ;
        RECT 1200.910 717.905 1201.210 718.255 ;
        RECT 1200.665 717.590 1201.210 717.905 ;
        RECT 1200.665 717.575 1200.995 717.590 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 38.660 133.790 38.720 ;
        RECT 1214.470 38.660 1214.790 38.720 ;
        RECT 133.470 38.520 1214.790 38.660 ;
        RECT 133.470 38.460 133.790 38.520 ;
        RECT 1214.470 38.460 1214.790 38.520 ;
      LAYER via ;
        RECT 133.500 38.460 133.760 38.720 ;
        RECT 1214.500 38.460 1214.760 38.720 ;
      LAYER met2 ;
        RECT 1217.180 1700.410 1217.460 1702.400 ;
        RECT 1214.560 1700.270 1217.460 1700.410 ;
        RECT 1214.560 38.750 1214.700 1700.270 ;
        RECT 1217.180 1700.000 1217.460 1700.270 ;
        RECT 133.500 38.430 133.760 38.750 ;
        RECT 1214.500 38.430 1214.760 38.750 ;
        RECT 133.560 2.400 133.700 38.430 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1221.905 234.685 1222.075 282.795 ;
      LAYER mcon ;
        RECT 1221.905 282.625 1222.075 282.795 ;
      LAYER met1 ;
        RECT 1222.290 1400.700 1222.610 1400.760 ;
        RECT 1222.750 1400.700 1223.070 1400.760 ;
        RECT 1222.290 1400.560 1223.070 1400.700 ;
        RECT 1222.290 1400.500 1222.610 1400.560 ;
        RECT 1222.750 1400.500 1223.070 1400.560 ;
        RECT 1222.290 1303.940 1222.610 1304.200 ;
        RECT 1222.380 1303.800 1222.520 1303.940 ;
        RECT 1222.750 1303.800 1223.070 1303.860 ;
        RECT 1222.380 1303.660 1223.070 1303.800 ;
        RECT 1222.750 1303.600 1223.070 1303.660 ;
        RECT 1222.290 934.900 1222.610 934.960 ;
        RECT 1223.210 934.900 1223.530 934.960 ;
        RECT 1222.290 934.760 1223.530 934.900 ;
        RECT 1222.290 934.700 1222.610 934.760 ;
        RECT 1223.210 934.700 1223.530 934.760 ;
        RECT 1222.290 689.900 1222.610 690.160 ;
        RECT 1222.380 689.480 1222.520 689.900 ;
        RECT 1222.290 689.220 1222.610 689.480 ;
        RECT 1222.290 400.220 1222.610 400.480 ;
        RECT 1222.380 399.800 1222.520 400.220 ;
        RECT 1222.290 399.540 1222.610 399.800 ;
        RECT 1221.845 282.780 1222.135 282.825 ;
        RECT 1222.290 282.780 1222.610 282.840 ;
        RECT 1221.845 282.640 1222.610 282.780 ;
        RECT 1221.845 282.595 1222.135 282.640 ;
        RECT 1222.290 282.580 1222.610 282.640 ;
        RECT 1221.830 234.840 1222.150 234.900 ;
        RECT 1221.635 234.700 1222.150 234.840 ;
        RECT 1221.830 234.640 1222.150 234.700 ;
        RECT 1222.290 144.740 1222.610 144.800 ;
        RECT 1222.750 144.740 1223.070 144.800 ;
        RECT 1222.290 144.600 1223.070 144.740 ;
        RECT 1222.290 144.540 1222.610 144.600 ;
        RECT 1222.750 144.540 1223.070 144.600 ;
        RECT 1221.370 48.520 1221.690 48.580 ;
        RECT 1222.750 48.520 1223.070 48.580 ;
        RECT 1221.370 48.380 1223.070 48.520 ;
        RECT 1221.370 48.320 1221.690 48.380 ;
        RECT 1222.750 48.320 1223.070 48.380 ;
        RECT 151.410 39.000 151.730 39.060 ;
        RECT 1221.370 39.000 1221.690 39.060 ;
        RECT 151.410 38.860 1221.690 39.000 ;
        RECT 151.410 38.800 151.730 38.860 ;
        RECT 1221.370 38.800 1221.690 38.860 ;
      LAYER via ;
        RECT 1222.320 1400.500 1222.580 1400.760 ;
        RECT 1222.780 1400.500 1223.040 1400.760 ;
        RECT 1222.320 1303.940 1222.580 1304.200 ;
        RECT 1222.780 1303.600 1223.040 1303.860 ;
        RECT 1222.320 934.700 1222.580 934.960 ;
        RECT 1223.240 934.700 1223.500 934.960 ;
        RECT 1222.320 689.900 1222.580 690.160 ;
        RECT 1222.320 689.220 1222.580 689.480 ;
        RECT 1222.320 400.220 1222.580 400.480 ;
        RECT 1222.320 399.540 1222.580 399.800 ;
        RECT 1222.320 282.580 1222.580 282.840 ;
        RECT 1221.860 234.640 1222.120 234.900 ;
        RECT 1222.320 144.540 1222.580 144.800 ;
        RECT 1222.780 144.540 1223.040 144.800 ;
        RECT 1221.400 48.320 1221.660 48.580 ;
        RECT 1222.780 48.320 1223.040 48.580 ;
        RECT 151.440 38.800 151.700 39.060 ;
        RECT 1221.400 38.800 1221.660 39.060 ;
      LAYER met2 ;
        RECT 1226.380 1700.410 1226.660 1702.400 ;
        RECT 1224.220 1700.270 1226.660 1700.410 ;
        RECT 1224.220 1656.210 1224.360 1700.270 ;
        RECT 1226.380 1700.000 1226.660 1700.270 ;
        RECT 1222.380 1656.070 1224.360 1656.210 ;
        RECT 1222.380 1559.650 1222.520 1656.070 ;
        RECT 1221.920 1559.510 1222.520 1559.650 ;
        RECT 1221.920 1558.970 1222.060 1559.510 ;
        RECT 1221.920 1558.830 1222.520 1558.970 ;
        RECT 1222.380 1400.790 1222.520 1558.830 ;
        RECT 1222.320 1400.470 1222.580 1400.790 ;
        RECT 1222.780 1400.470 1223.040 1400.790 ;
        RECT 1222.840 1365.850 1222.980 1400.470 ;
        RECT 1222.380 1365.710 1222.980 1365.850 ;
        RECT 1222.380 1304.230 1222.520 1365.710 ;
        RECT 1222.320 1303.910 1222.580 1304.230 ;
        RECT 1222.780 1303.570 1223.040 1303.890 ;
        RECT 1222.840 1269.290 1222.980 1303.570 ;
        RECT 1222.380 1269.150 1222.980 1269.290 ;
        RECT 1222.380 980.290 1222.520 1269.150 ;
        RECT 1221.920 980.150 1222.520 980.290 ;
        RECT 1221.920 979.610 1222.060 980.150 ;
        RECT 1221.920 979.470 1222.520 979.610 ;
        RECT 1222.380 934.990 1222.520 979.470 ;
        RECT 1222.320 934.670 1222.580 934.990 ;
        RECT 1223.240 934.670 1223.500 934.990 ;
        RECT 1223.300 911.045 1223.440 934.670 ;
        RECT 1222.310 910.675 1222.590 911.045 ;
        RECT 1223.230 910.675 1223.510 911.045 ;
        RECT 1222.380 787.170 1222.520 910.675 ;
        RECT 1221.920 787.030 1222.520 787.170 ;
        RECT 1221.920 786.490 1222.060 787.030 ;
        RECT 1221.920 786.350 1222.520 786.490 ;
        RECT 1222.380 690.190 1222.520 786.350 ;
        RECT 1222.320 689.870 1222.580 690.190 ;
        RECT 1222.320 689.190 1222.580 689.510 ;
        RECT 1222.380 400.510 1222.520 689.190 ;
        RECT 1222.320 400.190 1222.580 400.510 ;
        RECT 1222.320 399.510 1222.580 399.830 ;
        RECT 1222.380 303.690 1222.520 399.510 ;
        RECT 1221.920 303.550 1222.520 303.690 ;
        RECT 1221.920 303.010 1222.060 303.550 ;
        RECT 1221.920 302.870 1222.520 303.010 ;
        RECT 1222.380 282.870 1222.520 302.870 ;
        RECT 1222.320 282.550 1222.580 282.870 ;
        RECT 1221.860 234.610 1222.120 234.930 ;
        RECT 1221.920 210.530 1222.060 234.610 ;
        RECT 1221.920 210.390 1222.520 210.530 ;
        RECT 1222.380 144.830 1222.520 210.390 ;
        RECT 1222.320 144.510 1222.580 144.830 ;
        RECT 1222.780 144.510 1223.040 144.830 ;
        RECT 1222.840 48.610 1222.980 144.510 ;
        RECT 1221.400 48.290 1221.660 48.610 ;
        RECT 1222.780 48.290 1223.040 48.610 ;
        RECT 1221.460 39.090 1221.600 48.290 ;
        RECT 151.440 38.770 151.700 39.090 ;
        RECT 1221.400 38.770 1221.660 39.090 ;
        RECT 151.500 2.400 151.640 38.770 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 1222.310 910.720 1222.590 911.000 ;
        RECT 1223.230 910.720 1223.510 911.000 ;
      LAYER met3 ;
        RECT 1222.285 911.010 1222.615 911.025 ;
        RECT 1223.205 911.010 1223.535 911.025 ;
        RECT 1222.285 910.710 1223.535 911.010 ;
        RECT 1222.285 910.695 1222.615 910.710 ;
        RECT 1223.205 910.695 1223.535 910.710 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 39.340 169.670 39.400 ;
        RECT 1236.090 39.340 1236.410 39.400 ;
        RECT 169.350 39.200 1236.410 39.340 ;
        RECT 169.350 39.140 169.670 39.200 ;
        RECT 1236.090 39.140 1236.410 39.200 ;
      LAYER via ;
        RECT 169.380 39.140 169.640 39.400 ;
        RECT 1236.120 39.140 1236.380 39.400 ;
      LAYER met2 ;
        RECT 1235.580 1700.410 1235.860 1702.400 ;
        RECT 1235.580 1700.270 1236.320 1700.410 ;
        RECT 1235.580 1700.000 1235.860 1700.270 ;
        RECT 1236.180 39.430 1236.320 1700.270 ;
        RECT 169.380 39.110 169.640 39.430 ;
        RECT 1236.120 39.110 1236.380 39.430 ;
        RECT 169.440 2.400 169.580 39.110 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 39.680 187.150 39.740 ;
        RECT 1242.530 39.680 1242.850 39.740 ;
        RECT 186.830 39.540 1242.850 39.680 ;
        RECT 186.830 39.480 187.150 39.540 ;
        RECT 1242.530 39.480 1242.850 39.540 ;
      LAYER via ;
        RECT 186.860 39.480 187.120 39.740 ;
        RECT 1242.560 39.480 1242.820 39.740 ;
      LAYER met2 ;
        RECT 1244.780 1700.410 1245.060 1702.400 ;
        RECT 1242.620 1700.270 1245.060 1700.410 ;
        RECT 1242.620 39.770 1242.760 1700.270 ;
        RECT 1244.780 1700.000 1245.060 1700.270 ;
        RECT 186.860 39.450 187.120 39.770 ;
        RECT 1242.560 39.450 1242.820 39.770 ;
        RECT 186.920 2.400 187.060 39.450 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1249.965 1587.205 1250.135 1608.455 ;
        RECT 1249.505 1442.025 1249.675 1490.475 ;
        RECT 1249.505 1393.745 1249.675 1429.275 ;
        RECT 1249.965 234.685 1250.135 282.795 ;
      LAYER mcon ;
        RECT 1249.965 1608.285 1250.135 1608.455 ;
        RECT 1249.505 1490.305 1249.675 1490.475 ;
        RECT 1249.505 1429.105 1249.675 1429.275 ;
        RECT 1249.965 282.625 1250.135 282.795 ;
      LAYER met1 ;
        RECT 1249.890 1688.680 1250.210 1688.740 ;
        RECT 1254.030 1688.680 1254.350 1688.740 ;
        RECT 1249.890 1688.540 1254.350 1688.680 ;
        RECT 1249.890 1688.480 1250.210 1688.540 ;
        RECT 1254.030 1688.480 1254.350 1688.540 ;
        RECT 1249.890 1608.440 1250.210 1608.500 ;
        RECT 1249.695 1608.300 1250.210 1608.440 ;
        RECT 1249.890 1608.240 1250.210 1608.300 ;
        RECT 1249.890 1587.360 1250.210 1587.420 ;
        RECT 1249.695 1587.220 1250.210 1587.360 ;
        RECT 1249.890 1587.160 1250.210 1587.220 ;
        RECT 1249.890 1559.480 1250.210 1559.540 ;
        RECT 1249.520 1559.340 1250.210 1559.480 ;
        RECT 1249.520 1559.200 1249.660 1559.340 ;
        RECT 1249.890 1559.280 1250.210 1559.340 ;
        RECT 1249.430 1558.940 1249.750 1559.200 ;
        RECT 1249.430 1490.460 1249.750 1490.520 ;
        RECT 1249.235 1490.320 1249.750 1490.460 ;
        RECT 1249.430 1490.260 1249.750 1490.320 ;
        RECT 1249.430 1442.180 1249.750 1442.240 ;
        RECT 1249.235 1442.040 1249.750 1442.180 ;
        RECT 1249.430 1441.980 1249.750 1442.040 ;
        RECT 1249.430 1429.260 1249.750 1429.320 ;
        RECT 1249.235 1429.120 1249.750 1429.260 ;
        RECT 1249.430 1429.060 1249.750 1429.120 ;
        RECT 1249.445 1393.900 1249.735 1393.945 ;
        RECT 1250.350 1393.900 1250.670 1393.960 ;
        RECT 1249.445 1393.760 1250.670 1393.900 ;
        RECT 1249.445 1393.715 1249.735 1393.760 ;
        RECT 1250.350 1393.700 1250.670 1393.760 ;
        RECT 1249.890 1303.940 1250.210 1304.200 ;
        RECT 1249.980 1303.800 1250.120 1303.940 ;
        RECT 1250.350 1303.800 1250.670 1303.860 ;
        RECT 1249.980 1303.660 1250.670 1303.800 ;
        RECT 1250.350 1303.600 1250.670 1303.660 ;
        RECT 1250.350 869.960 1250.670 870.020 ;
        RECT 1249.980 869.820 1250.670 869.960 ;
        RECT 1249.980 869.340 1250.120 869.820 ;
        RECT 1250.350 869.760 1250.670 869.820 ;
        RECT 1249.890 869.080 1250.210 869.340 ;
        RECT 1249.890 689.900 1250.210 690.160 ;
        RECT 1249.980 689.480 1250.120 689.900 ;
        RECT 1249.890 689.220 1250.210 689.480 ;
        RECT 1249.890 282.780 1250.210 282.840 ;
        RECT 1249.695 282.640 1250.210 282.780 ;
        RECT 1249.890 282.580 1250.210 282.640 ;
        RECT 1249.890 234.840 1250.210 234.900 ;
        RECT 1249.695 234.700 1250.210 234.840 ;
        RECT 1249.890 234.640 1250.210 234.700 ;
        RECT 1249.890 48.520 1250.210 48.580 ;
        RECT 1250.350 48.520 1250.670 48.580 ;
        RECT 1249.890 48.380 1250.670 48.520 ;
        RECT 1249.890 48.320 1250.210 48.380 ;
        RECT 1250.350 48.320 1250.670 48.380 ;
        RECT 204.770 40.020 205.090 40.080 ;
        RECT 1249.890 40.020 1250.210 40.080 ;
        RECT 204.770 39.880 1250.210 40.020 ;
        RECT 204.770 39.820 205.090 39.880 ;
        RECT 1249.890 39.820 1250.210 39.880 ;
      LAYER via ;
        RECT 1249.920 1688.480 1250.180 1688.740 ;
        RECT 1254.060 1688.480 1254.320 1688.740 ;
        RECT 1249.920 1608.240 1250.180 1608.500 ;
        RECT 1249.920 1587.160 1250.180 1587.420 ;
        RECT 1249.920 1559.280 1250.180 1559.540 ;
        RECT 1249.460 1558.940 1249.720 1559.200 ;
        RECT 1249.460 1490.260 1249.720 1490.520 ;
        RECT 1249.460 1441.980 1249.720 1442.240 ;
        RECT 1249.460 1429.060 1249.720 1429.320 ;
        RECT 1250.380 1393.700 1250.640 1393.960 ;
        RECT 1249.920 1303.940 1250.180 1304.200 ;
        RECT 1250.380 1303.600 1250.640 1303.860 ;
        RECT 1250.380 869.760 1250.640 870.020 ;
        RECT 1249.920 869.080 1250.180 869.340 ;
        RECT 1249.920 689.900 1250.180 690.160 ;
        RECT 1249.920 689.220 1250.180 689.480 ;
        RECT 1249.920 282.580 1250.180 282.840 ;
        RECT 1249.920 234.640 1250.180 234.900 ;
        RECT 1249.920 48.320 1250.180 48.580 ;
        RECT 1250.380 48.320 1250.640 48.580 ;
        RECT 204.800 39.820 205.060 40.080 ;
        RECT 1249.920 39.820 1250.180 40.080 ;
      LAYER met2 ;
        RECT 1253.980 1700.000 1254.260 1702.400 ;
        RECT 1254.120 1688.770 1254.260 1700.000 ;
        RECT 1249.920 1688.450 1250.180 1688.770 ;
        RECT 1254.060 1688.450 1254.320 1688.770 ;
        RECT 1249.980 1608.530 1250.120 1688.450 ;
        RECT 1249.920 1608.210 1250.180 1608.530 ;
        RECT 1249.920 1587.130 1250.180 1587.450 ;
        RECT 1249.980 1559.570 1250.120 1587.130 ;
        RECT 1249.920 1559.250 1250.180 1559.570 ;
        RECT 1249.460 1558.910 1249.720 1559.230 ;
        RECT 1249.520 1512.050 1249.660 1558.910 ;
        RECT 1249.520 1511.910 1250.580 1512.050 ;
        RECT 1250.440 1497.090 1250.580 1511.910 ;
        RECT 1249.520 1496.950 1250.580 1497.090 ;
        RECT 1249.520 1490.550 1249.660 1496.950 ;
        RECT 1249.460 1490.230 1249.720 1490.550 ;
        RECT 1249.460 1441.950 1249.720 1442.270 ;
        RECT 1249.520 1429.350 1249.660 1441.950 ;
        RECT 1249.460 1429.030 1249.720 1429.350 ;
        RECT 1250.380 1393.670 1250.640 1393.990 ;
        RECT 1250.440 1365.850 1250.580 1393.670 ;
        RECT 1249.980 1365.710 1250.580 1365.850 ;
        RECT 1249.980 1304.230 1250.120 1365.710 ;
        RECT 1249.920 1303.910 1250.180 1304.230 ;
        RECT 1250.380 1303.570 1250.640 1303.890 ;
        RECT 1250.440 1269.290 1250.580 1303.570 ;
        RECT 1249.980 1269.150 1250.580 1269.290 ;
        RECT 1249.980 980.290 1250.120 1269.150 ;
        RECT 1249.520 980.150 1250.120 980.290 ;
        RECT 1249.520 979.610 1249.660 980.150 ;
        RECT 1249.520 979.470 1250.120 979.610 ;
        RECT 1249.980 934.730 1250.120 979.470 ;
        RECT 1249.980 934.590 1250.580 934.730 ;
        RECT 1250.440 870.050 1250.580 934.590 ;
        RECT 1250.380 869.730 1250.640 870.050 ;
        RECT 1249.920 869.050 1250.180 869.370 ;
        RECT 1249.980 787.170 1250.120 869.050 ;
        RECT 1249.520 787.030 1250.120 787.170 ;
        RECT 1249.520 786.490 1249.660 787.030 ;
        RECT 1249.520 786.350 1250.120 786.490 ;
        RECT 1249.980 690.190 1250.120 786.350 ;
        RECT 1249.920 689.870 1250.180 690.190 ;
        RECT 1249.920 689.190 1250.180 689.510 ;
        RECT 1249.980 303.690 1250.120 689.190 ;
        RECT 1249.520 303.550 1250.120 303.690 ;
        RECT 1249.520 303.010 1249.660 303.550 ;
        RECT 1249.520 302.870 1250.120 303.010 ;
        RECT 1249.980 282.870 1250.120 302.870 ;
        RECT 1249.920 282.550 1250.180 282.870 ;
        RECT 1249.920 234.610 1250.180 234.930 ;
        RECT 1249.980 144.570 1250.120 234.610 ;
        RECT 1249.980 144.430 1250.580 144.570 ;
        RECT 1250.440 48.610 1250.580 144.430 ;
        RECT 1249.920 48.290 1250.180 48.610 ;
        RECT 1250.380 48.290 1250.640 48.610 ;
        RECT 1249.980 40.110 1250.120 48.290 ;
        RECT 204.800 39.790 205.060 40.110 ;
        RECT 1249.920 39.790 1250.180 40.110 ;
        RECT 204.860 2.400 205.000 39.790 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1263.305 1600.465 1263.475 1642.115 ;
      LAYER mcon ;
        RECT 1263.305 1641.945 1263.475 1642.115 ;
      LAYER met1 ;
        RECT 1263.230 1642.100 1263.550 1642.160 ;
        RECT 1263.035 1641.960 1263.550 1642.100 ;
        RECT 1263.230 1641.900 1263.550 1641.960 ;
        RECT 1263.230 1600.620 1263.550 1600.680 ;
        RECT 1263.035 1600.480 1263.550 1600.620 ;
        RECT 1263.230 1600.420 1263.550 1600.480 ;
        RECT 222.710 40.360 223.030 40.420 ;
        RECT 1263.230 40.360 1263.550 40.420 ;
        RECT 222.710 40.220 1263.550 40.360 ;
        RECT 222.710 40.160 223.030 40.220 ;
        RECT 1263.230 40.160 1263.550 40.220 ;
      LAYER via ;
        RECT 1263.260 1641.900 1263.520 1642.160 ;
        RECT 1263.260 1600.420 1263.520 1600.680 ;
        RECT 222.740 40.160 223.000 40.420 ;
        RECT 1263.260 40.160 1263.520 40.420 ;
      LAYER met2 ;
        RECT 1263.180 1700.000 1263.460 1702.400 ;
        RECT 1263.320 1642.190 1263.460 1700.000 ;
        RECT 1263.260 1641.870 1263.520 1642.190 ;
        RECT 1263.260 1600.390 1263.520 1600.710 ;
        RECT 1263.320 40.450 1263.460 1600.390 ;
        RECT 222.740 40.130 223.000 40.450 ;
        RECT 1263.260 40.130 1263.520 40.450 ;
        RECT 222.800 2.400 222.940 40.130 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1153.365 1594.005 1153.535 1627.835 ;
        RECT 1153.365 1497.445 1153.535 1521.415 ;
        RECT 1154.285 1366.205 1154.455 1400.715 ;
        RECT 1154.745 1220.685 1154.915 1272.195 ;
        RECT 1154.285 448.205 1154.455 483.055 ;
        RECT 1154.745 386.325 1154.915 400.775 ;
        RECT 1154.745 331.245 1154.915 379.355 ;
        RECT 1153.365 41.565 1153.535 131.155 ;
      LAYER mcon ;
        RECT 1153.365 1627.665 1153.535 1627.835 ;
        RECT 1153.365 1521.245 1153.535 1521.415 ;
        RECT 1154.285 1400.545 1154.455 1400.715 ;
        RECT 1154.745 1272.025 1154.915 1272.195 ;
        RECT 1154.285 482.885 1154.455 483.055 ;
        RECT 1154.745 400.605 1154.915 400.775 ;
        RECT 1154.745 379.185 1154.915 379.355 ;
        RECT 1153.365 130.985 1153.535 131.155 ;
      LAYER met1 ;
        RECT 1153.290 1627.820 1153.610 1627.880 ;
        RECT 1153.095 1627.680 1153.610 1627.820 ;
        RECT 1153.290 1627.620 1153.610 1627.680 ;
        RECT 1153.305 1594.160 1153.595 1594.205 ;
        RECT 1154.210 1594.160 1154.530 1594.220 ;
        RECT 1153.305 1594.020 1154.530 1594.160 ;
        RECT 1153.305 1593.975 1153.595 1594.020 ;
        RECT 1154.210 1593.960 1154.530 1594.020 ;
        RECT 1153.290 1559.480 1153.610 1559.540 ;
        RECT 1154.210 1559.480 1154.530 1559.540 ;
        RECT 1153.290 1559.340 1154.530 1559.480 ;
        RECT 1153.290 1559.280 1153.610 1559.340 ;
        RECT 1154.210 1559.280 1154.530 1559.340 ;
        RECT 1153.290 1521.400 1153.610 1521.460 ;
        RECT 1153.095 1521.260 1153.610 1521.400 ;
        RECT 1153.290 1521.200 1153.610 1521.260 ;
        RECT 1153.305 1497.600 1153.595 1497.645 ;
        RECT 1154.210 1497.600 1154.530 1497.660 ;
        RECT 1153.305 1497.460 1154.530 1497.600 ;
        RECT 1153.305 1497.415 1153.595 1497.460 ;
        RECT 1154.210 1497.400 1154.530 1497.460 ;
        RECT 1153.290 1462.920 1153.610 1462.980 ;
        RECT 1154.210 1462.920 1154.530 1462.980 ;
        RECT 1153.290 1462.780 1154.530 1462.920 ;
        RECT 1153.290 1462.720 1153.610 1462.780 ;
        RECT 1154.210 1462.720 1154.530 1462.780 ;
        RECT 1153.290 1414.780 1153.610 1415.040 ;
        RECT 1153.380 1414.360 1153.520 1414.780 ;
        RECT 1153.290 1414.100 1153.610 1414.360 ;
        RECT 1153.290 1400.700 1153.610 1400.760 ;
        RECT 1154.225 1400.700 1154.515 1400.745 ;
        RECT 1153.290 1400.560 1154.515 1400.700 ;
        RECT 1153.290 1400.500 1153.610 1400.560 ;
        RECT 1154.225 1400.515 1154.515 1400.560 ;
        RECT 1154.210 1366.360 1154.530 1366.420 ;
        RECT 1154.015 1366.220 1154.530 1366.360 ;
        RECT 1154.210 1366.160 1154.530 1366.220 ;
        RECT 1154.210 1317.880 1154.530 1318.140 ;
        RECT 1154.300 1317.400 1154.440 1317.880 ;
        RECT 1154.670 1317.400 1154.990 1317.460 ;
        RECT 1154.300 1317.260 1154.990 1317.400 ;
        RECT 1154.670 1317.200 1154.990 1317.260 ;
        RECT 1154.670 1272.180 1154.990 1272.240 ;
        RECT 1154.475 1272.040 1154.990 1272.180 ;
        RECT 1154.670 1271.980 1154.990 1272.040 ;
        RECT 1154.670 1220.840 1154.990 1220.900 ;
        RECT 1154.475 1220.700 1154.990 1220.840 ;
        RECT 1154.670 1220.640 1154.990 1220.700 ;
        RECT 1154.670 1173.580 1154.990 1173.640 ;
        RECT 1154.300 1173.440 1154.990 1173.580 ;
        RECT 1154.300 1172.960 1154.440 1173.440 ;
        RECT 1154.670 1173.380 1154.990 1173.440 ;
        RECT 1154.210 1172.700 1154.530 1172.960 ;
        RECT 1153.290 1111.020 1153.610 1111.080 ;
        RECT 1154.670 1111.020 1154.990 1111.080 ;
        RECT 1153.290 1110.880 1154.990 1111.020 ;
        RECT 1153.290 1110.820 1153.610 1110.880 ;
        RECT 1154.670 1110.820 1154.990 1110.880 ;
        RECT 1154.670 1077.020 1154.990 1077.080 ;
        RECT 1154.300 1076.880 1154.990 1077.020 ;
        RECT 1154.300 1076.400 1154.440 1076.880 ;
        RECT 1154.670 1076.820 1154.990 1076.880 ;
        RECT 1154.210 1076.140 1154.530 1076.400 ;
        RECT 1153.290 1014.460 1153.610 1014.520 ;
        RECT 1154.670 1014.460 1154.990 1014.520 ;
        RECT 1153.290 1014.320 1154.990 1014.460 ;
        RECT 1153.290 1014.260 1153.610 1014.320 ;
        RECT 1154.670 1014.260 1154.990 1014.320 ;
        RECT 1154.670 980.460 1154.990 980.520 ;
        RECT 1154.300 980.320 1154.990 980.460 ;
        RECT 1154.300 979.840 1154.440 980.320 ;
        RECT 1154.670 980.260 1154.990 980.320 ;
        RECT 1154.210 979.580 1154.530 979.840 ;
        RECT 1153.290 917.900 1153.610 917.960 ;
        RECT 1154.670 917.900 1154.990 917.960 ;
        RECT 1153.290 917.760 1154.990 917.900 ;
        RECT 1153.290 917.700 1153.610 917.760 ;
        RECT 1154.670 917.700 1154.990 917.760 ;
        RECT 1153.750 872.000 1154.070 872.060 ;
        RECT 1154.670 872.000 1154.990 872.060 ;
        RECT 1153.750 871.860 1154.990 872.000 ;
        RECT 1153.750 871.800 1154.070 871.860 ;
        RECT 1154.670 871.800 1154.990 871.860 ;
        RECT 1153.750 834.940 1154.070 835.000 ;
        RECT 1154.670 834.940 1154.990 835.000 ;
        RECT 1153.750 834.800 1154.990 834.940 ;
        RECT 1153.750 834.740 1154.070 834.800 ;
        RECT 1154.670 834.740 1154.990 834.800 ;
        RECT 1153.290 821.000 1153.610 821.060 ;
        RECT 1154.670 821.000 1154.990 821.060 ;
        RECT 1153.290 820.860 1154.990 821.000 ;
        RECT 1153.290 820.800 1153.610 820.860 ;
        RECT 1154.670 820.800 1154.990 820.860 ;
        RECT 1154.210 772.720 1154.530 772.780 ;
        RECT 1155.130 772.720 1155.450 772.780 ;
        RECT 1154.210 772.580 1155.450 772.720 ;
        RECT 1154.210 772.520 1154.530 772.580 ;
        RECT 1155.130 772.520 1155.450 772.580 ;
        RECT 1153.750 689.900 1154.070 690.160 ;
        RECT 1153.840 689.760 1153.980 689.900 ;
        RECT 1154.210 689.760 1154.530 689.820 ;
        RECT 1153.840 689.620 1154.530 689.760 ;
        RECT 1154.210 689.560 1154.530 689.620 ;
        RECT 1154.210 676.160 1154.530 676.220 ;
        RECT 1155.130 676.160 1155.450 676.220 ;
        RECT 1154.210 676.020 1155.450 676.160 ;
        RECT 1154.210 675.960 1154.530 676.020 ;
        RECT 1155.130 675.960 1155.450 676.020 ;
        RECT 1153.750 593.340 1154.070 593.600 ;
        RECT 1153.840 593.200 1153.980 593.340 ;
        RECT 1154.210 593.200 1154.530 593.260 ;
        RECT 1153.840 593.060 1154.530 593.200 ;
        RECT 1154.210 593.000 1154.530 593.060 ;
        RECT 1154.210 579.600 1154.530 579.660 ;
        RECT 1155.130 579.600 1155.450 579.660 ;
        RECT 1154.210 579.460 1155.450 579.600 ;
        RECT 1154.210 579.400 1154.530 579.460 ;
        RECT 1155.130 579.400 1155.450 579.460 ;
        RECT 1153.750 496.780 1154.070 497.040 ;
        RECT 1153.840 496.640 1153.980 496.780 ;
        RECT 1154.210 496.640 1154.530 496.700 ;
        RECT 1153.840 496.500 1154.530 496.640 ;
        RECT 1154.210 496.440 1154.530 496.500 ;
        RECT 1154.210 483.040 1154.530 483.100 ;
        RECT 1154.015 482.900 1154.530 483.040 ;
        RECT 1154.210 482.840 1154.530 482.900 ;
        RECT 1154.210 448.360 1154.530 448.420 ;
        RECT 1154.015 448.220 1154.530 448.360 ;
        RECT 1154.210 448.160 1154.530 448.220 ;
        RECT 1154.670 400.760 1154.990 400.820 ;
        RECT 1154.475 400.620 1154.990 400.760 ;
        RECT 1154.670 400.560 1154.990 400.620 ;
        RECT 1154.670 386.480 1154.990 386.540 ;
        RECT 1154.475 386.340 1154.990 386.480 ;
        RECT 1154.670 386.280 1154.990 386.340 ;
        RECT 1154.670 379.340 1154.990 379.400 ;
        RECT 1154.475 379.200 1154.990 379.340 ;
        RECT 1154.670 379.140 1154.990 379.200 ;
        RECT 1154.685 331.400 1154.975 331.445 ;
        RECT 1155.130 331.400 1155.450 331.460 ;
        RECT 1154.685 331.260 1155.450 331.400 ;
        RECT 1154.685 331.215 1154.975 331.260 ;
        RECT 1155.130 331.200 1155.450 331.260 ;
        RECT 1153.290 217.500 1153.610 217.560 ;
        RECT 1154.210 217.500 1154.530 217.560 ;
        RECT 1153.290 217.360 1154.530 217.500 ;
        RECT 1153.290 217.300 1153.610 217.360 ;
        RECT 1154.210 217.300 1154.530 217.360 ;
        RECT 1153.290 186.220 1153.610 186.280 ;
        RECT 1153.750 186.220 1154.070 186.280 ;
        RECT 1153.290 186.080 1154.070 186.220 ;
        RECT 1153.290 186.020 1153.610 186.080 ;
        RECT 1153.750 186.020 1154.070 186.080 ;
        RECT 1153.750 137.940 1154.070 138.000 ;
        RECT 1154.210 137.940 1154.530 138.000 ;
        RECT 1153.750 137.800 1154.530 137.940 ;
        RECT 1153.750 137.740 1154.070 137.800 ;
        RECT 1154.210 137.740 1154.530 137.800 ;
        RECT 1153.305 131.140 1153.595 131.185 ;
        RECT 1153.750 131.140 1154.070 131.200 ;
        RECT 1153.305 131.000 1154.070 131.140 ;
        RECT 1153.305 130.955 1153.595 131.000 ;
        RECT 1153.750 130.940 1154.070 131.000 ;
        RECT 1153.290 41.720 1153.610 41.780 ;
        RECT 1153.095 41.580 1153.610 41.720 ;
        RECT 1153.290 41.520 1153.610 41.580 ;
        RECT 19.850 37.980 20.170 38.040 ;
        RECT 1153.290 37.980 1153.610 38.040 ;
        RECT 19.850 37.840 1153.610 37.980 ;
        RECT 19.850 37.780 20.170 37.840 ;
        RECT 1153.290 37.780 1153.610 37.840 ;
      LAYER via ;
        RECT 1153.320 1627.620 1153.580 1627.880 ;
        RECT 1154.240 1593.960 1154.500 1594.220 ;
        RECT 1153.320 1559.280 1153.580 1559.540 ;
        RECT 1154.240 1559.280 1154.500 1559.540 ;
        RECT 1153.320 1521.200 1153.580 1521.460 ;
        RECT 1154.240 1497.400 1154.500 1497.660 ;
        RECT 1153.320 1462.720 1153.580 1462.980 ;
        RECT 1154.240 1462.720 1154.500 1462.980 ;
        RECT 1153.320 1414.780 1153.580 1415.040 ;
        RECT 1153.320 1414.100 1153.580 1414.360 ;
        RECT 1153.320 1400.500 1153.580 1400.760 ;
        RECT 1154.240 1366.160 1154.500 1366.420 ;
        RECT 1154.240 1317.880 1154.500 1318.140 ;
        RECT 1154.700 1317.200 1154.960 1317.460 ;
        RECT 1154.700 1271.980 1154.960 1272.240 ;
        RECT 1154.700 1220.640 1154.960 1220.900 ;
        RECT 1154.700 1173.380 1154.960 1173.640 ;
        RECT 1154.240 1172.700 1154.500 1172.960 ;
        RECT 1153.320 1110.820 1153.580 1111.080 ;
        RECT 1154.700 1110.820 1154.960 1111.080 ;
        RECT 1154.700 1076.820 1154.960 1077.080 ;
        RECT 1154.240 1076.140 1154.500 1076.400 ;
        RECT 1153.320 1014.260 1153.580 1014.520 ;
        RECT 1154.700 1014.260 1154.960 1014.520 ;
        RECT 1154.700 980.260 1154.960 980.520 ;
        RECT 1154.240 979.580 1154.500 979.840 ;
        RECT 1153.320 917.700 1153.580 917.960 ;
        RECT 1154.700 917.700 1154.960 917.960 ;
        RECT 1153.780 871.800 1154.040 872.060 ;
        RECT 1154.700 871.800 1154.960 872.060 ;
        RECT 1153.780 834.740 1154.040 835.000 ;
        RECT 1154.700 834.740 1154.960 835.000 ;
        RECT 1153.320 820.800 1153.580 821.060 ;
        RECT 1154.700 820.800 1154.960 821.060 ;
        RECT 1154.240 772.520 1154.500 772.780 ;
        RECT 1155.160 772.520 1155.420 772.780 ;
        RECT 1153.780 689.900 1154.040 690.160 ;
        RECT 1154.240 689.560 1154.500 689.820 ;
        RECT 1154.240 675.960 1154.500 676.220 ;
        RECT 1155.160 675.960 1155.420 676.220 ;
        RECT 1153.780 593.340 1154.040 593.600 ;
        RECT 1154.240 593.000 1154.500 593.260 ;
        RECT 1154.240 579.400 1154.500 579.660 ;
        RECT 1155.160 579.400 1155.420 579.660 ;
        RECT 1153.780 496.780 1154.040 497.040 ;
        RECT 1154.240 496.440 1154.500 496.700 ;
        RECT 1154.240 482.840 1154.500 483.100 ;
        RECT 1154.240 448.160 1154.500 448.420 ;
        RECT 1154.700 400.560 1154.960 400.820 ;
        RECT 1154.700 386.280 1154.960 386.540 ;
        RECT 1154.700 379.140 1154.960 379.400 ;
        RECT 1155.160 331.200 1155.420 331.460 ;
        RECT 1153.320 217.300 1153.580 217.560 ;
        RECT 1154.240 217.300 1154.500 217.560 ;
        RECT 1153.320 186.020 1153.580 186.280 ;
        RECT 1153.780 186.020 1154.040 186.280 ;
        RECT 1153.780 137.740 1154.040 138.000 ;
        RECT 1154.240 137.740 1154.500 138.000 ;
        RECT 1153.780 130.940 1154.040 131.200 ;
        RECT 1153.320 41.520 1153.580 41.780 ;
        RECT 19.880 37.780 20.140 38.040 ;
        RECT 1153.320 37.780 1153.580 38.040 ;
      LAYER met2 ;
        RECT 1158.760 1701.090 1159.040 1702.400 ;
        RECT 1156.600 1700.950 1159.040 1701.090 ;
        RECT 1156.600 1677.290 1156.740 1700.950 ;
        RECT 1158.760 1700.000 1159.040 1700.950 ;
        RECT 1153.380 1677.150 1156.740 1677.290 ;
        RECT 1153.380 1627.910 1153.520 1677.150 ;
        RECT 1153.320 1627.590 1153.580 1627.910 ;
        RECT 1154.240 1593.930 1154.500 1594.250 ;
        RECT 1154.300 1559.570 1154.440 1593.930 ;
        RECT 1153.320 1559.250 1153.580 1559.570 ;
        RECT 1154.240 1559.250 1154.500 1559.570 ;
        RECT 1153.380 1521.490 1153.520 1559.250 ;
        RECT 1153.320 1521.170 1153.580 1521.490 ;
        RECT 1154.240 1497.370 1154.500 1497.690 ;
        RECT 1154.300 1463.010 1154.440 1497.370 ;
        RECT 1153.320 1462.690 1153.580 1463.010 ;
        RECT 1154.240 1462.690 1154.500 1463.010 ;
        RECT 1153.380 1415.070 1153.520 1462.690 ;
        RECT 1153.320 1414.750 1153.580 1415.070 ;
        RECT 1153.320 1414.070 1153.580 1414.390 ;
        RECT 1153.380 1400.790 1153.520 1414.070 ;
        RECT 1153.320 1400.470 1153.580 1400.790 ;
        RECT 1154.240 1366.130 1154.500 1366.450 ;
        RECT 1154.300 1318.170 1154.440 1366.130 ;
        RECT 1154.240 1317.850 1154.500 1318.170 ;
        RECT 1154.700 1317.170 1154.960 1317.490 ;
        RECT 1154.760 1272.270 1154.900 1317.170 ;
        RECT 1154.700 1271.950 1154.960 1272.270 ;
        RECT 1154.700 1220.610 1154.960 1220.930 ;
        RECT 1154.760 1173.670 1154.900 1220.610 ;
        RECT 1154.700 1173.350 1154.960 1173.670 ;
        RECT 1154.240 1172.670 1154.500 1172.990 ;
        RECT 1154.300 1159.245 1154.440 1172.670 ;
        RECT 1153.310 1158.875 1153.590 1159.245 ;
        RECT 1154.230 1158.875 1154.510 1159.245 ;
        RECT 1153.380 1111.110 1153.520 1158.875 ;
        RECT 1153.320 1110.790 1153.580 1111.110 ;
        RECT 1154.700 1110.790 1154.960 1111.110 ;
        RECT 1154.760 1077.110 1154.900 1110.790 ;
        RECT 1154.700 1076.790 1154.960 1077.110 ;
        RECT 1154.240 1076.110 1154.500 1076.430 ;
        RECT 1154.300 1062.685 1154.440 1076.110 ;
        RECT 1153.310 1062.315 1153.590 1062.685 ;
        RECT 1154.230 1062.315 1154.510 1062.685 ;
        RECT 1153.380 1014.550 1153.520 1062.315 ;
        RECT 1153.320 1014.230 1153.580 1014.550 ;
        RECT 1154.700 1014.230 1154.960 1014.550 ;
        RECT 1154.760 980.550 1154.900 1014.230 ;
        RECT 1154.700 980.230 1154.960 980.550 ;
        RECT 1154.240 979.550 1154.500 979.870 ;
        RECT 1154.300 966.125 1154.440 979.550 ;
        RECT 1153.310 965.755 1153.590 966.125 ;
        RECT 1154.230 965.755 1154.510 966.125 ;
        RECT 1153.380 917.990 1153.520 965.755 ;
        RECT 1153.320 917.670 1153.580 917.990 ;
        RECT 1154.700 917.670 1154.960 917.990 ;
        RECT 1154.760 872.090 1154.900 917.670 ;
        RECT 1153.780 871.770 1154.040 872.090 ;
        RECT 1154.700 871.770 1154.960 872.090 ;
        RECT 1153.840 835.030 1153.980 871.770 ;
        RECT 1153.780 834.710 1154.040 835.030 ;
        RECT 1154.700 834.710 1154.960 835.030 ;
        RECT 1154.760 821.090 1154.900 834.710 ;
        RECT 1153.320 820.770 1153.580 821.090 ;
        RECT 1154.700 820.770 1154.960 821.090 ;
        RECT 1153.380 773.005 1153.520 820.770 ;
        RECT 1153.310 772.635 1153.590 773.005 ;
        RECT 1154.230 772.635 1154.510 773.005 ;
        RECT 1154.240 772.490 1154.500 772.635 ;
        RECT 1155.160 772.490 1155.420 772.810 ;
        RECT 1155.220 724.725 1155.360 772.490 ;
        RECT 1153.770 724.355 1154.050 724.725 ;
        RECT 1155.150 724.355 1155.430 724.725 ;
        RECT 1153.840 690.190 1153.980 724.355 ;
        RECT 1153.780 689.870 1154.040 690.190 ;
        RECT 1154.240 689.530 1154.500 689.850 ;
        RECT 1154.300 676.250 1154.440 689.530 ;
        RECT 1154.240 675.930 1154.500 676.250 ;
        RECT 1155.160 675.930 1155.420 676.250 ;
        RECT 1155.220 628.165 1155.360 675.930 ;
        RECT 1153.770 627.795 1154.050 628.165 ;
        RECT 1155.150 627.795 1155.430 628.165 ;
        RECT 1153.840 593.630 1153.980 627.795 ;
        RECT 1153.780 593.310 1154.040 593.630 ;
        RECT 1154.240 592.970 1154.500 593.290 ;
        RECT 1154.300 579.690 1154.440 592.970 ;
        RECT 1154.240 579.370 1154.500 579.690 ;
        RECT 1155.160 579.370 1155.420 579.690 ;
        RECT 1155.220 531.605 1155.360 579.370 ;
        RECT 1153.770 531.235 1154.050 531.605 ;
        RECT 1155.150 531.235 1155.430 531.605 ;
        RECT 1153.840 497.070 1153.980 531.235 ;
        RECT 1153.780 496.750 1154.040 497.070 ;
        RECT 1154.240 496.410 1154.500 496.730 ;
        RECT 1154.300 483.130 1154.440 496.410 ;
        RECT 1154.240 482.810 1154.500 483.130 ;
        RECT 1154.240 448.130 1154.500 448.450 ;
        RECT 1154.300 434.930 1154.440 448.130 ;
        RECT 1154.300 434.790 1154.900 434.930 ;
        RECT 1154.760 400.850 1154.900 434.790 ;
        RECT 1154.700 400.530 1154.960 400.850 ;
        RECT 1154.700 386.250 1154.960 386.570 ;
        RECT 1154.760 379.430 1154.900 386.250 ;
        RECT 1154.700 379.110 1154.960 379.430 ;
        RECT 1155.160 331.170 1155.420 331.490 ;
        RECT 1155.220 307.090 1155.360 331.170 ;
        RECT 1153.840 306.950 1155.360 307.090 ;
        RECT 1153.840 255.410 1153.980 306.950 ;
        RECT 1153.840 255.270 1154.440 255.410 ;
        RECT 1154.300 217.590 1154.440 255.270 ;
        RECT 1153.320 217.270 1153.580 217.590 ;
        RECT 1154.240 217.270 1154.500 217.590 ;
        RECT 1153.380 186.310 1153.520 217.270 ;
        RECT 1153.320 185.990 1153.580 186.310 ;
        RECT 1153.780 185.990 1154.040 186.310 ;
        RECT 1153.840 138.450 1153.980 185.990 ;
        RECT 1153.840 138.310 1154.440 138.450 ;
        RECT 1154.300 138.030 1154.440 138.310 ;
        RECT 1153.780 137.710 1154.040 138.030 ;
        RECT 1154.240 137.710 1154.500 138.030 ;
        RECT 1153.840 131.230 1153.980 137.710 ;
        RECT 1153.780 130.910 1154.040 131.230 ;
        RECT 1153.320 41.490 1153.580 41.810 ;
        RECT 1153.380 38.070 1153.520 41.490 ;
        RECT 19.880 37.750 20.140 38.070 ;
        RECT 1153.320 37.750 1153.580 38.070 ;
        RECT 19.940 3.130 20.080 37.750 ;
        RECT 19.940 2.990 20.540 3.130 ;
        RECT 20.400 2.400 20.540 2.990 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 1153.310 1158.920 1153.590 1159.200 ;
        RECT 1154.230 1158.920 1154.510 1159.200 ;
        RECT 1153.310 1062.360 1153.590 1062.640 ;
        RECT 1154.230 1062.360 1154.510 1062.640 ;
        RECT 1153.310 965.800 1153.590 966.080 ;
        RECT 1154.230 965.800 1154.510 966.080 ;
        RECT 1153.310 772.680 1153.590 772.960 ;
        RECT 1154.230 772.680 1154.510 772.960 ;
        RECT 1153.770 724.400 1154.050 724.680 ;
        RECT 1155.150 724.400 1155.430 724.680 ;
        RECT 1153.770 627.840 1154.050 628.120 ;
        RECT 1155.150 627.840 1155.430 628.120 ;
        RECT 1153.770 531.280 1154.050 531.560 ;
        RECT 1155.150 531.280 1155.430 531.560 ;
      LAYER met3 ;
        RECT 1153.285 1159.210 1153.615 1159.225 ;
        RECT 1154.205 1159.210 1154.535 1159.225 ;
        RECT 1153.285 1158.910 1154.535 1159.210 ;
        RECT 1153.285 1158.895 1153.615 1158.910 ;
        RECT 1154.205 1158.895 1154.535 1158.910 ;
        RECT 1153.285 1062.650 1153.615 1062.665 ;
        RECT 1154.205 1062.650 1154.535 1062.665 ;
        RECT 1153.285 1062.350 1154.535 1062.650 ;
        RECT 1153.285 1062.335 1153.615 1062.350 ;
        RECT 1154.205 1062.335 1154.535 1062.350 ;
        RECT 1153.285 966.090 1153.615 966.105 ;
        RECT 1154.205 966.090 1154.535 966.105 ;
        RECT 1153.285 965.790 1154.535 966.090 ;
        RECT 1153.285 965.775 1153.615 965.790 ;
        RECT 1154.205 965.775 1154.535 965.790 ;
        RECT 1153.285 772.970 1153.615 772.985 ;
        RECT 1154.205 772.970 1154.535 772.985 ;
        RECT 1153.285 772.670 1154.535 772.970 ;
        RECT 1153.285 772.655 1153.615 772.670 ;
        RECT 1154.205 772.655 1154.535 772.670 ;
        RECT 1153.745 724.690 1154.075 724.705 ;
        RECT 1155.125 724.690 1155.455 724.705 ;
        RECT 1153.745 724.390 1155.455 724.690 ;
        RECT 1153.745 724.375 1154.075 724.390 ;
        RECT 1155.125 724.375 1155.455 724.390 ;
        RECT 1153.745 628.130 1154.075 628.145 ;
        RECT 1155.125 628.130 1155.455 628.145 ;
        RECT 1153.745 627.830 1155.455 628.130 ;
        RECT 1153.745 627.815 1154.075 627.830 ;
        RECT 1155.125 627.815 1155.455 627.830 ;
        RECT 1153.745 531.570 1154.075 531.585 ;
        RECT 1155.125 531.570 1155.455 531.585 ;
        RECT 1153.745 531.270 1155.455 531.570 ;
        RECT 1153.745 531.255 1154.075 531.270 ;
        RECT 1155.125 531.255 1155.455 531.270 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1166.630 1400.700 1166.950 1400.760 ;
        RECT 1167.550 1400.700 1167.870 1400.760 ;
        RECT 1166.630 1400.560 1167.870 1400.700 ;
        RECT 1166.630 1400.500 1166.950 1400.560 ;
        RECT 1167.550 1400.500 1167.870 1400.560 ;
        RECT 1166.630 1221.520 1166.950 1221.580 ;
        RECT 1167.550 1221.520 1167.870 1221.580 ;
        RECT 1166.630 1221.380 1167.870 1221.520 ;
        RECT 1166.630 1221.320 1166.950 1221.380 ;
        RECT 1167.550 1221.320 1167.870 1221.380 ;
        RECT 1166.630 1124.960 1166.950 1125.020 ;
        RECT 1167.550 1124.960 1167.870 1125.020 ;
        RECT 1166.630 1124.820 1167.870 1124.960 ;
        RECT 1166.630 1124.760 1166.950 1124.820 ;
        RECT 1167.550 1124.760 1167.870 1124.820 ;
        RECT 1166.630 1076.340 1166.950 1076.400 ;
        RECT 1167.550 1076.340 1167.870 1076.400 ;
        RECT 1166.630 1076.200 1167.870 1076.340 ;
        RECT 1166.630 1076.140 1166.950 1076.200 ;
        RECT 1167.550 1076.140 1167.870 1076.200 ;
        RECT 1167.550 1025.820 1167.870 1026.080 ;
        RECT 1167.640 1025.400 1167.780 1025.820 ;
        RECT 1167.550 1025.140 1167.870 1025.400 ;
        RECT 1166.630 931.840 1166.950 931.900 ;
        RECT 1167.550 931.840 1167.870 931.900 ;
        RECT 1166.630 931.700 1167.870 931.840 ;
        RECT 1166.630 931.640 1166.950 931.700 ;
        RECT 1167.550 931.640 1167.870 931.700 ;
        RECT 1166.630 641.820 1166.950 641.880 ;
        RECT 1167.550 641.820 1167.870 641.880 ;
        RECT 1166.630 641.680 1167.870 641.820 ;
        RECT 1166.630 641.620 1166.950 641.680 ;
        RECT 1167.550 641.620 1167.870 641.680 ;
        RECT 1166.630 545.260 1166.950 545.320 ;
        RECT 1167.550 545.260 1167.870 545.320 ;
        RECT 1166.630 545.120 1167.870 545.260 ;
        RECT 1166.630 545.060 1166.950 545.120 ;
        RECT 1167.550 545.060 1167.870 545.120 ;
        RECT 1166.630 448.700 1166.950 448.760 ;
        RECT 1167.550 448.700 1167.870 448.760 ;
        RECT 1166.630 448.560 1167.870 448.700 ;
        RECT 1166.630 448.500 1166.950 448.560 ;
        RECT 1167.550 448.500 1167.870 448.560 ;
        RECT 1166.630 158.680 1166.950 158.740 ;
        RECT 1167.550 158.680 1167.870 158.740 ;
        RECT 1166.630 158.540 1167.870 158.680 ;
        RECT 1166.630 158.480 1166.950 158.540 ;
        RECT 1167.550 158.480 1167.870 158.540 ;
        RECT 1166.630 96.460 1166.950 96.520 ;
        RECT 1167.090 96.460 1167.410 96.520 ;
        RECT 1166.630 96.320 1167.410 96.460 ;
        RECT 1166.630 96.260 1166.950 96.320 ;
        RECT 1167.090 96.260 1167.410 96.320 ;
        RECT 44.230 38.320 44.550 38.380 ;
        RECT 1166.630 38.320 1166.950 38.380 ;
        RECT 44.230 38.180 1166.950 38.320 ;
        RECT 44.230 38.120 44.550 38.180 ;
        RECT 1166.630 38.120 1166.950 38.180 ;
      LAYER via ;
        RECT 1166.660 1400.500 1166.920 1400.760 ;
        RECT 1167.580 1400.500 1167.840 1400.760 ;
        RECT 1166.660 1221.320 1166.920 1221.580 ;
        RECT 1167.580 1221.320 1167.840 1221.580 ;
        RECT 1166.660 1124.760 1166.920 1125.020 ;
        RECT 1167.580 1124.760 1167.840 1125.020 ;
        RECT 1166.660 1076.140 1166.920 1076.400 ;
        RECT 1167.580 1076.140 1167.840 1076.400 ;
        RECT 1167.580 1025.820 1167.840 1026.080 ;
        RECT 1167.580 1025.140 1167.840 1025.400 ;
        RECT 1166.660 931.640 1166.920 931.900 ;
        RECT 1167.580 931.640 1167.840 931.900 ;
        RECT 1166.660 641.620 1166.920 641.880 ;
        RECT 1167.580 641.620 1167.840 641.880 ;
        RECT 1166.660 545.060 1166.920 545.320 ;
        RECT 1167.580 545.060 1167.840 545.320 ;
        RECT 1166.660 448.500 1166.920 448.760 ;
        RECT 1167.580 448.500 1167.840 448.760 ;
        RECT 1166.660 158.480 1166.920 158.740 ;
        RECT 1167.580 158.480 1167.840 158.740 ;
        RECT 1166.660 96.260 1166.920 96.520 ;
        RECT 1167.120 96.260 1167.380 96.520 ;
        RECT 44.260 38.120 44.520 38.380 ;
        RECT 1166.660 38.120 1166.920 38.380 ;
      LAYER met2 ;
        RECT 1171.180 1700.410 1171.460 1702.400 ;
        RECT 1169.020 1700.270 1171.460 1700.410 ;
        RECT 1169.020 1656.210 1169.160 1700.270 ;
        RECT 1171.180 1700.000 1171.460 1700.270 ;
        RECT 1166.720 1656.070 1169.160 1656.210 ;
        RECT 1166.720 1400.790 1166.860 1656.070 ;
        RECT 1166.660 1400.470 1166.920 1400.790 ;
        RECT 1167.580 1400.470 1167.840 1400.790 ;
        RECT 1167.640 1221.610 1167.780 1400.470 ;
        RECT 1166.660 1221.290 1166.920 1221.610 ;
        RECT 1167.580 1221.290 1167.840 1221.610 ;
        RECT 1166.720 1221.010 1166.860 1221.290 ;
        RECT 1166.720 1220.870 1167.320 1221.010 ;
        RECT 1167.180 1173.410 1167.320 1220.870 ;
        RECT 1167.180 1173.270 1167.780 1173.410 ;
        RECT 1167.640 1125.050 1167.780 1173.270 ;
        RECT 1166.660 1124.730 1166.920 1125.050 ;
        RECT 1167.580 1124.730 1167.840 1125.050 ;
        RECT 1166.720 1076.430 1166.860 1124.730 ;
        RECT 1166.660 1076.110 1166.920 1076.430 ;
        RECT 1167.580 1076.110 1167.840 1076.430 ;
        RECT 1167.640 1026.110 1167.780 1076.110 ;
        RECT 1167.580 1025.790 1167.840 1026.110 ;
        RECT 1167.580 1025.110 1167.840 1025.430 ;
        RECT 1167.640 931.930 1167.780 1025.110 ;
        RECT 1166.660 931.610 1166.920 931.930 ;
        RECT 1167.580 931.610 1167.840 931.930 ;
        RECT 1166.720 883.050 1166.860 931.610 ;
        RECT 1166.720 882.910 1167.320 883.050 ;
        RECT 1167.180 869.450 1167.320 882.910 ;
        RECT 1167.180 869.310 1167.780 869.450 ;
        RECT 1167.640 772.210 1167.780 869.310 ;
        RECT 1167.180 772.070 1167.780 772.210 ;
        RECT 1167.180 748.410 1167.320 772.070 ;
        RECT 1166.720 748.270 1167.320 748.410 ;
        RECT 1166.720 689.930 1166.860 748.270 ;
        RECT 1166.720 689.790 1167.780 689.930 ;
        RECT 1167.640 641.910 1167.780 689.790 ;
        RECT 1166.660 641.590 1166.920 641.910 ;
        RECT 1167.580 641.590 1167.840 641.910 ;
        RECT 1166.720 593.370 1166.860 641.590 ;
        RECT 1166.720 593.230 1167.780 593.370 ;
        RECT 1167.640 545.350 1167.780 593.230 ;
        RECT 1166.660 545.030 1166.920 545.350 ;
        RECT 1167.580 545.030 1167.840 545.350 ;
        RECT 1166.720 496.810 1166.860 545.030 ;
        RECT 1166.720 496.670 1167.780 496.810 ;
        RECT 1167.640 448.790 1167.780 496.670 ;
        RECT 1166.660 448.470 1166.920 448.790 ;
        RECT 1167.580 448.470 1167.840 448.790 ;
        RECT 1166.720 400.250 1166.860 448.470 ;
        RECT 1166.720 400.110 1167.780 400.250 ;
        RECT 1167.640 255.410 1167.780 400.110 ;
        RECT 1167.640 255.270 1168.240 255.410 ;
        RECT 1168.100 254.050 1168.240 255.270 ;
        RECT 1167.640 253.910 1168.240 254.050 ;
        RECT 1167.640 207.130 1167.780 253.910 ;
        RECT 1166.720 206.990 1167.780 207.130 ;
        RECT 1166.720 158.770 1166.860 206.990 ;
        RECT 1166.660 158.450 1166.920 158.770 ;
        RECT 1167.580 158.450 1167.840 158.770 ;
        RECT 1167.640 96.970 1167.780 158.450 ;
        RECT 1167.180 96.830 1167.780 96.970 ;
        RECT 1167.180 96.550 1167.320 96.830 ;
        RECT 1166.660 96.230 1166.920 96.550 ;
        RECT 1167.120 96.230 1167.380 96.550 ;
        RECT 1166.720 38.410 1166.860 96.230 ;
        RECT 44.260 38.090 44.520 38.410 ;
        RECT 1166.660 38.090 1166.920 38.410 ;
        RECT 44.320 2.400 44.460 38.090 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1270.665 862.665 1270.835 886.635 ;
        RECT 1270.665 544.765 1270.835 579.615 ;
        RECT 1270.665 386.325 1270.835 434.435 ;
      LAYER mcon ;
        RECT 1270.665 886.465 1270.835 886.635 ;
        RECT 1270.665 579.445 1270.835 579.615 ;
        RECT 1270.665 434.265 1270.835 434.435 ;
      LAYER met1 ;
        RECT 1270.590 1675.760 1270.910 1675.820 ;
        RECT 1275.190 1675.760 1275.510 1675.820 ;
        RECT 1270.590 1675.620 1275.510 1675.760 ;
        RECT 1270.590 1675.560 1270.910 1675.620 ;
        RECT 1275.190 1675.560 1275.510 1675.620 ;
        RECT 1271.050 1490.460 1271.370 1490.520 ;
        RECT 1272.430 1490.460 1272.750 1490.520 ;
        RECT 1271.050 1490.320 1272.750 1490.460 ;
        RECT 1271.050 1490.260 1271.370 1490.320 ;
        RECT 1272.430 1490.260 1272.750 1490.320 ;
        RECT 1271.050 1393.900 1271.370 1393.960 ;
        RECT 1272.430 1393.900 1272.750 1393.960 ;
        RECT 1271.050 1393.760 1272.750 1393.900 ;
        RECT 1271.050 1393.700 1271.370 1393.760 ;
        RECT 1272.430 1393.700 1272.750 1393.760 ;
        RECT 1271.050 1366.700 1271.370 1366.760 ;
        RECT 1270.680 1366.560 1271.370 1366.700 ;
        RECT 1270.680 1366.080 1270.820 1366.560 ;
        RECT 1271.050 1366.500 1271.370 1366.560 ;
        RECT 1270.590 1365.820 1270.910 1366.080 ;
        RECT 1270.130 1304.140 1270.450 1304.200 ;
        RECT 1271.050 1304.140 1271.370 1304.200 ;
        RECT 1270.130 1304.000 1271.370 1304.140 ;
        RECT 1270.130 1303.940 1270.450 1304.000 ;
        RECT 1271.050 1303.940 1271.370 1304.000 ;
        RECT 1270.130 1255.520 1270.450 1255.580 ;
        RECT 1271.050 1255.520 1271.370 1255.580 ;
        RECT 1270.130 1255.380 1271.370 1255.520 ;
        RECT 1270.130 1255.320 1270.450 1255.380 ;
        RECT 1271.050 1255.320 1271.370 1255.380 ;
        RECT 1270.130 1207.580 1270.450 1207.640 ;
        RECT 1271.050 1207.580 1271.370 1207.640 ;
        RECT 1270.130 1207.440 1271.370 1207.580 ;
        RECT 1270.130 1207.380 1270.450 1207.440 ;
        RECT 1271.050 1207.380 1271.370 1207.440 ;
        RECT 1270.590 1124.760 1270.910 1125.020 ;
        RECT 1270.680 1124.280 1270.820 1124.760 ;
        RECT 1271.050 1124.280 1271.370 1124.340 ;
        RECT 1270.680 1124.140 1271.370 1124.280 ;
        RECT 1271.050 1124.080 1271.370 1124.140 ;
        RECT 1271.050 1087.220 1271.370 1087.280 ;
        RECT 1270.680 1087.080 1271.370 1087.220 ;
        RECT 1270.680 1086.940 1270.820 1087.080 ;
        RECT 1271.050 1087.020 1271.370 1087.080 ;
        RECT 1270.590 1086.680 1270.910 1086.940 ;
        RECT 1270.590 966.180 1270.910 966.240 ;
        RECT 1271.510 966.180 1271.830 966.240 ;
        RECT 1270.590 966.040 1271.830 966.180 ;
        RECT 1270.590 965.980 1270.910 966.040 ;
        RECT 1271.510 965.980 1271.830 966.040 ;
        RECT 1271.510 917.900 1271.830 917.960 ;
        RECT 1271.140 917.760 1271.830 917.900 ;
        RECT 1271.140 917.620 1271.280 917.760 ;
        RECT 1271.510 917.700 1271.830 917.760 ;
        RECT 1271.050 917.360 1271.370 917.620 ;
        RECT 1270.605 886.620 1270.895 886.665 ;
        RECT 1271.050 886.620 1271.370 886.680 ;
        RECT 1270.605 886.480 1271.370 886.620 ;
        RECT 1270.605 886.435 1270.895 886.480 ;
        RECT 1271.050 886.420 1271.370 886.480 ;
        RECT 1270.590 862.820 1270.910 862.880 ;
        RECT 1270.395 862.680 1270.910 862.820 ;
        RECT 1270.590 862.620 1270.910 862.680 ;
        RECT 1270.590 821.000 1270.910 821.060 ;
        RECT 1271.510 821.000 1271.830 821.060 ;
        RECT 1270.590 820.860 1271.830 821.000 ;
        RECT 1270.590 820.800 1270.910 820.860 ;
        RECT 1271.510 820.800 1271.830 820.860 ;
        RECT 1271.050 724.440 1271.370 724.500 ;
        RECT 1271.510 724.440 1271.830 724.500 ;
        RECT 1271.050 724.300 1271.830 724.440 ;
        RECT 1271.050 724.240 1271.370 724.300 ;
        RECT 1271.510 724.240 1271.830 724.300 ;
        RECT 1271.050 627.880 1271.370 627.940 ;
        RECT 1271.510 627.880 1271.830 627.940 ;
        RECT 1271.050 627.740 1271.830 627.880 ;
        RECT 1271.050 627.680 1271.370 627.740 ;
        RECT 1271.510 627.680 1271.830 627.740 ;
        RECT 1270.590 579.600 1270.910 579.660 ;
        RECT 1270.395 579.460 1270.910 579.600 ;
        RECT 1270.590 579.400 1270.910 579.460 ;
        RECT 1270.590 544.920 1270.910 544.980 ;
        RECT 1270.395 544.780 1270.910 544.920 ;
        RECT 1270.590 544.720 1270.910 544.780 ;
        RECT 1270.590 531.320 1270.910 531.380 ;
        RECT 1271.050 531.320 1271.370 531.380 ;
        RECT 1270.590 531.180 1271.370 531.320 ;
        RECT 1270.590 531.120 1270.910 531.180 ;
        RECT 1271.050 531.120 1271.370 531.180 ;
        RECT 1270.590 434.420 1270.910 434.480 ;
        RECT 1270.395 434.280 1270.910 434.420 ;
        RECT 1270.590 434.220 1270.910 434.280 ;
        RECT 1270.590 386.480 1270.910 386.540 ;
        RECT 1270.395 386.340 1270.910 386.480 ;
        RECT 1270.590 386.280 1270.910 386.340 ;
        RECT 1270.590 241.780 1270.910 242.040 ;
        RECT 1270.680 241.640 1270.820 241.780 ;
        RECT 1271.050 241.640 1271.370 241.700 ;
        RECT 1270.680 241.500 1271.370 241.640 ;
        RECT 1271.050 241.440 1271.370 241.500 ;
        RECT 1270.130 144.740 1270.450 144.800 ;
        RECT 1271.050 144.740 1271.370 144.800 ;
        RECT 1270.130 144.600 1271.370 144.740 ;
        RECT 1270.130 144.540 1270.450 144.600 ;
        RECT 1271.050 144.540 1271.370 144.600 ;
        RECT 246.630 40.700 246.950 40.760 ;
        RECT 1270.130 40.700 1270.450 40.760 ;
        RECT 246.630 40.560 1270.450 40.700 ;
        RECT 246.630 40.500 246.950 40.560 ;
        RECT 1270.130 40.500 1270.450 40.560 ;
      LAYER via ;
        RECT 1270.620 1675.560 1270.880 1675.820 ;
        RECT 1275.220 1675.560 1275.480 1675.820 ;
        RECT 1271.080 1490.260 1271.340 1490.520 ;
        RECT 1272.460 1490.260 1272.720 1490.520 ;
        RECT 1271.080 1393.700 1271.340 1393.960 ;
        RECT 1272.460 1393.700 1272.720 1393.960 ;
        RECT 1271.080 1366.500 1271.340 1366.760 ;
        RECT 1270.620 1365.820 1270.880 1366.080 ;
        RECT 1270.160 1303.940 1270.420 1304.200 ;
        RECT 1271.080 1303.940 1271.340 1304.200 ;
        RECT 1270.160 1255.320 1270.420 1255.580 ;
        RECT 1271.080 1255.320 1271.340 1255.580 ;
        RECT 1270.160 1207.380 1270.420 1207.640 ;
        RECT 1271.080 1207.380 1271.340 1207.640 ;
        RECT 1270.620 1124.760 1270.880 1125.020 ;
        RECT 1271.080 1124.080 1271.340 1124.340 ;
        RECT 1271.080 1087.020 1271.340 1087.280 ;
        RECT 1270.620 1086.680 1270.880 1086.940 ;
        RECT 1270.620 965.980 1270.880 966.240 ;
        RECT 1271.540 965.980 1271.800 966.240 ;
        RECT 1271.540 917.700 1271.800 917.960 ;
        RECT 1271.080 917.360 1271.340 917.620 ;
        RECT 1271.080 886.420 1271.340 886.680 ;
        RECT 1270.620 862.620 1270.880 862.880 ;
        RECT 1270.620 820.800 1270.880 821.060 ;
        RECT 1271.540 820.800 1271.800 821.060 ;
        RECT 1271.080 724.240 1271.340 724.500 ;
        RECT 1271.540 724.240 1271.800 724.500 ;
        RECT 1271.080 627.680 1271.340 627.940 ;
        RECT 1271.540 627.680 1271.800 627.940 ;
        RECT 1270.620 579.400 1270.880 579.660 ;
        RECT 1270.620 544.720 1270.880 544.980 ;
        RECT 1270.620 531.120 1270.880 531.380 ;
        RECT 1271.080 531.120 1271.340 531.380 ;
        RECT 1270.620 434.220 1270.880 434.480 ;
        RECT 1270.620 386.280 1270.880 386.540 ;
        RECT 1270.620 241.780 1270.880 242.040 ;
        RECT 1271.080 241.440 1271.340 241.700 ;
        RECT 1270.160 144.540 1270.420 144.800 ;
        RECT 1271.080 144.540 1271.340 144.800 ;
        RECT 246.660 40.500 246.920 40.760 ;
        RECT 1270.160 40.500 1270.420 40.760 ;
      LAYER met2 ;
        RECT 1275.140 1700.000 1275.420 1702.400 ;
        RECT 1275.280 1675.850 1275.420 1700.000 ;
        RECT 1270.620 1675.530 1270.880 1675.850 ;
        RECT 1275.220 1675.530 1275.480 1675.850 ;
        RECT 1270.680 1655.530 1270.820 1675.530 ;
        RECT 1270.680 1655.390 1271.280 1655.530 ;
        RECT 1271.140 1606.570 1271.280 1655.390 ;
        RECT 1270.680 1606.430 1271.280 1606.570 ;
        RECT 1270.680 1593.650 1270.820 1606.430 ;
        RECT 1270.680 1593.510 1271.280 1593.650 ;
        RECT 1271.140 1490.550 1271.280 1593.510 ;
        RECT 1271.080 1490.230 1271.340 1490.550 ;
        RECT 1272.460 1490.230 1272.720 1490.550 ;
        RECT 1272.520 1483.605 1272.660 1490.230 ;
        RECT 1271.530 1483.235 1271.810 1483.605 ;
        RECT 1272.450 1483.235 1272.730 1483.605 ;
        RECT 1271.600 1440.650 1271.740 1483.235 ;
        RECT 1271.600 1440.510 1272.660 1440.650 ;
        RECT 1272.520 1393.990 1272.660 1440.510 ;
        RECT 1271.080 1393.670 1271.340 1393.990 ;
        RECT 1272.460 1393.670 1272.720 1393.990 ;
        RECT 1271.140 1366.790 1271.280 1393.670 ;
        RECT 1271.080 1366.470 1271.340 1366.790 ;
        RECT 1270.620 1365.790 1270.880 1366.110 ;
        RECT 1270.680 1328.450 1270.820 1365.790 ;
        RECT 1270.680 1328.310 1271.280 1328.450 ;
        RECT 1271.140 1304.230 1271.280 1328.310 ;
        RECT 1270.160 1303.910 1270.420 1304.230 ;
        RECT 1271.080 1303.910 1271.340 1304.230 ;
        RECT 1270.220 1297.285 1270.360 1303.910 ;
        RECT 1270.150 1296.915 1270.430 1297.285 ;
        RECT 1271.070 1296.915 1271.350 1297.285 ;
        RECT 1271.140 1255.610 1271.280 1296.915 ;
        RECT 1270.160 1255.290 1270.420 1255.610 ;
        RECT 1271.080 1255.290 1271.340 1255.610 ;
        RECT 1270.220 1207.670 1270.360 1255.290 ;
        RECT 1270.160 1207.525 1270.420 1207.670 ;
        RECT 1271.080 1207.525 1271.340 1207.670 ;
        RECT 1270.150 1207.155 1270.430 1207.525 ;
        RECT 1271.070 1207.155 1271.350 1207.525 ;
        RECT 1270.220 1182.930 1270.360 1207.155 ;
        RECT 1270.220 1182.790 1270.820 1182.930 ;
        RECT 1270.680 1125.050 1270.820 1182.790 ;
        RECT 1270.620 1124.730 1270.880 1125.050 ;
        RECT 1271.080 1124.050 1271.340 1124.370 ;
        RECT 1271.140 1087.310 1271.280 1124.050 ;
        RECT 1271.080 1086.990 1271.340 1087.310 ;
        RECT 1270.620 1086.650 1270.880 1086.970 ;
        RECT 1270.680 1062.570 1270.820 1086.650 ;
        RECT 1270.680 1062.430 1271.740 1062.570 ;
        RECT 1271.600 1027.890 1271.740 1062.430 ;
        RECT 1271.140 1027.750 1271.740 1027.890 ;
        RECT 1271.140 1014.290 1271.280 1027.750 ;
        RECT 1271.140 1014.150 1271.740 1014.290 ;
        RECT 1271.600 966.270 1271.740 1014.150 ;
        RECT 1270.620 966.125 1270.880 966.270 ;
        RECT 1271.540 966.125 1271.800 966.270 ;
        RECT 1270.610 965.755 1270.890 966.125 ;
        RECT 1271.530 965.755 1271.810 966.125 ;
        RECT 1271.600 917.990 1271.740 965.755 ;
        RECT 1271.540 917.670 1271.800 917.990 ;
        RECT 1271.080 917.330 1271.340 917.650 ;
        RECT 1271.140 886.710 1271.280 917.330 ;
        RECT 1271.080 886.390 1271.340 886.710 ;
        RECT 1270.620 862.590 1270.880 862.910 ;
        RECT 1270.680 821.090 1270.820 862.590 ;
        RECT 1270.620 820.770 1270.880 821.090 ;
        RECT 1271.540 820.770 1271.800 821.090 ;
        RECT 1271.600 773.005 1271.740 820.770 ;
        RECT 1271.530 772.635 1271.810 773.005 ;
        RECT 1271.530 771.955 1271.810 772.325 ;
        RECT 1271.600 737.530 1271.740 771.955 ;
        RECT 1271.140 737.390 1271.740 737.530 ;
        RECT 1271.140 724.530 1271.280 737.390 ;
        RECT 1271.080 724.210 1271.340 724.530 ;
        RECT 1271.540 724.210 1271.800 724.530 ;
        RECT 1271.600 676.445 1271.740 724.210 ;
        RECT 1270.610 676.075 1270.890 676.445 ;
        RECT 1271.530 676.075 1271.810 676.445 ;
        RECT 1270.680 651.850 1270.820 676.075 ;
        RECT 1270.680 651.710 1271.280 651.850 ;
        RECT 1271.140 627.970 1271.280 651.710 ;
        RECT 1271.080 627.650 1271.340 627.970 ;
        RECT 1271.540 627.650 1271.800 627.970 ;
        RECT 1271.600 579.885 1271.740 627.650 ;
        RECT 1270.610 579.515 1270.890 579.885 ;
        RECT 1271.530 579.515 1271.810 579.885 ;
        RECT 1270.620 579.370 1270.880 579.515 ;
        RECT 1270.620 544.690 1270.880 545.010 ;
        RECT 1270.680 531.490 1270.820 544.690 ;
        RECT 1270.680 531.410 1271.280 531.490 ;
        RECT 1270.620 531.350 1271.340 531.410 ;
        RECT 1270.620 531.090 1270.880 531.350 ;
        RECT 1271.080 531.090 1271.340 531.350 ;
        RECT 1270.680 434.510 1270.820 531.090 ;
        RECT 1270.620 434.190 1270.880 434.510 ;
        RECT 1270.620 386.250 1270.880 386.570 ;
        RECT 1270.680 242.070 1270.820 386.250 ;
        RECT 1270.620 241.750 1270.880 242.070 ;
        RECT 1271.080 241.410 1271.340 241.730 ;
        RECT 1271.140 207.810 1271.280 241.410 ;
        RECT 1271.140 207.670 1271.740 207.810 ;
        RECT 1271.600 196.930 1271.740 207.670 ;
        RECT 1271.140 196.790 1271.740 196.930 ;
        RECT 1271.140 144.830 1271.280 196.790 ;
        RECT 1270.160 144.510 1270.420 144.830 ;
        RECT 1271.080 144.510 1271.340 144.830 ;
        RECT 1270.220 96.970 1270.360 144.510 ;
        RECT 1270.220 96.830 1270.820 96.970 ;
        RECT 1270.680 48.520 1270.820 96.830 ;
        RECT 1270.220 48.380 1270.820 48.520 ;
        RECT 1270.220 40.790 1270.360 48.380 ;
        RECT 246.660 40.470 246.920 40.790 ;
        RECT 1270.160 40.470 1270.420 40.790 ;
        RECT 246.720 2.400 246.860 40.470 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 1271.530 1483.280 1271.810 1483.560 ;
        RECT 1272.450 1483.280 1272.730 1483.560 ;
        RECT 1270.150 1296.960 1270.430 1297.240 ;
        RECT 1271.070 1296.960 1271.350 1297.240 ;
        RECT 1270.150 1207.200 1270.430 1207.480 ;
        RECT 1271.070 1207.200 1271.350 1207.480 ;
        RECT 1270.610 965.800 1270.890 966.080 ;
        RECT 1271.530 965.800 1271.810 966.080 ;
        RECT 1271.530 772.680 1271.810 772.960 ;
        RECT 1271.530 772.000 1271.810 772.280 ;
        RECT 1270.610 676.120 1270.890 676.400 ;
        RECT 1271.530 676.120 1271.810 676.400 ;
        RECT 1270.610 579.560 1270.890 579.840 ;
        RECT 1271.530 579.560 1271.810 579.840 ;
      LAYER met3 ;
        RECT 1271.505 1483.570 1271.835 1483.585 ;
        RECT 1272.425 1483.570 1272.755 1483.585 ;
        RECT 1271.505 1483.270 1272.755 1483.570 ;
        RECT 1271.505 1483.255 1271.835 1483.270 ;
        RECT 1272.425 1483.255 1272.755 1483.270 ;
        RECT 1270.125 1297.250 1270.455 1297.265 ;
        RECT 1271.045 1297.250 1271.375 1297.265 ;
        RECT 1270.125 1296.950 1271.375 1297.250 ;
        RECT 1270.125 1296.935 1270.455 1296.950 ;
        RECT 1271.045 1296.935 1271.375 1296.950 ;
        RECT 1270.125 1207.490 1270.455 1207.505 ;
        RECT 1271.045 1207.490 1271.375 1207.505 ;
        RECT 1270.125 1207.190 1271.375 1207.490 ;
        RECT 1270.125 1207.175 1270.455 1207.190 ;
        RECT 1271.045 1207.175 1271.375 1207.190 ;
        RECT 1270.585 966.090 1270.915 966.105 ;
        RECT 1271.505 966.090 1271.835 966.105 ;
        RECT 1270.585 965.790 1271.835 966.090 ;
        RECT 1270.585 965.775 1270.915 965.790 ;
        RECT 1271.505 965.775 1271.835 965.790 ;
        RECT 1271.505 772.970 1271.835 772.985 ;
        RECT 1270.830 772.670 1271.835 772.970 ;
        RECT 1270.830 772.290 1271.130 772.670 ;
        RECT 1271.505 772.655 1271.835 772.670 ;
        RECT 1271.505 772.290 1271.835 772.305 ;
        RECT 1270.830 771.990 1271.835 772.290 ;
        RECT 1271.505 771.975 1271.835 771.990 ;
        RECT 1270.585 676.410 1270.915 676.425 ;
        RECT 1271.505 676.410 1271.835 676.425 ;
        RECT 1270.585 676.110 1271.835 676.410 ;
        RECT 1270.585 676.095 1270.915 676.110 ;
        RECT 1271.505 676.095 1271.835 676.110 ;
        RECT 1270.585 579.850 1270.915 579.865 ;
        RECT 1271.505 579.850 1271.835 579.865 ;
        RECT 1270.585 579.550 1271.835 579.850 ;
        RECT 1270.585 579.535 1270.915 579.550 ;
        RECT 1271.505 579.535 1271.835 579.550 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 41.040 264.430 41.100 ;
        RECT 1283.930 41.040 1284.250 41.100 ;
        RECT 264.110 40.900 1284.250 41.040 ;
        RECT 264.110 40.840 264.430 40.900 ;
        RECT 1283.930 40.840 1284.250 40.900 ;
      LAYER via ;
        RECT 264.140 40.840 264.400 41.100 ;
        RECT 1283.960 40.840 1284.220 41.100 ;
      LAYER met2 ;
        RECT 1284.340 1700.410 1284.620 1702.400 ;
        RECT 1284.020 1700.270 1284.620 1700.410 ;
        RECT 1284.020 41.130 1284.160 1700.270 ;
        RECT 1284.340 1700.000 1284.620 1700.270 ;
        RECT 264.140 40.810 264.400 41.130 ;
        RECT 1283.960 40.810 1284.220 41.130 ;
        RECT 264.200 2.400 264.340 40.810 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 41.380 282.370 41.440 ;
        RECT 1291.750 41.380 1292.070 41.440 ;
        RECT 282.050 41.240 1292.070 41.380 ;
        RECT 282.050 41.180 282.370 41.240 ;
        RECT 1291.750 41.180 1292.070 41.240 ;
      LAYER via ;
        RECT 282.080 41.180 282.340 41.440 ;
        RECT 1291.780 41.180 1292.040 41.440 ;
      LAYER met2 ;
        RECT 1293.540 1700.410 1293.820 1702.400 ;
        RECT 1291.840 1700.270 1293.820 1700.410 ;
        RECT 1291.840 41.470 1291.980 1700.270 ;
        RECT 1293.540 1700.000 1293.820 1700.270 ;
        RECT 282.080 41.150 282.340 41.470 ;
        RECT 1291.780 41.150 1292.040 41.470 ;
        RECT 282.140 2.400 282.280 41.150 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1298.265 1594.005 1298.435 1608.115 ;
        RECT 1298.265 1413.805 1298.435 1448.995 ;
        RECT 1298.265 1110.865 1298.435 1158.975 ;
        RECT 1298.265 772.905 1298.435 821.015 ;
        RECT 1298.265 386.325 1298.435 434.435 ;
        RECT 1298.265 241.485 1298.435 298.775 ;
        RECT 1299.185 89.845 1299.355 137.955 ;
      LAYER mcon ;
        RECT 1298.265 1607.945 1298.435 1608.115 ;
        RECT 1298.265 1448.825 1298.435 1448.995 ;
        RECT 1298.265 1158.805 1298.435 1158.975 ;
        RECT 1298.265 820.845 1298.435 821.015 ;
        RECT 1298.265 434.265 1298.435 434.435 ;
        RECT 1298.265 298.605 1298.435 298.775 ;
        RECT 1299.185 137.785 1299.355 137.955 ;
      LAYER met1 ;
        RECT 1298.190 1678.140 1298.510 1678.200 ;
        RECT 1301.410 1678.140 1301.730 1678.200 ;
        RECT 1298.190 1678.000 1301.730 1678.140 ;
        RECT 1298.190 1677.940 1298.510 1678.000 ;
        RECT 1301.410 1677.940 1301.730 1678.000 ;
        RECT 1298.205 1608.100 1298.495 1608.145 ;
        RECT 1298.650 1608.100 1298.970 1608.160 ;
        RECT 1298.205 1607.960 1298.970 1608.100 ;
        RECT 1298.205 1607.915 1298.495 1607.960 ;
        RECT 1298.650 1607.900 1298.970 1607.960 ;
        RECT 1298.190 1594.160 1298.510 1594.220 ;
        RECT 1297.995 1594.020 1298.510 1594.160 ;
        RECT 1298.190 1593.960 1298.510 1594.020 ;
        RECT 1298.190 1448.980 1298.510 1449.040 ;
        RECT 1297.995 1448.840 1298.510 1448.980 ;
        RECT 1298.190 1448.780 1298.510 1448.840 ;
        RECT 1298.205 1413.960 1298.495 1414.005 ;
        RECT 1298.650 1413.960 1298.970 1414.020 ;
        RECT 1298.205 1413.820 1298.970 1413.960 ;
        RECT 1298.205 1413.775 1298.495 1413.820 ;
        RECT 1298.650 1413.760 1298.970 1413.820 ;
        RECT 1296.810 1338.820 1297.130 1338.880 ;
        RECT 1297.730 1338.820 1298.050 1338.880 ;
        RECT 1296.810 1338.680 1298.050 1338.820 ;
        RECT 1296.810 1338.620 1297.130 1338.680 ;
        RECT 1297.730 1338.620 1298.050 1338.680 ;
        RECT 1297.730 1249.060 1298.050 1249.120 ;
        RECT 1298.650 1249.060 1298.970 1249.120 ;
        RECT 1297.730 1248.920 1298.970 1249.060 ;
        RECT 1297.730 1248.860 1298.050 1248.920 ;
        RECT 1298.650 1248.860 1298.970 1248.920 ;
        RECT 1297.730 1207.580 1298.050 1207.640 ;
        RECT 1298.650 1207.580 1298.970 1207.640 ;
        RECT 1297.730 1207.440 1298.970 1207.580 ;
        RECT 1297.730 1207.380 1298.050 1207.440 ;
        RECT 1298.650 1207.380 1298.970 1207.440 ;
        RECT 1298.190 1158.960 1298.510 1159.020 ;
        RECT 1297.995 1158.820 1298.510 1158.960 ;
        RECT 1298.190 1158.760 1298.510 1158.820 ;
        RECT 1298.205 1111.020 1298.495 1111.065 ;
        RECT 1298.650 1111.020 1298.970 1111.080 ;
        RECT 1298.205 1110.880 1298.970 1111.020 ;
        RECT 1298.205 1110.835 1298.495 1110.880 ;
        RECT 1298.650 1110.820 1298.970 1110.880 ;
        RECT 1298.650 1087.220 1298.970 1087.280 ;
        RECT 1298.280 1087.080 1298.970 1087.220 ;
        RECT 1298.280 1086.940 1298.420 1087.080 ;
        RECT 1298.650 1087.020 1298.970 1087.080 ;
        RECT 1298.190 1086.680 1298.510 1086.940 ;
        RECT 1298.190 1028.200 1298.510 1028.460 ;
        RECT 1298.280 1027.720 1298.420 1028.200 ;
        RECT 1298.650 1027.720 1298.970 1027.780 ;
        RECT 1298.280 1027.580 1298.970 1027.720 ;
        RECT 1298.650 1027.520 1298.970 1027.580 ;
        RECT 1298.650 966.180 1298.970 966.240 ;
        RECT 1298.280 966.040 1298.970 966.180 ;
        RECT 1298.280 965.900 1298.420 966.040 ;
        RECT 1298.650 965.980 1298.970 966.040 ;
        RECT 1298.190 965.640 1298.510 965.900 ;
        RECT 1298.650 910.760 1298.970 910.820 ;
        RECT 1299.570 910.760 1299.890 910.820 ;
        RECT 1298.650 910.620 1299.890 910.760 ;
        RECT 1298.650 910.560 1298.970 910.620 ;
        RECT 1299.570 910.560 1299.890 910.620 ;
        RECT 1298.190 821.000 1298.510 821.060 ;
        RECT 1297.995 820.860 1298.510 821.000 ;
        RECT 1298.190 820.800 1298.510 820.860 ;
        RECT 1298.190 773.060 1298.510 773.120 ;
        RECT 1297.995 772.920 1298.510 773.060 ;
        RECT 1298.190 772.860 1298.510 772.920 ;
        RECT 1298.190 738.180 1298.510 738.440 ;
        RECT 1298.280 738.040 1298.420 738.180 ;
        RECT 1298.650 738.040 1298.970 738.100 ;
        RECT 1298.280 737.900 1298.970 738.040 ;
        RECT 1298.650 737.840 1298.970 737.900 ;
        RECT 1298.650 724.440 1298.970 724.500 ;
        RECT 1299.110 724.440 1299.430 724.500 ;
        RECT 1298.650 724.300 1299.430 724.440 ;
        RECT 1298.650 724.240 1298.970 724.300 ;
        RECT 1299.110 724.240 1299.430 724.300 ;
        RECT 1298.190 676.160 1298.510 676.220 ;
        RECT 1299.110 676.160 1299.430 676.220 ;
        RECT 1298.190 676.020 1299.430 676.160 ;
        RECT 1298.190 675.960 1298.510 676.020 ;
        RECT 1299.110 675.960 1299.430 676.020 ;
        RECT 1298.650 627.880 1298.970 627.940 ;
        RECT 1299.110 627.880 1299.430 627.940 ;
        RECT 1298.650 627.740 1299.430 627.880 ;
        RECT 1298.650 627.680 1298.970 627.740 ;
        RECT 1299.110 627.680 1299.430 627.740 ;
        RECT 1298.190 579.600 1298.510 579.660 ;
        RECT 1299.110 579.600 1299.430 579.660 ;
        RECT 1298.190 579.460 1299.430 579.600 ;
        RECT 1298.190 579.400 1298.510 579.460 ;
        RECT 1299.110 579.400 1299.430 579.460 ;
        RECT 1298.190 434.420 1298.510 434.480 ;
        RECT 1297.995 434.280 1298.510 434.420 ;
        RECT 1298.190 434.220 1298.510 434.280 ;
        RECT 1298.190 386.480 1298.510 386.540 ;
        RECT 1297.995 386.340 1298.510 386.480 ;
        RECT 1298.190 386.280 1298.510 386.340 ;
        RECT 1298.190 298.760 1298.510 298.820 ;
        RECT 1297.995 298.620 1298.510 298.760 ;
        RECT 1298.190 298.560 1298.510 298.620 ;
        RECT 1298.205 241.640 1298.495 241.685 ;
        RECT 1298.650 241.640 1298.970 241.700 ;
        RECT 1298.205 241.500 1298.970 241.640 ;
        RECT 1298.205 241.455 1298.495 241.500 ;
        RECT 1298.650 241.440 1298.970 241.500 ;
        RECT 1298.650 144.740 1298.970 144.800 ;
        RECT 1299.110 144.740 1299.430 144.800 ;
        RECT 1298.650 144.600 1299.430 144.740 ;
        RECT 1298.650 144.540 1298.970 144.600 ;
        RECT 1299.110 144.540 1299.430 144.600 ;
        RECT 1299.110 137.940 1299.430 138.000 ;
        RECT 1298.915 137.800 1299.430 137.940 ;
        RECT 1299.110 137.740 1299.430 137.800 ;
        RECT 1299.110 90.000 1299.430 90.060 ;
        RECT 1298.915 89.860 1299.430 90.000 ;
        RECT 1299.110 89.800 1299.430 89.860 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 1298.220 1677.940 1298.480 1678.200 ;
        RECT 1301.440 1677.940 1301.700 1678.200 ;
        RECT 1298.680 1607.900 1298.940 1608.160 ;
        RECT 1298.220 1593.960 1298.480 1594.220 ;
        RECT 1298.220 1448.780 1298.480 1449.040 ;
        RECT 1298.680 1413.760 1298.940 1414.020 ;
        RECT 1296.840 1338.620 1297.100 1338.880 ;
        RECT 1297.760 1338.620 1298.020 1338.880 ;
        RECT 1297.760 1248.860 1298.020 1249.120 ;
        RECT 1298.680 1248.860 1298.940 1249.120 ;
        RECT 1297.760 1207.380 1298.020 1207.640 ;
        RECT 1298.680 1207.380 1298.940 1207.640 ;
        RECT 1298.220 1158.760 1298.480 1159.020 ;
        RECT 1298.680 1110.820 1298.940 1111.080 ;
        RECT 1298.680 1087.020 1298.940 1087.280 ;
        RECT 1298.220 1086.680 1298.480 1086.940 ;
        RECT 1298.220 1028.200 1298.480 1028.460 ;
        RECT 1298.680 1027.520 1298.940 1027.780 ;
        RECT 1298.680 965.980 1298.940 966.240 ;
        RECT 1298.220 965.640 1298.480 965.900 ;
        RECT 1298.680 910.560 1298.940 910.820 ;
        RECT 1299.600 910.560 1299.860 910.820 ;
        RECT 1298.220 820.800 1298.480 821.060 ;
        RECT 1298.220 772.860 1298.480 773.120 ;
        RECT 1298.220 738.180 1298.480 738.440 ;
        RECT 1298.680 737.840 1298.940 738.100 ;
        RECT 1298.680 724.240 1298.940 724.500 ;
        RECT 1299.140 724.240 1299.400 724.500 ;
        RECT 1298.220 675.960 1298.480 676.220 ;
        RECT 1299.140 675.960 1299.400 676.220 ;
        RECT 1298.680 627.680 1298.940 627.940 ;
        RECT 1299.140 627.680 1299.400 627.940 ;
        RECT 1298.220 579.400 1298.480 579.660 ;
        RECT 1299.140 579.400 1299.400 579.660 ;
        RECT 1298.220 434.220 1298.480 434.480 ;
        RECT 1298.220 386.280 1298.480 386.540 ;
        RECT 1298.220 298.560 1298.480 298.820 ;
        RECT 1298.680 241.440 1298.940 241.700 ;
        RECT 1298.680 144.540 1298.940 144.800 ;
        RECT 1299.140 144.540 1299.400 144.800 ;
        RECT 1299.140 137.740 1299.400 138.000 ;
        RECT 1299.140 89.800 1299.400 90.060 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 1302.740 1700.410 1303.020 1702.400 ;
        RECT 1301.500 1700.270 1303.020 1700.410 ;
        RECT 1301.500 1678.230 1301.640 1700.270 ;
        RECT 1302.740 1700.000 1303.020 1700.270 ;
        RECT 1298.220 1677.910 1298.480 1678.230 ;
        RECT 1301.440 1677.910 1301.700 1678.230 ;
        RECT 1298.280 1655.530 1298.420 1677.910 ;
        RECT 1298.280 1655.390 1298.880 1655.530 ;
        RECT 1298.740 1608.190 1298.880 1655.390 ;
        RECT 1298.680 1607.870 1298.940 1608.190 ;
        RECT 1298.220 1593.930 1298.480 1594.250 ;
        RECT 1298.280 1593.650 1298.420 1593.930 ;
        RECT 1298.280 1593.510 1298.880 1593.650 ;
        RECT 1298.740 1463.090 1298.880 1593.510 ;
        RECT 1298.280 1462.950 1298.880 1463.090 ;
        RECT 1298.280 1449.070 1298.420 1462.950 ;
        RECT 1298.220 1448.750 1298.480 1449.070 ;
        RECT 1298.680 1413.730 1298.940 1414.050 ;
        RECT 1298.740 1387.045 1298.880 1413.730 ;
        RECT 1296.830 1386.675 1297.110 1387.045 ;
        RECT 1298.670 1386.675 1298.950 1387.045 ;
        RECT 1296.900 1338.910 1297.040 1386.675 ;
        RECT 1296.840 1338.590 1297.100 1338.910 ;
        RECT 1297.760 1338.590 1298.020 1338.910 ;
        RECT 1297.820 1297.285 1297.960 1338.590 ;
        RECT 1297.750 1296.915 1298.030 1297.285 ;
        RECT 1298.670 1296.915 1298.950 1297.285 ;
        RECT 1298.740 1249.150 1298.880 1296.915 ;
        RECT 1297.760 1248.830 1298.020 1249.150 ;
        RECT 1298.680 1248.830 1298.940 1249.150 ;
        RECT 1297.820 1207.670 1297.960 1248.830 ;
        RECT 1297.760 1207.525 1298.020 1207.670 ;
        RECT 1298.680 1207.525 1298.940 1207.670 ;
        RECT 1297.750 1207.155 1298.030 1207.525 ;
        RECT 1298.670 1207.155 1298.950 1207.525 ;
        RECT 1297.820 1182.930 1297.960 1207.155 ;
        RECT 1297.820 1182.790 1298.420 1182.930 ;
        RECT 1298.280 1159.050 1298.420 1182.790 ;
        RECT 1298.220 1158.730 1298.480 1159.050 ;
        RECT 1298.680 1110.790 1298.940 1111.110 ;
        RECT 1298.740 1087.310 1298.880 1110.790 ;
        RECT 1298.680 1086.990 1298.940 1087.310 ;
        RECT 1298.220 1086.650 1298.480 1086.970 ;
        RECT 1298.280 1028.490 1298.420 1086.650 ;
        RECT 1298.220 1028.170 1298.480 1028.490 ;
        RECT 1298.680 1027.490 1298.940 1027.810 ;
        RECT 1298.740 966.270 1298.880 1027.490 ;
        RECT 1298.680 965.950 1298.940 966.270 ;
        RECT 1298.220 965.610 1298.480 965.930 ;
        RECT 1298.280 911.725 1298.420 965.610 ;
        RECT 1298.210 911.355 1298.490 911.725 ;
        RECT 1298.670 910.675 1298.950 911.045 ;
        RECT 1298.680 910.530 1298.940 910.675 ;
        RECT 1299.600 910.530 1299.860 910.850 ;
        RECT 1299.660 862.765 1299.800 910.530 ;
        RECT 1298.210 862.395 1298.490 862.765 ;
        RECT 1299.590 862.395 1299.870 862.765 ;
        RECT 1298.280 821.090 1298.420 862.395 ;
        RECT 1298.220 820.770 1298.480 821.090 ;
        RECT 1298.220 772.830 1298.480 773.150 ;
        RECT 1298.280 738.470 1298.420 772.830 ;
        RECT 1298.220 738.150 1298.480 738.470 ;
        RECT 1298.680 737.810 1298.940 738.130 ;
        RECT 1298.740 724.530 1298.880 737.810 ;
        RECT 1298.680 724.210 1298.940 724.530 ;
        RECT 1299.140 724.210 1299.400 724.530 ;
        RECT 1299.200 676.445 1299.340 724.210 ;
        RECT 1298.210 676.075 1298.490 676.445 ;
        RECT 1299.130 676.075 1299.410 676.445 ;
        RECT 1298.220 675.930 1298.480 676.075 ;
        RECT 1299.140 675.930 1299.400 676.075 ;
        RECT 1299.200 628.050 1299.340 675.930 ;
        RECT 1298.740 627.970 1299.340 628.050 ;
        RECT 1298.680 627.910 1299.400 627.970 ;
        RECT 1298.680 627.650 1298.940 627.910 ;
        RECT 1299.140 627.650 1299.400 627.910 ;
        RECT 1299.200 579.885 1299.340 627.650 ;
        RECT 1298.210 579.515 1298.490 579.885 ;
        RECT 1299.130 579.515 1299.410 579.885 ;
        RECT 1298.220 579.370 1298.480 579.515 ;
        RECT 1299.140 579.370 1299.400 579.515 ;
        RECT 1299.200 483.325 1299.340 579.370 ;
        RECT 1298.210 482.955 1298.490 483.325 ;
        RECT 1299.130 482.955 1299.410 483.325 ;
        RECT 1298.280 434.510 1298.420 482.955 ;
        RECT 1298.220 434.190 1298.480 434.510 ;
        RECT 1298.220 386.250 1298.480 386.570 ;
        RECT 1298.280 298.850 1298.420 386.250 ;
        RECT 1298.220 298.530 1298.480 298.850 ;
        RECT 1298.680 241.410 1298.940 241.730 ;
        RECT 1298.740 144.830 1298.880 241.410 ;
        RECT 1298.680 144.510 1298.940 144.830 ;
        RECT 1299.140 144.510 1299.400 144.830 ;
        RECT 1299.200 138.030 1299.340 144.510 ;
        RECT 1299.140 137.710 1299.400 138.030 ;
        RECT 1299.140 89.770 1299.400 90.090 ;
        RECT 1299.200 51.525 1299.340 89.770 ;
        RECT 303.230 51.155 303.510 51.525 ;
        RECT 1299.130 51.155 1299.410 51.525 ;
        RECT 303.300 16.990 303.440 51.155 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
      LAYER via2 ;
        RECT 1296.830 1386.720 1297.110 1387.000 ;
        RECT 1298.670 1386.720 1298.950 1387.000 ;
        RECT 1297.750 1296.960 1298.030 1297.240 ;
        RECT 1298.670 1296.960 1298.950 1297.240 ;
        RECT 1297.750 1207.200 1298.030 1207.480 ;
        RECT 1298.670 1207.200 1298.950 1207.480 ;
        RECT 1298.210 911.400 1298.490 911.680 ;
        RECT 1298.670 910.720 1298.950 911.000 ;
        RECT 1298.210 862.440 1298.490 862.720 ;
        RECT 1299.590 862.440 1299.870 862.720 ;
        RECT 1298.210 676.120 1298.490 676.400 ;
        RECT 1299.130 676.120 1299.410 676.400 ;
        RECT 1298.210 579.560 1298.490 579.840 ;
        RECT 1299.130 579.560 1299.410 579.840 ;
        RECT 1298.210 483.000 1298.490 483.280 ;
        RECT 1299.130 483.000 1299.410 483.280 ;
        RECT 303.230 51.200 303.510 51.480 ;
        RECT 1299.130 51.200 1299.410 51.480 ;
      LAYER met3 ;
        RECT 1296.805 1387.010 1297.135 1387.025 ;
        RECT 1298.645 1387.010 1298.975 1387.025 ;
        RECT 1296.805 1386.710 1298.975 1387.010 ;
        RECT 1296.805 1386.695 1297.135 1386.710 ;
        RECT 1298.645 1386.695 1298.975 1386.710 ;
        RECT 1297.725 1297.250 1298.055 1297.265 ;
        RECT 1298.645 1297.250 1298.975 1297.265 ;
        RECT 1297.725 1296.950 1298.975 1297.250 ;
        RECT 1297.725 1296.935 1298.055 1296.950 ;
        RECT 1298.645 1296.935 1298.975 1296.950 ;
        RECT 1297.725 1207.490 1298.055 1207.505 ;
        RECT 1298.645 1207.490 1298.975 1207.505 ;
        RECT 1297.725 1207.190 1298.975 1207.490 ;
        RECT 1297.725 1207.175 1298.055 1207.190 ;
        RECT 1298.645 1207.175 1298.975 1207.190 ;
        RECT 1298.185 911.690 1298.515 911.705 ;
        RECT 1298.185 911.375 1298.730 911.690 ;
        RECT 1298.430 911.025 1298.730 911.375 ;
        RECT 1298.430 910.710 1298.975 911.025 ;
        RECT 1298.645 910.695 1298.975 910.710 ;
        RECT 1298.185 862.730 1298.515 862.745 ;
        RECT 1299.565 862.730 1299.895 862.745 ;
        RECT 1298.185 862.430 1299.895 862.730 ;
        RECT 1298.185 862.415 1298.515 862.430 ;
        RECT 1299.565 862.415 1299.895 862.430 ;
        RECT 1298.185 676.410 1298.515 676.425 ;
        RECT 1299.105 676.410 1299.435 676.425 ;
        RECT 1298.185 676.110 1299.435 676.410 ;
        RECT 1298.185 676.095 1298.515 676.110 ;
        RECT 1299.105 676.095 1299.435 676.110 ;
        RECT 1298.185 579.850 1298.515 579.865 ;
        RECT 1299.105 579.850 1299.435 579.865 ;
        RECT 1298.185 579.550 1299.435 579.850 ;
        RECT 1298.185 579.535 1298.515 579.550 ;
        RECT 1299.105 579.535 1299.435 579.550 ;
        RECT 1298.185 483.290 1298.515 483.305 ;
        RECT 1299.105 483.290 1299.435 483.305 ;
        RECT 1298.185 482.990 1299.435 483.290 ;
        RECT 1298.185 482.975 1298.515 482.990 ;
        RECT 1299.105 482.975 1299.435 482.990 ;
        RECT 303.205 51.490 303.535 51.505 ;
        RECT 1299.105 51.490 1299.435 51.505 ;
        RECT 303.205 51.190 1299.435 51.490 ;
        RECT 303.205 51.175 303.535 51.190 ;
        RECT 1299.105 51.175 1299.435 51.190 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.910 51.580 324.230 51.640 ;
        RECT 1311.530 51.580 1311.850 51.640 ;
        RECT 323.910 51.440 1311.850 51.580 ;
        RECT 323.910 51.380 324.230 51.440 ;
        RECT 1311.530 51.380 1311.850 51.440 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 323.910 16.900 324.230 16.960 ;
        RECT 317.930 16.760 324.230 16.900 ;
        RECT 317.930 16.700 318.250 16.760 ;
        RECT 323.910 16.700 324.230 16.760 ;
      LAYER via ;
        RECT 323.940 51.380 324.200 51.640 ;
        RECT 1311.560 51.380 1311.820 51.640 ;
        RECT 317.960 16.700 318.220 16.960 ;
        RECT 323.940 16.700 324.200 16.960 ;
      LAYER met2 ;
        RECT 1311.940 1700.410 1312.220 1702.400 ;
        RECT 1311.620 1700.270 1312.220 1700.410 ;
        RECT 1311.620 51.670 1311.760 1700.270 ;
        RECT 1311.940 1700.000 1312.220 1700.270 ;
        RECT 323.940 51.350 324.200 51.670 ;
        RECT 1311.560 51.350 1311.820 51.670 ;
        RECT 324.000 16.990 324.140 51.350 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 323.940 16.670 324.200 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 335.870 26.420 336.190 26.480 ;
        RECT 1318.890 26.420 1319.210 26.480 ;
        RECT 335.870 26.280 1319.210 26.420 ;
        RECT 335.870 26.220 336.190 26.280 ;
        RECT 1318.890 26.220 1319.210 26.280 ;
      LAYER via ;
        RECT 335.900 26.220 336.160 26.480 ;
        RECT 1318.920 26.220 1319.180 26.480 ;
      LAYER met2 ;
        RECT 1321.140 1700.410 1321.420 1702.400 ;
        RECT 1318.980 1700.270 1321.420 1700.410 ;
        RECT 1318.980 26.510 1319.120 1700.270 ;
        RECT 1321.140 1700.000 1321.420 1700.270 ;
        RECT 335.900 26.190 336.160 26.510 ;
        RECT 1318.920 26.190 1319.180 26.510 ;
        RECT 335.960 2.400 336.100 26.190 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1326.325 1442.025 1326.495 1490.475 ;
        RECT 1325.865 1013.965 1326.035 1048.815 ;
        RECT 1326.325 758.965 1326.495 807.075 ;
        RECT 1326.785 622.965 1326.955 662.235 ;
        RECT 1325.865 427.805 1326.035 475.915 ;
      LAYER mcon ;
        RECT 1326.325 1490.305 1326.495 1490.475 ;
        RECT 1325.865 1048.645 1326.035 1048.815 ;
        RECT 1326.325 806.905 1326.495 807.075 ;
        RECT 1326.785 662.065 1326.955 662.235 ;
        RECT 1325.865 475.745 1326.035 475.915 ;
      LAYER met1 ;
        RECT 1326.250 1642.440 1326.570 1642.500 ;
        RECT 1327.630 1642.440 1327.950 1642.500 ;
        RECT 1326.250 1642.300 1327.950 1642.440 ;
        RECT 1326.250 1642.240 1326.570 1642.300 ;
        RECT 1327.630 1642.240 1327.950 1642.300 ;
        RECT 1325.790 1497.600 1326.110 1497.660 ;
        RECT 1326.250 1497.600 1326.570 1497.660 ;
        RECT 1325.790 1497.460 1326.570 1497.600 ;
        RECT 1325.790 1497.400 1326.110 1497.460 ;
        RECT 1326.250 1497.400 1326.570 1497.460 ;
        RECT 1326.250 1490.460 1326.570 1490.520 ;
        RECT 1326.055 1490.320 1326.570 1490.460 ;
        RECT 1326.250 1490.260 1326.570 1490.320 ;
        RECT 1326.250 1442.180 1326.570 1442.240 ;
        RECT 1326.055 1442.040 1326.570 1442.180 ;
        RECT 1326.250 1441.980 1326.570 1442.040 ;
        RECT 1325.790 1400.700 1326.110 1400.760 ;
        RECT 1326.250 1400.700 1326.570 1400.760 ;
        RECT 1325.790 1400.560 1326.570 1400.700 ;
        RECT 1325.790 1400.500 1326.110 1400.560 ;
        RECT 1326.250 1400.500 1326.570 1400.560 ;
        RECT 1325.790 1152.840 1326.110 1152.900 ;
        RECT 1326.250 1152.840 1326.570 1152.900 ;
        RECT 1325.790 1152.700 1326.570 1152.840 ;
        RECT 1325.790 1152.640 1326.110 1152.700 ;
        RECT 1326.250 1152.640 1326.570 1152.700 ;
        RECT 1325.790 1124.280 1326.110 1124.340 ;
        RECT 1326.710 1124.280 1327.030 1124.340 ;
        RECT 1325.790 1124.140 1327.030 1124.280 ;
        RECT 1325.790 1124.080 1326.110 1124.140 ;
        RECT 1326.710 1124.080 1327.030 1124.140 ;
        RECT 1325.790 1048.800 1326.110 1048.860 ;
        RECT 1325.595 1048.660 1326.110 1048.800 ;
        RECT 1325.790 1048.600 1326.110 1048.660 ;
        RECT 1325.805 1014.120 1326.095 1014.165 ;
        RECT 1326.250 1014.120 1326.570 1014.180 ;
        RECT 1325.805 1013.980 1326.570 1014.120 ;
        RECT 1325.805 1013.935 1326.095 1013.980 ;
        RECT 1326.250 1013.920 1326.570 1013.980 ;
        RECT 1325.790 966.520 1326.110 966.580 ;
        RECT 1326.710 966.520 1327.030 966.580 ;
        RECT 1325.790 966.380 1327.030 966.520 ;
        RECT 1325.790 966.320 1326.110 966.380 ;
        RECT 1326.710 966.320 1327.030 966.380 ;
        RECT 1326.250 870.100 1326.570 870.360 ;
        RECT 1326.340 869.680 1326.480 870.100 ;
        RECT 1326.250 869.420 1326.570 869.680 ;
        RECT 1326.250 807.060 1326.570 807.120 ;
        RECT 1326.055 806.920 1326.570 807.060 ;
        RECT 1326.250 806.860 1326.570 806.920 ;
        RECT 1326.250 759.120 1326.570 759.180 ;
        RECT 1326.055 758.980 1326.570 759.120 ;
        RECT 1326.250 758.920 1326.570 758.980 ;
        RECT 1326.710 662.220 1327.030 662.280 ;
        RECT 1326.515 662.080 1327.030 662.220 ;
        RECT 1326.710 662.020 1327.030 662.080 ;
        RECT 1326.710 623.120 1327.030 623.180 ;
        RECT 1326.515 622.980 1327.030 623.120 ;
        RECT 1326.710 622.920 1327.030 622.980 ;
        RECT 1325.790 579.600 1326.110 579.660 ;
        RECT 1326.250 579.600 1326.570 579.660 ;
        RECT 1325.790 579.460 1326.570 579.600 ;
        RECT 1325.790 579.400 1326.110 579.460 ;
        RECT 1326.250 579.400 1326.570 579.460 ;
        RECT 1325.790 475.900 1326.110 475.960 ;
        RECT 1325.595 475.760 1326.110 475.900 ;
        RECT 1325.790 475.700 1326.110 475.760 ;
        RECT 1325.790 427.960 1326.110 428.020 ;
        RECT 1325.595 427.820 1326.110 427.960 ;
        RECT 1325.790 427.760 1326.110 427.820 ;
        RECT 1325.790 241.640 1326.110 241.700 ;
        RECT 1326.710 241.640 1327.030 241.700 ;
        RECT 1325.790 241.500 1327.030 241.640 ;
        RECT 1325.790 241.440 1326.110 241.500 ;
        RECT 1326.710 241.440 1327.030 241.500 ;
        RECT 1325.790 144.740 1326.110 144.800 ;
        RECT 1326.250 144.740 1326.570 144.800 ;
        RECT 1325.790 144.600 1326.570 144.740 ;
        RECT 1325.790 144.540 1326.110 144.600 ;
        RECT 1326.250 144.540 1326.570 144.600 ;
        RECT 358.410 72.660 358.730 72.720 ;
        RECT 1325.790 72.660 1326.110 72.720 ;
        RECT 358.410 72.520 1326.110 72.660 ;
        RECT 358.410 72.460 358.730 72.520 ;
        RECT 1325.790 72.460 1326.110 72.520 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 358.410 16.900 358.730 16.960 ;
        RECT 353.350 16.760 358.730 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 358.410 16.700 358.730 16.760 ;
      LAYER via ;
        RECT 1326.280 1642.240 1326.540 1642.500 ;
        RECT 1327.660 1642.240 1327.920 1642.500 ;
        RECT 1325.820 1497.400 1326.080 1497.660 ;
        RECT 1326.280 1497.400 1326.540 1497.660 ;
        RECT 1326.280 1490.260 1326.540 1490.520 ;
        RECT 1326.280 1441.980 1326.540 1442.240 ;
        RECT 1325.820 1400.500 1326.080 1400.760 ;
        RECT 1326.280 1400.500 1326.540 1400.760 ;
        RECT 1325.820 1152.640 1326.080 1152.900 ;
        RECT 1326.280 1152.640 1326.540 1152.900 ;
        RECT 1325.820 1124.080 1326.080 1124.340 ;
        RECT 1326.740 1124.080 1327.000 1124.340 ;
        RECT 1325.820 1048.600 1326.080 1048.860 ;
        RECT 1326.280 1013.920 1326.540 1014.180 ;
        RECT 1325.820 966.320 1326.080 966.580 ;
        RECT 1326.740 966.320 1327.000 966.580 ;
        RECT 1326.280 870.100 1326.540 870.360 ;
        RECT 1326.280 869.420 1326.540 869.680 ;
        RECT 1326.280 806.860 1326.540 807.120 ;
        RECT 1326.280 758.920 1326.540 759.180 ;
        RECT 1326.740 662.020 1327.000 662.280 ;
        RECT 1326.740 622.920 1327.000 623.180 ;
        RECT 1325.820 579.400 1326.080 579.660 ;
        RECT 1326.280 579.400 1326.540 579.660 ;
        RECT 1325.820 475.700 1326.080 475.960 ;
        RECT 1325.820 427.760 1326.080 428.020 ;
        RECT 1325.820 241.440 1326.080 241.700 ;
        RECT 1326.740 241.440 1327.000 241.700 ;
        RECT 1325.820 144.540 1326.080 144.800 ;
        RECT 1326.280 144.540 1326.540 144.800 ;
        RECT 358.440 72.460 358.700 72.720 ;
        RECT 1325.820 72.460 1326.080 72.720 ;
        RECT 353.380 16.700 353.640 16.960 ;
        RECT 358.440 16.700 358.700 16.960 ;
      LAYER met2 ;
        RECT 1330.340 1701.090 1330.620 1702.400 ;
        RECT 1327.720 1700.950 1330.620 1701.090 ;
        RECT 1327.720 1642.530 1327.860 1700.950 ;
        RECT 1330.340 1700.000 1330.620 1700.950 ;
        RECT 1326.280 1642.210 1326.540 1642.530 ;
        RECT 1327.660 1642.210 1327.920 1642.530 ;
        RECT 1326.340 1559.650 1326.480 1642.210 ;
        RECT 1325.880 1559.510 1326.480 1559.650 ;
        RECT 1325.880 1497.690 1326.020 1559.510 ;
        RECT 1325.820 1497.370 1326.080 1497.690 ;
        RECT 1326.280 1497.370 1326.540 1497.690 ;
        RECT 1326.340 1490.550 1326.480 1497.370 ;
        RECT 1326.280 1490.230 1326.540 1490.550 ;
        RECT 1326.280 1441.950 1326.540 1442.270 ;
        RECT 1326.340 1424.330 1326.480 1441.950 ;
        RECT 1326.340 1424.190 1326.940 1424.330 ;
        RECT 1326.800 1414.130 1326.940 1424.190 ;
        RECT 1326.340 1413.990 1326.940 1414.130 ;
        RECT 1326.340 1400.790 1326.480 1413.990 ;
        RECT 1325.820 1400.470 1326.080 1400.790 ;
        RECT 1326.280 1400.470 1326.540 1400.790 ;
        RECT 1325.880 1345.565 1326.020 1400.470 ;
        RECT 1325.810 1345.195 1326.090 1345.565 ;
        RECT 1327.190 1345.195 1327.470 1345.565 ;
        RECT 1327.260 1269.970 1327.400 1345.195 ;
        RECT 1326.340 1269.830 1327.400 1269.970 ;
        RECT 1326.340 1152.930 1326.480 1269.830 ;
        RECT 1325.820 1152.610 1326.080 1152.930 ;
        RECT 1326.280 1152.610 1326.540 1152.930 ;
        RECT 1325.880 1152.445 1326.020 1152.610 ;
        RECT 1325.810 1152.075 1326.090 1152.445 ;
        RECT 1326.730 1152.075 1327.010 1152.445 ;
        RECT 1326.800 1124.370 1326.940 1152.075 ;
        RECT 1325.820 1124.050 1326.080 1124.370 ;
        RECT 1326.740 1124.050 1327.000 1124.370 ;
        RECT 1325.880 1048.890 1326.020 1124.050 ;
        RECT 1325.820 1048.570 1326.080 1048.890 ;
        RECT 1326.280 1013.890 1326.540 1014.210 ;
        RECT 1326.340 1000.690 1326.480 1013.890 ;
        RECT 1326.340 1000.550 1326.940 1000.690 ;
        RECT 1326.800 966.610 1326.940 1000.550 ;
        RECT 1325.820 966.290 1326.080 966.610 ;
        RECT 1326.740 966.290 1327.000 966.610 ;
        RECT 1325.880 966.010 1326.020 966.290 ;
        RECT 1325.880 965.870 1326.480 966.010 ;
        RECT 1326.340 870.390 1326.480 965.870 ;
        RECT 1326.280 870.070 1326.540 870.390 ;
        RECT 1326.280 869.620 1326.540 869.710 ;
        RECT 1325.880 869.480 1326.540 869.620 ;
        RECT 1325.880 821.965 1326.020 869.480 ;
        RECT 1326.280 869.390 1326.540 869.480 ;
        RECT 1325.810 821.595 1326.090 821.965 ;
        RECT 1326.270 820.915 1326.550 821.285 ;
        RECT 1326.340 807.150 1326.480 820.915 ;
        RECT 1326.280 806.830 1326.540 807.150 ;
        RECT 1326.280 758.890 1326.540 759.210 ;
        RECT 1326.340 717.925 1326.480 758.890 ;
        RECT 1326.270 717.555 1326.550 717.925 ;
        RECT 1327.190 716.875 1327.470 717.245 ;
        RECT 1327.260 662.730 1327.400 716.875 ;
        RECT 1326.800 662.590 1327.400 662.730 ;
        RECT 1326.800 662.310 1326.940 662.590 ;
        RECT 1326.740 661.990 1327.000 662.310 ;
        RECT 1326.740 622.890 1327.000 623.210 ;
        RECT 1326.800 579.885 1326.940 622.890 ;
        RECT 1325.810 579.515 1326.090 579.885 ;
        RECT 1325.820 579.370 1326.080 579.515 ;
        RECT 1326.280 579.370 1326.540 579.690 ;
        RECT 1326.730 579.515 1327.010 579.885 ;
        RECT 1326.340 476.410 1326.480 579.370 ;
        RECT 1325.880 476.270 1326.480 476.410 ;
        RECT 1325.880 475.990 1326.020 476.270 ;
        RECT 1325.820 475.670 1326.080 475.990 ;
        RECT 1325.820 427.730 1326.080 428.050 ;
        RECT 1325.880 385.970 1326.020 427.730 ;
        RECT 1325.880 385.830 1326.480 385.970 ;
        RECT 1326.340 364.890 1326.480 385.830 ;
        RECT 1326.340 364.750 1326.940 364.890 ;
        RECT 1326.800 241.730 1326.940 364.750 ;
        RECT 1325.820 241.410 1326.080 241.730 ;
        RECT 1326.740 241.410 1327.000 241.730 ;
        RECT 1325.880 192.170 1326.020 241.410 ;
        RECT 1325.880 192.030 1326.480 192.170 ;
        RECT 1326.340 144.830 1326.480 192.030 ;
        RECT 1325.820 144.510 1326.080 144.830 ;
        RECT 1326.280 144.510 1326.540 144.830 ;
        RECT 1325.880 72.750 1326.020 144.510 ;
        RECT 358.440 72.430 358.700 72.750 ;
        RECT 1325.820 72.430 1326.080 72.750 ;
        RECT 358.500 16.990 358.640 72.430 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 358.440 16.670 358.700 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
      LAYER via2 ;
        RECT 1325.810 1345.240 1326.090 1345.520 ;
        RECT 1327.190 1345.240 1327.470 1345.520 ;
        RECT 1325.810 1152.120 1326.090 1152.400 ;
        RECT 1326.730 1152.120 1327.010 1152.400 ;
        RECT 1325.810 821.640 1326.090 821.920 ;
        RECT 1326.270 820.960 1326.550 821.240 ;
        RECT 1326.270 717.600 1326.550 717.880 ;
        RECT 1327.190 716.920 1327.470 717.200 ;
        RECT 1325.810 579.560 1326.090 579.840 ;
        RECT 1326.730 579.560 1327.010 579.840 ;
      LAYER met3 ;
        RECT 1325.785 1345.530 1326.115 1345.545 ;
        RECT 1327.165 1345.530 1327.495 1345.545 ;
        RECT 1325.785 1345.230 1327.495 1345.530 ;
        RECT 1325.785 1345.215 1326.115 1345.230 ;
        RECT 1327.165 1345.215 1327.495 1345.230 ;
        RECT 1325.785 1152.410 1326.115 1152.425 ;
        RECT 1326.705 1152.410 1327.035 1152.425 ;
        RECT 1325.785 1152.110 1327.035 1152.410 ;
        RECT 1325.785 1152.095 1326.115 1152.110 ;
        RECT 1326.705 1152.095 1327.035 1152.110 ;
        RECT 1325.785 821.930 1326.115 821.945 ;
        RECT 1325.785 821.615 1326.330 821.930 ;
        RECT 1326.030 821.265 1326.330 821.615 ;
        RECT 1326.030 820.950 1326.575 821.265 ;
        RECT 1326.245 820.935 1326.575 820.950 ;
        RECT 1326.245 717.890 1326.575 717.905 ;
        RECT 1326.030 717.575 1326.575 717.890 ;
        RECT 1326.030 717.210 1326.330 717.575 ;
        RECT 1327.165 717.210 1327.495 717.225 ;
        RECT 1326.030 716.910 1327.495 717.210 ;
        RECT 1327.165 716.895 1327.495 716.910 ;
        RECT 1325.785 579.850 1326.115 579.865 ;
        RECT 1326.705 579.850 1327.035 579.865 ;
        RECT 1325.785 579.550 1327.035 579.850 ;
        RECT 1325.785 579.535 1326.115 579.550 ;
        RECT 1326.705 579.535 1327.035 579.550 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 73.000 372.530 73.060 ;
        RECT 1339.130 73.000 1339.450 73.060 ;
        RECT 372.210 72.860 1339.450 73.000 ;
        RECT 372.210 72.800 372.530 72.860 ;
        RECT 1339.130 72.800 1339.450 72.860 ;
      LAYER via ;
        RECT 372.240 72.800 372.500 73.060 ;
        RECT 1339.160 72.800 1339.420 73.060 ;
      LAYER met2 ;
        RECT 1339.540 1700.410 1339.820 1702.400 ;
        RECT 1339.220 1700.270 1339.820 1700.410 ;
        RECT 1339.220 73.090 1339.360 1700.270 ;
        RECT 1339.540 1700.000 1339.820 1700.270 ;
        RECT 372.240 72.770 372.500 73.090 ;
        RECT 1339.160 72.770 1339.420 73.090 ;
        RECT 372.300 16.900 372.440 72.770 ;
        RECT 371.380 16.760 372.440 16.900 ;
        RECT 371.380 2.400 371.520 16.760 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 73.340 393.230 73.400 ;
        RECT 1346.030 73.340 1346.350 73.400 ;
        RECT 392.910 73.200 1346.350 73.340 ;
        RECT 392.910 73.140 393.230 73.200 ;
        RECT 1346.030 73.140 1346.350 73.200 ;
        RECT 389.230 16.220 389.550 16.280 ;
        RECT 392.910 16.220 393.230 16.280 ;
        RECT 389.230 16.080 393.230 16.220 ;
        RECT 389.230 16.020 389.550 16.080 ;
        RECT 392.910 16.020 393.230 16.080 ;
      LAYER via ;
        RECT 392.940 73.140 393.200 73.400 ;
        RECT 1346.060 73.140 1346.320 73.400 ;
        RECT 389.260 16.020 389.520 16.280 ;
        RECT 392.940 16.020 393.200 16.280 ;
      LAYER met2 ;
        RECT 1348.740 1700.410 1349.020 1702.400 ;
        RECT 1346.120 1700.270 1349.020 1700.410 ;
        RECT 1346.120 73.430 1346.260 1700.270 ;
        RECT 1348.740 1700.000 1349.020 1700.270 ;
        RECT 392.940 73.110 393.200 73.430 ;
        RECT 1346.060 73.110 1346.320 73.430 ;
        RECT 393.000 16.310 393.140 73.110 ;
        RECT 389.260 15.990 389.520 16.310 ;
        RECT 392.940 15.990 393.200 16.310 ;
        RECT 389.320 2.400 389.460 15.990 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1353.465 1497.445 1353.635 1545.555 ;
        RECT 1353.005 1345.465 1353.175 1393.575 ;
        RECT 1353.925 965.685 1354.095 980.475 ;
        RECT 1353.465 737.885 1353.635 772.735 ;
        RECT 1353.465 641.325 1353.635 676.175 ;
        RECT 1354.385 462.485 1354.555 510.595 ;
        RECT 1353.465 324.445 1353.635 414.035 ;
        RECT 1353.005 234.685 1353.175 287.895 ;
        RECT 1353.465 73.525 1353.635 113.135 ;
      LAYER mcon ;
        RECT 1353.465 1545.385 1353.635 1545.555 ;
        RECT 1353.005 1393.405 1353.175 1393.575 ;
        RECT 1353.925 980.305 1354.095 980.475 ;
        RECT 1353.465 772.565 1353.635 772.735 ;
        RECT 1353.465 676.005 1353.635 676.175 ;
        RECT 1354.385 510.425 1354.555 510.595 ;
        RECT 1353.465 413.865 1353.635 414.035 ;
        RECT 1353.005 287.725 1353.175 287.895 ;
        RECT 1353.465 112.965 1353.635 113.135 ;
      LAYER met1 ;
        RECT 1353.850 1642.440 1354.170 1642.500 ;
        RECT 1355.230 1642.440 1355.550 1642.500 ;
        RECT 1353.850 1642.300 1355.550 1642.440 ;
        RECT 1353.850 1642.240 1354.170 1642.300 ;
        RECT 1355.230 1642.240 1355.550 1642.300 ;
        RECT 1353.390 1545.540 1353.710 1545.600 ;
        RECT 1353.195 1545.400 1353.710 1545.540 ;
        RECT 1353.390 1545.340 1353.710 1545.400 ;
        RECT 1353.405 1497.600 1353.695 1497.645 ;
        RECT 1353.850 1497.600 1354.170 1497.660 ;
        RECT 1353.405 1497.460 1354.170 1497.600 ;
        RECT 1353.405 1497.415 1353.695 1497.460 ;
        RECT 1353.850 1497.400 1354.170 1497.460 ;
        RECT 1353.850 1490.460 1354.170 1490.520 ;
        RECT 1354.310 1490.460 1354.630 1490.520 ;
        RECT 1353.850 1490.320 1354.630 1490.460 ;
        RECT 1353.850 1490.260 1354.170 1490.320 ;
        RECT 1354.310 1490.260 1354.630 1490.320 ;
        RECT 1352.930 1400.700 1353.250 1400.760 ;
        RECT 1354.310 1400.700 1354.630 1400.760 ;
        RECT 1352.930 1400.560 1354.630 1400.700 ;
        RECT 1352.930 1400.500 1353.250 1400.560 ;
        RECT 1354.310 1400.500 1354.630 1400.560 ;
        RECT 1352.930 1393.560 1353.250 1393.620 ;
        RECT 1352.735 1393.420 1353.250 1393.560 ;
        RECT 1352.930 1393.360 1353.250 1393.420 ;
        RECT 1352.945 1345.620 1353.235 1345.665 ;
        RECT 1353.850 1345.620 1354.170 1345.680 ;
        RECT 1352.945 1345.480 1354.170 1345.620 ;
        RECT 1352.945 1345.435 1353.235 1345.480 ;
        RECT 1353.850 1345.420 1354.170 1345.480 ;
        RECT 1352.930 1255.860 1353.250 1255.920 ;
        RECT 1354.770 1255.860 1355.090 1255.920 ;
        RECT 1352.930 1255.720 1355.090 1255.860 ;
        RECT 1352.930 1255.660 1353.250 1255.720 ;
        RECT 1354.770 1255.660 1355.090 1255.720 ;
        RECT 1353.850 1062.740 1354.170 1062.800 ;
        RECT 1354.770 1062.740 1355.090 1062.800 ;
        RECT 1353.850 1062.600 1355.090 1062.740 ;
        RECT 1353.850 1062.540 1354.170 1062.600 ;
        RECT 1354.770 1062.540 1355.090 1062.600 ;
        RECT 1353.850 980.460 1354.170 980.520 ;
        RECT 1353.655 980.320 1354.170 980.460 ;
        RECT 1353.850 980.260 1354.170 980.320 ;
        RECT 1353.850 965.840 1354.170 965.900 ;
        RECT 1353.655 965.700 1354.170 965.840 ;
        RECT 1353.850 965.640 1354.170 965.700 ;
        RECT 1352.010 959.040 1352.330 959.100 ;
        RECT 1353.850 959.040 1354.170 959.100 ;
        RECT 1352.010 958.900 1354.170 959.040 ;
        RECT 1352.010 958.840 1352.330 958.900 ;
        RECT 1353.850 958.840 1354.170 958.900 ;
        RECT 1352.930 910.760 1353.250 910.820 ;
        RECT 1354.310 910.760 1354.630 910.820 ;
        RECT 1352.930 910.620 1354.630 910.760 ;
        RECT 1352.930 910.560 1353.250 910.620 ;
        RECT 1354.310 910.560 1354.630 910.620 ;
        RECT 1353.390 835.080 1353.710 835.340 ;
        RECT 1353.480 834.600 1353.620 835.080 ;
        RECT 1353.850 834.600 1354.170 834.660 ;
        RECT 1353.480 834.460 1354.170 834.600 ;
        RECT 1353.850 834.400 1354.170 834.460 ;
        RECT 1353.390 772.720 1353.710 772.780 ;
        RECT 1353.195 772.580 1353.710 772.720 ;
        RECT 1353.390 772.520 1353.710 772.580 ;
        RECT 1353.390 738.040 1353.710 738.100 ;
        RECT 1353.195 737.900 1353.710 738.040 ;
        RECT 1353.390 737.840 1353.710 737.900 ;
        RECT 1353.390 676.160 1353.710 676.220 ;
        RECT 1353.195 676.020 1353.710 676.160 ;
        RECT 1353.390 675.960 1353.710 676.020 ;
        RECT 1353.390 641.480 1353.710 641.540 ;
        RECT 1353.195 641.340 1353.710 641.480 ;
        RECT 1353.390 641.280 1353.710 641.340 ;
        RECT 1353.850 603.540 1354.170 603.800 ;
        RECT 1353.940 603.120 1354.080 603.540 ;
        RECT 1353.850 602.860 1354.170 603.120 ;
        RECT 1354.310 510.580 1354.630 510.640 ;
        RECT 1354.115 510.440 1354.630 510.580 ;
        RECT 1354.310 510.380 1354.630 510.440 ;
        RECT 1354.325 462.640 1354.615 462.685 ;
        RECT 1354.770 462.640 1355.090 462.700 ;
        RECT 1354.325 462.500 1355.090 462.640 ;
        RECT 1354.325 462.455 1354.615 462.500 ;
        RECT 1354.770 462.440 1355.090 462.500 ;
        RECT 1353.405 414.020 1353.695 414.065 ;
        RECT 1354.770 414.020 1355.090 414.080 ;
        RECT 1353.405 413.880 1355.090 414.020 ;
        RECT 1353.405 413.835 1353.695 413.880 ;
        RECT 1354.770 413.820 1355.090 413.880 ;
        RECT 1353.390 324.600 1353.710 324.660 ;
        RECT 1353.195 324.460 1353.710 324.600 ;
        RECT 1353.390 324.400 1353.710 324.460 ;
        RECT 1352.945 287.880 1353.235 287.925 ;
        RECT 1353.390 287.880 1353.710 287.940 ;
        RECT 1352.945 287.740 1353.710 287.880 ;
        RECT 1352.945 287.695 1353.235 287.740 ;
        RECT 1353.390 287.680 1353.710 287.740 ;
        RECT 1352.930 234.840 1353.250 234.900 ;
        RECT 1352.735 234.700 1353.250 234.840 ;
        RECT 1352.930 234.640 1353.250 234.700 ;
        RECT 1353.390 145.220 1353.710 145.480 ;
        RECT 1353.480 145.080 1353.620 145.220 ;
        RECT 1353.850 145.080 1354.170 145.140 ;
        RECT 1353.480 144.940 1354.170 145.080 ;
        RECT 1353.850 144.880 1354.170 144.940 ;
        RECT 1353.405 113.120 1353.695 113.165 ;
        RECT 1353.850 113.120 1354.170 113.180 ;
        RECT 1353.405 112.980 1354.170 113.120 ;
        RECT 1353.405 112.935 1353.695 112.980 ;
        RECT 1353.850 112.920 1354.170 112.980 ;
        RECT 413.610 73.680 413.930 73.740 ;
        RECT 1353.405 73.680 1353.695 73.725 ;
        RECT 413.610 73.540 1353.695 73.680 ;
        RECT 413.610 73.480 413.930 73.540 ;
        RECT 1353.405 73.495 1353.695 73.540 ;
        RECT 407.170 16.220 407.490 16.280 ;
        RECT 413.610 16.220 413.930 16.280 ;
        RECT 407.170 16.080 413.930 16.220 ;
        RECT 407.170 16.020 407.490 16.080 ;
        RECT 413.610 16.020 413.930 16.080 ;
      LAYER via ;
        RECT 1353.880 1642.240 1354.140 1642.500 ;
        RECT 1355.260 1642.240 1355.520 1642.500 ;
        RECT 1353.420 1545.340 1353.680 1545.600 ;
        RECT 1353.880 1497.400 1354.140 1497.660 ;
        RECT 1353.880 1490.260 1354.140 1490.520 ;
        RECT 1354.340 1490.260 1354.600 1490.520 ;
        RECT 1352.960 1400.500 1353.220 1400.760 ;
        RECT 1354.340 1400.500 1354.600 1400.760 ;
        RECT 1352.960 1393.360 1353.220 1393.620 ;
        RECT 1353.880 1345.420 1354.140 1345.680 ;
        RECT 1352.960 1255.660 1353.220 1255.920 ;
        RECT 1354.800 1255.660 1355.060 1255.920 ;
        RECT 1353.880 1062.540 1354.140 1062.800 ;
        RECT 1354.800 1062.540 1355.060 1062.800 ;
        RECT 1353.880 980.260 1354.140 980.520 ;
        RECT 1353.880 965.640 1354.140 965.900 ;
        RECT 1352.040 958.840 1352.300 959.100 ;
        RECT 1353.880 958.840 1354.140 959.100 ;
        RECT 1352.960 910.560 1353.220 910.820 ;
        RECT 1354.340 910.560 1354.600 910.820 ;
        RECT 1353.420 835.080 1353.680 835.340 ;
        RECT 1353.880 834.400 1354.140 834.660 ;
        RECT 1353.420 772.520 1353.680 772.780 ;
        RECT 1353.420 737.840 1353.680 738.100 ;
        RECT 1353.420 675.960 1353.680 676.220 ;
        RECT 1353.420 641.280 1353.680 641.540 ;
        RECT 1353.880 603.540 1354.140 603.800 ;
        RECT 1353.880 602.860 1354.140 603.120 ;
        RECT 1354.340 510.380 1354.600 510.640 ;
        RECT 1354.800 462.440 1355.060 462.700 ;
        RECT 1354.800 413.820 1355.060 414.080 ;
        RECT 1353.420 324.400 1353.680 324.660 ;
        RECT 1353.420 287.680 1353.680 287.940 ;
        RECT 1352.960 234.640 1353.220 234.900 ;
        RECT 1353.420 145.220 1353.680 145.480 ;
        RECT 1353.880 144.880 1354.140 145.140 ;
        RECT 1353.880 112.920 1354.140 113.180 ;
        RECT 413.640 73.480 413.900 73.740 ;
        RECT 407.200 16.020 407.460 16.280 ;
        RECT 413.640 16.020 413.900 16.280 ;
      LAYER met2 ;
        RECT 1357.940 1701.090 1358.220 1702.400 ;
        RECT 1355.320 1700.950 1358.220 1701.090 ;
        RECT 1355.320 1642.530 1355.460 1700.950 ;
        RECT 1357.940 1700.000 1358.220 1700.950 ;
        RECT 1353.880 1642.210 1354.140 1642.530 ;
        RECT 1355.260 1642.210 1355.520 1642.530 ;
        RECT 1353.940 1559.650 1354.080 1642.210 ;
        RECT 1353.480 1559.510 1354.080 1559.650 ;
        RECT 1353.480 1545.630 1353.620 1559.510 ;
        RECT 1353.420 1545.310 1353.680 1545.630 ;
        RECT 1353.880 1497.370 1354.140 1497.690 ;
        RECT 1353.940 1490.550 1354.080 1497.370 ;
        RECT 1353.880 1490.230 1354.140 1490.550 ;
        RECT 1354.340 1490.230 1354.600 1490.550 ;
        RECT 1354.400 1400.790 1354.540 1490.230 ;
        RECT 1352.960 1400.470 1353.220 1400.790 ;
        RECT 1354.340 1400.470 1354.600 1400.790 ;
        RECT 1353.020 1393.650 1353.160 1400.470 ;
        RECT 1352.960 1393.330 1353.220 1393.650 ;
        RECT 1353.880 1345.390 1354.140 1345.710 ;
        RECT 1353.940 1304.085 1354.080 1345.390 ;
        RECT 1353.870 1303.715 1354.150 1304.085 ;
        RECT 1352.950 1303.035 1353.230 1303.405 ;
        RECT 1353.020 1255.950 1353.160 1303.035 ;
        RECT 1352.960 1255.630 1353.220 1255.950 ;
        RECT 1354.800 1255.630 1355.060 1255.950 ;
        RECT 1354.860 1159.810 1355.000 1255.630 ;
        RECT 1353.940 1159.670 1355.000 1159.810 ;
        RECT 1353.940 1159.130 1354.080 1159.670 ;
        RECT 1353.940 1158.990 1355.000 1159.130 ;
        RECT 1354.860 1062.830 1355.000 1158.990 ;
        RECT 1353.880 1062.510 1354.140 1062.830 ;
        RECT 1354.800 1062.510 1355.060 1062.830 ;
        RECT 1353.940 1028.570 1354.080 1062.510 ;
        RECT 1353.020 1028.430 1354.080 1028.570 ;
        RECT 1353.020 1015.765 1353.160 1028.430 ;
        RECT 1352.950 1015.395 1353.230 1015.765 ;
        RECT 1353.870 1014.715 1354.150 1015.085 ;
        RECT 1353.940 980.550 1354.080 1014.715 ;
        RECT 1353.880 980.230 1354.140 980.550 ;
        RECT 1353.880 965.610 1354.140 965.930 ;
        RECT 1353.940 959.130 1354.080 965.610 ;
        RECT 1352.040 958.810 1352.300 959.130 ;
        RECT 1353.880 958.810 1354.140 959.130 ;
        RECT 1352.100 911.045 1352.240 958.810 ;
        RECT 1352.030 910.675 1352.310 911.045 ;
        RECT 1352.950 910.675 1353.230 911.045 ;
        RECT 1352.960 910.530 1353.220 910.675 ;
        RECT 1354.340 910.530 1354.600 910.850 ;
        RECT 1354.400 862.765 1354.540 910.530 ;
        RECT 1353.410 862.395 1353.690 862.765 ;
        RECT 1354.330 862.395 1354.610 862.765 ;
        RECT 1353.480 835.370 1353.620 862.395 ;
        RECT 1353.420 835.050 1353.680 835.370 ;
        RECT 1353.880 834.370 1354.140 834.690 ;
        RECT 1353.940 787.850 1354.080 834.370 ;
        RECT 1353.940 787.710 1354.540 787.850 ;
        RECT 1354.400 773.685 1354.540 787.710 ;
        RECT 1354.330 773.315 1354.610 773.685 ;
        RECT 1353.410 772.635 1353.690 773.005 ;
        RECT 1353.420 772.490 1353.680 772.635 ;
        RECT 1353.420 737.810 1353.680 738.130 ;
        RECT 1353.480 724.610 1353.620 737.810 ;
        RECT 1353.480 724.470 1354.080 724.610 ;
        RECT 1353.940 691.290 1354.080 724.470 ;
        RECT 1353.940 691.150 1354.540 691.290 ;
        RECT 1354.400 676.445 1354.540 691.150 ;
        RECT 1353.410 676.075 1353.690 676.445 ;
        RECT 1354.330 676.075 1354.610 676.445 ;
        RECT 1353.420 675.930 1353.680 676.075 ;
        RECT 1353.420 641.250 1353.680 641.570 ;
        RECT 1353.480 628.050 1353.620 641.250 ;
        RECT 1353.480 627.910 1354.080 628.050 ;
        RECT 1353.940 603.830 1354.080 627.910 ;
        RECT 1353.880 603.510 1354.140 603.830 ;
        RECT 1353.880 602.830 1354.140 603.150 ;
        RECT 1353.940 555.290 1354.080 602.830 ;
        RECT 1353.940 555.150 1354.540 555.290 ;
        RECT 1354.400 510.670 1354.540 555.150 ;
        RECT 1354.340 510.350 1354.600 510.670 ;
        RECT 1354.800 462.410 1355.060 462.730 ;
        RECT 1354.860 414.110 1355.000 462.410 ;
        RECT 1354.800 413.790 1355.060 414.110 ;
        RECT 1353.420 324.370 1353.680 324.690 ;
        RECT 1353.480 287.970 1353.620 324.370 ;
        RECT 1353.420 287.650 1353.680 287.970 ;
        RECT 1352.960 234.610 1353.220 234.930 ;
        RECT 1353.020 193.530 1353.160 234.610 ;
        RECT 1353.020 193.390 1353.620 193.530 ;
        RECT 1353.480 145.510 1353.620 193.390 ;
        RECT 1353.420 145.190 1353.680 145.510 ;
        RECT 1353.880 144.850 1354.140 145.170 ;
        RECT 1353.940 113.210 1354.080 144.850 ;
        RECT 1353.880 112.890 1354.140 113.210 ;
        RECT 413.640 73.450 413.900 73.770 ;
        RECT 413.700 16.310 413.840 73.450 ;
        RECT 407.200 15.990 407.460 16.310 ;
        RECT 413.640 15.990 413.900 16.310 ;
        RECT 407.260 2.400 407.400 15.990 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 1353.870 1303.760 1354.150 1304.040 ;
        RECT 1352.950 1303.080 1353.230 1303.360 ;
        RECT 1352.950 1015.440 1353.230 1015.720 ;
        RECT 1353.870 1014.760 1354.150 1015.040 ;
        RECT 1352.030 910.720 1352.310 911.000 ;
        RECT 1352.950 910.720 1353.230 911.000 ;
        RECT 1353.410 862.440 1353.690 862.720 ;
        RECT 1354.330 862.440 1354.610 862.720 ;
        RECT 1354.330 773.360 1354.610 773.640 ;
        RECT 1353.410 772.680 1353.690 772.960 ;
        RECT 1353.410 676.120 1353.690 676.400 ;
        RECT 1354.330 676.120 1354.610 676.400 ;
      LAYER met3 ;
        RECT 1353.845 1304.050 1354.175 1304.065 ;
        RECT 1353.845 1303.750 1354.850 1304.050 ;
        RECT 1353.845 1303.735 1354.175 1303.750 ;
        RECT 1352.925 1303.370 1353.255 1303.385 ;
        RECT 1354.550 1303.370 1354.850 1303.750 ;
        RECT 1352.925 1303.070 1354.850 1303.370 ;
        RECT 1352.925 1303.055 1353.255 1303.070 ;
        RECT 1352.925 1015.730 1353.255 1015.745 ;
        RECT 1352.925 1015.430 1354.850 1015.730 ;
        RECT 1352.925 1015.415 1353.255 1015.430 ;
        RECT 1353.845 1015.050 1354.175 1015.065 ;
        RECT 1354.550 1015.050 1354.850 1015.430 ;
        RECT 1353.845 1014.750 1354.850 1015.050 ;
        RECT 1353.845 1014.735 1354.175 1014.750 ;
        RECT 1352.005 911.010 1352.335 911.025 ;
        RECT 1352.925 911.010 1353.255 911.025 ;
        RECT 1352.005 910.710 1353.255 911.010 ;
        RECT 1352.005 910.695 1352.335 910.710 ;
        RECT 1352.925 910.695 1353.255 910.710 ;
        RECT 1353.385 862.730 1353.715 862.745 ;
        RECT 1354.305 862.730 1354.635 862.745 ;
        RECT 1353.385 862.430 1354.635 862.730 ;
        RECT 1353.385 862.415 1353.715 862.430 ;
        RECT 1354.305 862.415 1354.635 862.430 ;
        RECT 1354.305 773.650 1354.635 773.665 ;
        RECT 1352.710 773.350 1354.635 773.650 ;
        RECT 1352.710 772.970 1353.010 773.350 ;
        RECT 1354.305 773.335 1354.635 773.350 ;
        RECT 1353.385 772.970 1353.715 772.985 ;
        RECT 1352.710 772.670 1353.715 772.970 ;
        RECT 1353.385 772.655 1353.715 772.670 ;
        RECT 1353.385 676.410 1353.715 676.425 ;
        RECT 1354.305 676.410 1354.635 676.425 ;
        RECT 1353.385 676.110 1354.635 676.410 ;
        RECT 1353.385 676.095 1353.715 676.110 ;
        RECT 1354.305 676.095 1354.635 676.110 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1163.945 58.565 1164.115 62.475 ;
      LAYER mcon ;
        RECT 1163.945 62.305 1164.115 62.475 ;
      LAYER met1 ;
        RECT 1163.885 62.460 1164.175 62.505 ;
        RECT 1180.890 62.460 1181.210 62.520 ;
        RECT 1163.885 62.320 1181.210 62.460 ;
        RECT 1163.885 62.275 1164.175 62.320 ;
        RECT 1180.890 62.260 1181.210 62.320 ;
        RECT 68.150 58.720 68.470 58.780 ;
        RECT 1163.885 58.720 1164.175 58.765 ;
        RECT 68.150 58.580 1164.175 58.720 ;
        RECT 68.150 58.520 68.470 58.580 ;
        RECT 1163.885 58.535 1164.175 58.580 ;
      LAYER via ;
        RECT 1180.920 62.260 1181.180 62.520 ;
        RECT 68.180 58.520 68.440 58.780 ;
      LAYER met2 ;
        RECT 1183.600 1700.410 1183.880 1702.400 ;
        RECT 1180.980 1700.270 1183.880 1700.410 ;
        RECT 1180.980 62.550 1181.120 1700.270 ;
        RECT 1183.600 1700.000 1183.880 1700.270 ;
        RECT 1180.920 62.230 1181.180 62.550 ;
        RECT 68.180 58.490 68.440 58.810 ;
        RECT 68.240 2.400 68.380 58.490 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 74.020 427.730 74.080 ;
        RECT 1366.730 74.020 1367.050 74.080 ;
        RECT 427.410 73.880 1367.050 74.020 ;
        RECT 427.410 73.820 427.730 73.880 ;
        RECT 1366.730 73.820 1367.050 73.880 ;
        RECT 424.650 16.220 424.970 16.280 ;
        RECT 427.410 16.220 427.730 16.280 ;
        RECT 424.650 16.080 427.730 16.220 ;
        RECT 424.650 16.020 424.970 16.080 ;
        RECT 427.410 16.020 427.730 16.080 ;
      LAYER via ;
        RECT 427.440 73.820 427.700 74.080 ;
        RECT 1366.760 73.820 1367.020 74.080 ;
        RECT 424.680 16.020 424.940 16.280 ;
        RECT 427.440 16.020 427.700 16.280 ;
      LAYER met2 ;
        RECT 1367.140 1700.410 1367.420 1702.400 ;
        RECT 1366.820 1700.270 1367.420 1700.410 ;
        RECT 1366.820 74.110 1366.960 1700.270 ;
        RECT 1367.140 1700.000 1367.420 1700.270 ;
        RECT 427.440 73.790 427.700 74.110 ;
        RECT 1366.760 73.790 1367.020 74.110 ;
        RECT 427.500 16.310 427.640 73.790 ;
        RECT 424.680 15.990 424.940 16.310 ;
        RECT 427.440 15.990 427.700 16.310 ;
        RECT 424.740 2.400 424.880 15.990 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 74.360 448.430 74.420 ;
        RECT 1373.630 74.360 1373.950 74.420 ;
        RECT 448.110 74.220 1373.950 74.360 ;
        RECT 448.110 74.160 448.430 74.220 ;
        RECT 1373.630 74.160 1373.950 74.220 ;
        RECT 442.590 16.220 442.910 16.280 ;
        RECT 448.110 16.220 448.430 16.280 ;
        RECT 442.590 16.080 448.430 16.220 ;
        RECT 442.590 16.020 442.910 16.080 ;
        RECT 448.110 16.020 448.430 16.080 ;
      LAYER via ;
        RECT 448.140 74.160 448.400 74.420 ;
        RECT 1373.660 74.160 1373.920 74.420 ;
        RECT 442.620 16.020 442.880 16.280 ;
        RECT 448.140 16.020 448.400 16.280 ;
      LAYER met2 ;
        RECT 1376.340 1700.410 1376.620 1702.400 ;
        RECT 1373.720 1700.270 1376.620 1700.410 ;
        RECT 1373.720 74.450 1373.860 1700.270 ;
        RECT 1376.340 1700.000 1376.620 1700.270 ;
        RECT 448.140 74.130 448.400 74.450 ;
        RECT 1373.660 74.130 1373.920 74.450 ;
        RECT 448.200 16.310 448.340 74.130 ;
        RECT 442.620 15.990 442.880 16.310 ;
        RECT 448.140 15.990 448.400 16.310 ;
        RECT 442.680 2.400 442.820 15.990 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 74.700 462.230 74.760 ;
        RECT 1380.530 74.700 1380.850 74.760 ;
        RECT 461.910 74.560 1380.850 74.700 ;
        RECT 461.910 74.500 462.230 74.560 ;
        RECT 1380.530 74.500 1380.850 74.560 ;
      LAYER via ;
        RECT 461.940 74.500 462.200 74.760 ;
        RECT 1380.560 74.500 1380.820 74.760 ;
      LAYER met2 ;
        RECT 1385.540 1700.410 1385.820 1702.400 ;
        RECT 1382.920 1700.270 1385.820 1700.410 ;
        RECT 1382.920 1678.650 1383.060 1700.270 ;
        RECT 1385.540 1700.000 1385.820 1700.270 ;
        RECT 1380.620 1678.510 1383.060 1678.650 ;
        RECT 1380.620 74.790 1380.760 1678.510 ;
        RECT 461.940 74.470 462.200 74.790 ;
        RECT 1380.560 74.470 1380.820 74.790 ;
        RECT 462.000 17.410 462.140 74.470 ;
        RECT 460.620 17.270 462.140 17.410 ;
        RECT 460.620 2.400 460.760 17.270 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 75.040 482.930 75.100 ;
        RECT 1394.330 75.040 1394.650 75.100 ;
        RECT 482.610 74.900 1394.650 75.040 ;
        RECT 482.610 74.840 482.930 74.900 ;
        RECT 1394.330 74.840 1394.650 74.900 ;
        RECT 478.470 15.540 478.790 15.600 ;
        RECT 482.610 15.540 482.930 15.600 ;
        RECT 478.470 15.400 482.930 15.540 ;
        RECT 478.470 15.340 478.790 15.400 ;
        RECT 482.610 15.340 482.930 15.400 ;
      LAYER via ;
        RECT 482.640 74.840 482.900 75.100 ;
        RECT 1394.360 74.840 1394.620 75.100 ;
        RECT 478.500 15.340 478.760 15.600 ;
        RECT 482.640 15.340 482.900 15.600 ;
      LAYER met2 ;
        RECT 1394.740 1700.410 1395.020 1702.400 ;
        RECT 1394.420 1700.270 1395.020 1700.410 ;
        RECT 1394.420 75.130 1394.560 1700.270 ;
        RECT 1394.740 1700.000 1395.020 1700.270 ;
        RECT 482.640 74.810 482.900 75.130 ;
        RECT 1394.360 74.810 1394.620 75.130 ;
        RECT 482.700 15.630 482.840 74.810 ;
        RECT 478.500 15.310 478.760 15.630 ;
        RECT 482.640 15.310 482.900 15.630 ;
        RECT 478.560 2.400 478.700 15.310 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 75.380 496.730 75.440 ;
        RECT 1401.230 75.380 1401.550 75.440 ;
        RECT 496.410 75.240 1401.550 75.380 ;
        RECT 496.410 75.180 496.730 75.240 ;
        RECT 1401.230 75.180 1401.550 75.240 ;
      LAYER via ;
        RECT 496.440 75.180 496.700 75.440 ;
        RECT 1401.260 75.180 1401.520 75.440 ;
      LAYER met2 ;
        RECT 1403.940 1700.410 1404.220 1702.400 ;
        RECT 1401.320 1700.270 1404.220 1700.410 ;
        RECT 1401.320 75.470 1401.460 1700.270 ;
        RECT 1403.940 1700.000 1404.220 1700.270 ;
        RECT 496.440 75.150 496.700 75.470 ;
        RECT 1401.260 75.150 1401.520 75.470 ;
        RECT 496.500 2.400 496.640 75.150 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1408.205 1449.165 1408.375 1497.275 ;
        RECT 1409.585 1207.765 1409.755 1297.015 ;
        RECT 1409.585 1172.745 1409.755 1207.255 ;
        RECT 1409.585 1104.065 1409.755 1111.035 ;
        RECT 1408.665 1013.965 1408.835 1055.615 ;
        RECT 1408.205 645.065 1408.375 676.175 ;
        RECT 1408.665 282.965 1408.835 331.075 ;
      LAYER mcon ;
        RECT 1408.205 1497.105 1408.375 1497.275 ;
        RECT 1409.585 1296.845 1409.755 1297.015 ;
        RECT 1409.585 1207.085 1409.755 1207.255 ;
        RECT 1409.585 1110.865 1409.755 1111.035 ;
        RECT 1408.665 1055.445 1408.835 1055.615 ;
        RECT 1408.205 676.005 1408.375 676.175 ;
        RECT 1408.665 330.905 1408.835 331.075 ;
      LAYER met1 ;
        RECT 1408.145 1497.260 1408.435 1497.305 ;
        RECT 1409.050 1497.260 1409.370 1497.320 ;
        RECT 1408.145 1497.120 1409.370 1497.260 ;
        RECT 1408.145 1497.075 1408.435 1497.120 ;
        RECT 1409.050 1497.060 1409.370 1497.120 ;
        RECT 1408.130 1449.320 1408.450 1449.380 ;
        RECT 1407.935 1449.180 1408.450 1449.320 ;
        RECT 1408.130 1449.120 1408.450 1449.180 ;
        RECT 1408.590 1401.040 1408.910 1401.100 ;
        RECT 1409.510 1401.040 1409.830 1401.100 ;
        RECT 1408.590 1400.900 1409.830 1401.040 ;
        RECT 1408.590 1400.840 1408.910 1400.900 ;
        RECT 1409.510 1400.840 1409.830 1400.900 ;
        RECT 1409.525 1297.000 1409.815 1297.045 ;
        RECT 1409.970 1297.000 1410.290 1297.060 ;
        RECT 1409.525 1296.860 1410.290 1297.000 ;
        RECT 1409.525 1296.815 1409.815 1296.860 ;
        RECT 1409.970 1296.800 1410.290 1296.860 ;
        RECT 1409.510 1207.920 1409.830 1207.980 ;
        RECT 1409.315 1207.780 1409.830 1207.920 ;
        RECT 1409.510 1207.720 1409.830 1207.780 ;
        RECT 1409.510 1207.240 1409.830 1207.300 ;
        RECT 1409.315 1207.100 1409.830 1207.240 ;
        RECT 1409.510 1207.040 1409.830 1207.100 ;
        RECT 1409.510 1172.900 1409.830 1172.960 ;
        RECT 1409.315 1172.760 1409.830 1172.900 ;
        RECT 1409.510 1172.700 1409.830 1172.760 ;
        RECT 1409.510 1111.020 1409.830 1111.080 ;
        RECT 1409.315 1110.880 1409.830 1111.020 ;
        RECT 1409.510 1110.820 1409.830 1110.880 ;
        RECT 1409.510 1104.220 1409.830 1104.280 ;
        RECT 1409.315 1104.080 1409.830 1104.220 ;
        RECT 1409.510 1104.020 1409.830 1104.080 ;
        RECT 1409.510 1076.820 1409.830 1077.080 ;
        RECT 1409.600 1076.400 1409.740 1076.820 ;
        RECT 1409.510 1076.140 1409.830 1076.400 ;
        RECT 1408.590 1055.600 1408.910 1055.660 ;
        RECT 1408.395 1055.460 1408.910 1055.600 ;
        RECT 1408.590 1055.400 1408.910 1055.460 ;
        RECT 1408.605 1014.120 1408.895 1014.165 ;
        RECT 1409.050 1014.120 1409.370 1014.180 ;
        RECT 1408.605 1013.980 1409.370 1014.120 ;
        RECT 1408.605 1013.935 1408.895 1013.980 ;
        RECT 1409.050 1013.920 1409.370 1013.980 ;
        RECT 1409.510 980.460 1409.830 980.520 ;
        RECT 1409.140 980.320 1409.830 980.460 ;
        RECT 1409.140 979.840 1409.280 980.320 ;
        RECT 1409.510 980.260 1409.830 980.320 ;
        RECT 1409.050 979.580 1409.370 979.840 ;
        RECT 1408.590 834.940 1408.910 835.000 ;
        RECT 1409.510 834.940 1409.830 835.000 ;
        RECT 1408.590 834.800 1409.830 834.940 ;
        RECT 1408.590 834.740 1408.910 834.800 ;
        RECT 1409.510 834.740 1409.830 834.800 ;
        RECT 1409.510 787.000 1409.830 787.060 ;
        RECT 1409.140 786.860 1409.830 787.000 ;
        RECT 1409.140 786.720 1409.280 786.860 ;
        RECT 1409.510 786.800 1409.830 786.860 ;
        RECT 1409.050 786.460 1409.370 786.720 ;
        RECT 1408.130 676.160 1408.450 676.220 ;
        RECT 1407.935 676.020 1408.450 676.160 ;
        RECT 1408.130 675.960 1408.450 676.020 ;
        RECT 1408.145 645.220 1408.435 645.265 ;
        RECT 1409.050 645.220 1409.370 645.280 ;
        RECT 1408.145 645.080 1409.370 645.220 ;
        RECT 1408.145 645.035 1408.435 645.080 ;
        RECT 1409.050 645.020 1409.370 645.080 ;
        RECT 1409.050 531.320 1409.370 531.380 ;
        RECT 1409.510 531.320 1409.830 531.380 ;
        RECT 1409.050 531.180 1409.830 531.320 ;
        RECT 1409.050 531.120 1409.370 531.180 ;
        RECT 1409.510 531.120 1409.830 531.180 ;
        RECT 1409.050 483.040 1409.370 483.100 ;
        RECT 1409.970 483.040 1410.290 483.100 ;
        RECT 1409.050 482.900 1410.290 483.040 ;
        RECT 1409.050 482.840 1409.370 482.900 ;
        RECT 1409.970 482.840 1410.290 482.900 ;
        RECT 1409.050 386.820 1409.370 386.880 ;
        RECT 1409.970 386.820 1410.290 386.880 ;
        RECT 1409.050 386.680 1410.290 386.820 ;
        RECT 1409.050 386.620 1409.370 386.680 ;
        RECT 1409.970 386.620 1410.290 386.680 ;
        RECT 1409.050 362.340 1409.370 362.400 ;
        RECT 1409.970 362.340 1410.290 362.400 ;
        RECT 1409.050 362.200 1410.290 362.340 ;
        RECT 1409.050 362.140 1409.370 362.200 ;
        RECT 1409.970 362.140 1410.290 362.200 ;
        RECT 1408.590 331.060 1408.910 331.120 ;
        RECT 1408.395 330.920 1408.910 331.060 ;
        RECT 1408.590 330.860 1408.910 330.920 ;
        RECT 1408.590 283.120 1408.910 283.180 ;
        RECT 1408.395 282.980 1408.910 283.120 ;
        RECT 1408.590 282.920 1408.910 282.980 ;
        RECT 1408.590 241.640 1408.910 241.700 ;
        RECT 1409.050 241.640 1409.370 241.700 ;
        RECT 1408.590 241.500 1409.370 241.640 ;
        RECT 1408.590 241.440 1408.910 241.500 ;
        RECT 1409.050 241.440 1409.370 241.500 ;
        RECT 1408.130 193.360 1408.450 193.420 ;
        RECT 1409.050 193.360 1409.370 193.420 ;
        RECT 1408.130 193.220 1409.370 193.360 ;
        RECT 1408.130 193.160 1408.450 193.220 ;
        RECT 1409.050 193.160 1409.370 193.220 ;
        RECT 1408.130 158.680 1408.450 158.740 ;
        RECT 1409.050 158.680 1409.370 158.740 ;
        RECT 1408.130 158.540 1409.370 158.680 ;
        RECT 1408.130 158.480 1408.450 158.540 ;
        RECT 1409.050 158.480 1409.370 158.540 ;
        RECT 1409.050 110.740 1409.370 110.800 ;
        RECT 1408.680 110.600 1409.370 110.740 ;
        RECT 1408.680 110.460 1408.820 110.600 ;
        RECT 1409.050 110.540 1409.370 110.600 ;
        RECT 1408.590 110.200 1408.910 110.460 ;
        RECT 517.110 80.140 517.430 80.200 ;
        RECT 1408.590 80.140 1408.910 80.200 ;
        RECT 517.110 80.000 1408.910 80.140 ;
        RECT 517.110 79.940 517.430 80.000 ;
        RECT 1408.590 79.940 1408.910 80.000 ;
        RECT 513.890 15.540 514.210 15.600 ;
        RECT 517.110 15.540 517.430 15.600 ;
        RECT 513.890 15.400 517.430 15.540 ;
        RECT 513.890 15.340 514.210 15.400 ;
        RECT 517.110 15.340 517.430 15.400 ;
      LAYER via ;
        RECT 1409.080 1497.060 1409.340 1497.320 ;
        RECT 1408.160 1449.120 1408.420 1449.380 ;
        RECT 1408.620 1400.840 1408.880 1401.100 ;
        RECT 1409.540 1400.840 1409.800 1401.100 ;
        RECT 1410.000 1296.800 1410.260 1297.060 ;
        RECT 1409.540 1207.720 1409.800 1207.980 ;
        RECT 1409.540 1207.040 1409.800 1207.300 ;
        RECT 1409.540 1172.700 1409.800 1172.960 ;
        RECT 1409.540 1110.820 1409.800 1111.080 ;
        RECT 1409.540 1104.020 1409.800 1104.280 ;
        RECT 1409.540 1076.820 1409.800 1077.080 ;
        RECT 1409.540 1076.140 1409.800 1076.400 ;
        RECT 1408.620 1055.400 1408.880 1055.660 ;
        RECT 1409.080 1013.920 1409.340 1014.180 ;
        RECT 1409.540 980.260 1409.800 980.520 ;
        RECT 1409.080 979.580 1409.340 979.840 ;
        RECT 1408.620 834.740 1408.880 835.000 ;
        RECT 1409.540 834.740 1409.800 835.000 ;
        RECT 1409.540 786.800 1409.800 787.060 ;
        RECT 1409.080 786.460 1409.340 786.720 ;
        RECT 1408.160 675.960 1408.420 676.220 ;
        RECT 1409.080 645.020 1409.340 645.280 ;
        RECT 1409.080 531.120 1409.340 531.380 ;
        RECT 1409.540 531.120 1409.800 531.380 ;
        RECT 1409.080 482.840 1409.340 483.100 ;
        RECT 1410.000 482.840 1410.260 483.100 ;
        RECT 1409.080 386.620 1409.340 386.880 ;
        RECT 1410.000 386.620 1410.260 386.880 ;
        RECT 1409.080 362.140 1409.340 362.400 ;
        RECT 1410.000 362.140 1410.260 362.400 ;
        RECT 1408.620 330.860 1408.880 331.120 ;
        RECT 1408.620 282.920 1408.880 283.180 ;
        RECT 1408.620 241.440 1408.880 241.700 ;
        RECT 1409.080 241.440 1409.340 241.700 ;
        RECT 1408.160 193.160 1408.420 193.420 ;
        RECT 1409.080 193.160 1409.340 193.420 ;
        RECT 1408.160 158.480 1408.420 158.740 ;
        RECT 1409.080 158.480 1409.340 158.740 ;
        RECT 1409.080 110.540 1409.340 110.800 ;
        RECT 1408.620 110.200 1408.880 110.460 ;
        RECT 517.140 79.940 517.400 80.200 ;
        RECT 1408.620 79.940 1408.880 80.200 ;
        RECT 513.920 15.340 514.180 15.600 ;
        RECT 517.140 15.340 517.400 15.600 ;
      LAYER met2 ;
        RECT 1413.140 1700.410 1413.420 1702.400 ;
        RECT 1410.980 1700.270 1413.420 1700.410 ;
        RECT 1410.980 1656.210 1411.120 1700.270 ;
        RECT 1413.140 1700.000 1413.420 1700.270 ;
        RECT 1408.220 1656.070 1411.120 1656.210 ;
        RECT 1408.220 1607.250 1408.360 1656.070 ;
        RECT 1408.220 1607.110 1409.280 1607.250 ;
        RECT 1409.140 1546.050 1409.280 1607.110 ;
        RECT 1408.220 1545.910 1409.280 1546.050 ;
        RECT 1408.220 1510.010 1408.360 1545.910 ;
        RECT 1408.220 1509.870 1409.280 1510.010 ;
        RECT 1409.140 1497.350 1409.280 1509.870 ;
        RECT 1409.080 1497.030 1409.340 1497.350 ;
        RECT 1408.160 1449.090 1408.420 1449.410 ;
        RECT 1408.220 1448.925 1408.360 1449.090 ;
        RECT 1408.150 1448.555 1408.430 1448.925 ;
        RECT 1409.530 1448.555 1409.810 1448.925 ;
        RECT 1409.600 1401.130 1409.740 1448.555 ;
        RECT 1408.620 1400.810 1408.880 1401.130 ;
        RECT 1409.540 1400.810 1409.800 1401.130 ;
        RECT 1408.680 1400.645 1408.820 1400.810 ;
        RECT 1408.610 1400.275 1408.890 1400.645 ;
        RECT 1409.070 1399.595 1409.350 1399.965 ;
        RECT 1409.140 1317.570 1409.280 1399.595 ;
        RECT 1408.680 1317.430 1409.280 1317.570 ;
        RECT 1408.680 1303.970 1408.820 1317.430 ;
        RECT 1409.070 1303.970 1409.350 1304.085 ;
        RECT 1408.680 1303.830 1409.350 1303.970 ;
        RECT 1409.070 1303.715 1409.350 1303.830 ;
        RECT 1409.990 1303.715 1410.270 1304.085 ;
        RECT 1410.060 1297.090 1410.200 1303.715 ;
        RECT 1410.000 1296.770 1410.260 1297.090 ;
        RECT 1409.540 1207.690 1409.800 1208.010 ;
        RECT 1409.600 1207.330 1409.740 1207.690 ;
        RECT 1409.540 1207.010 1409.800 1207.330 ;
        RECT 1409.540 1172.670 1409.800 1172.990 ;
        RECT 1409.600 1111.110 1409.740 1172.670 ;
        RECT 1409.540 1110.790 1409.800 1111.110 ;
        RECT 1409.540 1103.990 1409.800 1104.310 ;
        RECT 1409.600 1077.110 1409.740 1103.990 ;
        RECT 1409.540 1076.790 1409.800 1077.110 ;
        RECT 1409.540 1076.110 1409.800 1076.430 ;
        RECT 1409.600 1055.885 1409.740 1076.110 ;
        RECT 1408.610 1055.515 1408.890 1055.885 ;
        RECT 1409.530 1055.515 1409.810 1055.885 ;
        RECT 1408.620 1055.370 1408.880 1055.515 ;
        RECT 1409.080 1013.890 1409.340 1014.210 ;
        RECT 1409.140 1007.490 1409.280 1013.890 ;
        RECT 1409.140 1007.350 1409.740 1007.490 ;
        RECT 1409.600 980.550 1409.740 1007.350 ;
        RECT 1409.540 980.230 1409.800 980.550 ;
        RECT 1409.080 979.550 1409.340 979.870 ;
        RECT 1409.140 931.330 1409.280 979.550 ;
        RECT 1409.140 931.190 1409.740 931.330 ;
        RECT 1409.600 917.730 1409.740 931.190 ;
        RECT 1408.680 917.590 1409.740 917.730 ;
        RECT 1408.680 835.030 1408.820 917.590 ;
        RECT 1408.620 834.710 1408.880 835.030 ;
        RECT 1409.540 834.710 1409.800 835.030 ;
        RECT 1409.600 787.090 1409.740 834.710 ;
        RECT 1409.540 786.770 1409.800 787.090 ;
        RECT 1409.080 786.430 1409.340 786.750 ;
        RECT 1409.140 717.925 1409.280 786.430 ;
        RECT 1408.150 717.555 1408.430 717.925 ;
        RECT 1409.070 717.555 1409.350 717.925 ;
        RECT 1408.220 676.250 1408.360 717.555 ;
        RECT 1408.160 675.930 1408.420 676.250 ;
        RECT 1409.080 644.990 1409.340 645.310 ;
        RECT 1409.140 531.410 1409.280 644.990 ;
        RECT 1409.080 531.090 1409.340 531.410 ;
        RECT 1409.540 531.090 1409.800 531.410 ;
        RECT 1409.600 483.210 1409.740 531.090 ;
        RECT 1409.140 483.130 1409.740 483.210 ;
        RECT 1409.080 483.070 1409.740 483.130 ;
        RECT 1409.080 482.810 1409.340 483.070 ;
        RECT 1410.000 482.810 1410.260 483.130 ;
        RECT 1409.140 482.655 1409.280 482.810 ;
        RECT 1410.060 386.910 1410.200 482.810 ;
        RECT 1409.080 386.590 1409.340 386.910 ;
        RECT 1410.000 386.590 1410.260 386.910 ;
        RECT 1409.140 362.430 1409.280 386.590 ;
        RECT 1409.080 362.110 1409.340 362.430 ;
        RECT 1410.000 362.110 1410.260 362.430 ;
        RECT 1410.060 338.485 1410.200 362.110 ;
        RECT 1409.070 338.370 1409.350 338.485 ;
        RECT 1408.680 338.230 1409.350 338.370 ;
        RECT 1408.680 331.150 1408.820 338.230 ;
        RECT 1409.070 338.115 1409.350 338.230 ;
        RECT 1409.990 338.115 1410.270 338.485 ;
        RECT 1408.620 330.830 1408.880 331.150 ;
        RECT 1408.620 282.890 1408.880 283.210 ;
        RECT 1408.680 241.730 1408.820 282.890 ;
        RECT 1408.620 241.410 1408.880 241.730 ;
        RECT 1409.080 241.410 1409.340 241.730 ;
        RECT 1409.140 193.450 1409.280 241.410 ;
        RECT 1408.160 193.130 1408.420 193.450 ;
        RECT 1409.080 193.130 1409.340 193.450 ;
        RECT 1408.220 158.770 1408.360 193.130 ;
        RECT 1408.160 158.450 1408.420 158.770 ;
        RECT 1409.080 158.450 1409.340 158.770 ;
        RECT 1409.140 110.830 1409.280 158.450 ;
        RECT 1409.080 110.510 1409.340 110.830 ;
        RECT 1408.620 110.170 1408.880 110.490 ;
        RECT 1408.680 80.230 1408.820 110.170 ;
        RECT 517.140 79.910 517.400 80.230 ;
        RECT 1408.620 79.910 1408.880 80.230 ;
        RECT 517.200 15.630 517.340 79.910 ;
        RECT 513.920 15.310 514.180 15.630 ;
        RECT 517.140 15.310 517.400 15.630 ;
        RECT 513.980 2.400 514.120 15.310 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 1408.150 1448.600 1408.430 1448.880 ;
        RECT 1409.530 1448.600 1409.810 1448.880 ;
        RECT 1408.610 1400.320 1408.890 1400.600 ;
        RECT 1409.070 1399.640 1409.350 1399.920 ;
        RECT 1409.070 1303.760 1409.350 1304.040 ;
        RECT 1409.990 1303.760 1410.270 1304.040 ;
        RECT 1408.610 1055.560 1408.890 1055.840 ;
        RECT 1409.530 1055.560 1409.810 1055.840 ;
        RECT 1408.150 717.600 1408.430 717.880 ;
        RECT 1409.070 717.600 1409.350 717.880 ;
        RECT 1409.070 338.160 1409.350 338.440 ;
        RECT 1409.990 338.160 1410.270 338.440 ;
      LAYER met3 ;
        RECT 1408.125 1448.890 1408.455 1448.905 ;
        RECT 1409.505 1448.890 1409.835 1448.905 ;
        RECT 1408.125 1448.590 1409.835 1448.890 ;
        RECT 1408.125 1448.575 1408.455 1448.590 ;
        RECT 1409.505 1448.575 1409.835 1448.590 ;
        RECT 1408.585 1400.610 1408.915 1400.625 ;
        RECT 1407.910 1400.310 1408.915 1400.610 ;
        RECT 1407.910 1399.930 1408.210 1400.310 ;
        RECT 1408.585 1400.295 1408.915 1400.310 ;
        RECT 1409.045 1399.930 1409.375 1399.945 ;
        RECT 1407.910 1399.630 1409.375 1399.930 ;
        RECT 1409.045 1399.615 1409.375 1399.630 ;
        RECT 1409.045 1304.050 1409.375 1304.065 ;
        RECT 1409.965 1304.050 1410.295 1304.065 ;
        RECT 1409.045 1303.750 1410.295 1304.050 ;
        RECT 1409.045 1303.735 1409.375 1303.750 ;
        RECT 1409.965 1303.735 1410.295 1303.750 ;
        RECT 1408.585 1055.850 1408.915 1055.865 ;
        RECT 1409.505 1055.850 1409.835 1055.865 ;
        RECT 1408.585 1055.550 1409.835 1055.850 ;
        RECT 1408.585 1055.535 1408.915 1055.550 ;
        RECT 1409.505 1055.535 1409.835 1055.550 ;
        RECT 1408.125 717.890 1408.455 717.905 ;
        RECT 1409.045 717.890 1409.375 717.905 ;
        RECT 1408.125 717.590 1409.375 717.890 ;
        RECT 1408.125 717.575 1408.455 717.590 ;
        RECT 1409.045 717.575 1409.375 717.590 ;
        RECT 1409.045 338.450 1409.375 338.465 ;
        RECT 1409.965 338.450 1410.295 338.465 ;
        RECT 1409.045 338.150 1410.295 338.450 ;
        RECT 1409.045 338.135 1409.375 338.150 ;
        RECT 1409.965 338.135 1410.295 338.150 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.810 80.480 538.130 80.540 ;
        RECT 1421.930 80.480 1422.250 80.540 ;
        RECT 537.810 80.340 1422.250 80.480 ;
        RECT 537.810 80.280 538.130 80.340 ;
        RECT 1421.930 80.280 1422.250 80.340 ;
        RECT 531.830 15.540 532.150 15.600 ;
        RECT 537.810 15.540 538.130 15.600 ;
        RECT 531.830 15.400 538.130 15.540 ;
        RECT 531.830 15.340 532.150 15.400 ;
        RECT 537.810 15.340 538.130 15.400 ;
      LAYER via ;
        RECT 537.840 80.280 538.100 80.540 ;
        RECT 1421.960 80.280 1422.220 80.540 ;
        RECT 531.860 15.340 532.120 15.600 ;
        RECT 537.840 15.340 538.100 15.600 ;
      LAYER met2 ;
        RECT 1422.340 1700.410 1422.620 1702.400 ;
        RECT 1422.020 1700.270 1422.620 1700.410 ;
        RECT 1422.020 80.570 1422.160 1700.270 ;
        RECT 1422.340 1700.000 1422.620 1700.270 ;
        RECT 537.840 80.250 538.100 80.570 ;
        RECT 1421.960 80.250 1422.220 80.570 ;
        RECT 537.900 15.630 538.040 80.250 ;
        RECT 531.860 15.310 532.120 15.630 ;
        RECT 537.840 15.310 538.100 15.630 ;
        RECT 531.920 2.400 532.060 15.310 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 80.820 551.930 80.880 ;
        RECT 1428.830 80.820 1429.150 80.880 ;
        RECT 551.610 80.680 1429.150 80.820 ;
        RECT 551.610 80.620 551.930 80.680 ;
        RECT 1428.830 80.620 1429.150 80.680 ;
      LAYER via ;
        RECT 551.640 80.620 551.900 80.880 ;
        RECT 1428.860 80.620 1429.120 80.880 ;
      LAYER met2 ;
        RECT 1431.540 1700.410 1431.820 1702.400 ;
        RECT 1428.920 1700.270 1431.820 1700.410 ;
        RECT 1428.920 80.910 1429.060 1700.270 ;
        RECT 1431.540 1700.000 1431.820 1700.270 ;
        RECT 551.640 80.590 551.900 80.910 ;
        RECT 1428.860 80.590 1429.120 80.910 ;
        RECT 551.700 16.730 551.840 80.590 ;
        RECT 549.860 16.590 551.840 16.730 ;
        RECT 549.860 2.400 550.000 16.590 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1436.265 1400.885 1436.435 1448.995 ;
        RECT 1436.265 1304.325 1436.435 1352.435 ;
        RECT 1436.265 1207.425 1436.435 1255.875 ;
      LAYER mcon ;
        RECT 1436.265 1448.825 1436.435 1448.995 ;
        RECT 1436.265 1352.265 1436.435 1352.435 ;
        RECT 1436.265 1255.705 1436.435 1255.875 ;
      LAYER met1 ;
        RECT 1435.730 1545.880 1436.050 1545.940 ;
        RECT 1436.190 1545.880 1436.510 1545.940 ;
        RECT 1435.730 1545.740 1436.510 1545.880 ;
        RECT 1435.730 1545.680 1436.050 1545.740 ;
        RECT 1436.190 1545.680 1436.510 1545.740 ;
        RECT 1436.190 1448.980 1436.510 1449.040 ;
        RECT 1435.995 1448.840 1436.510 1448.980 ;
        RECT 1436.190 1448.780 1436.510 1448.840 ;
        RECT 1436.190 1401.040 1436.510 1401.100 ;
        RECT 1435.995 1400.900 1436.510 1401.040 ;
        RECT 1436.190 1400.840 1436.510 1400.900 ;
        RECT 1436.190 1352.420 1436.510 1352.480 ;
        RECT 1435.995 1352.280 1436.510 1352.420 ;
        RECT 1436.190 1352.220 1436.510 1352.280 ;
        RECT 1436.190 1304.480 1436.510 1304.540 ;
        RECT 1435.995 1304.340 1436.510 1304.480 ;
        RECT 1436.190 1304.280 1436.510 1304.340 ;
        RECT 1436.190 1255.860 1436.510 1255.920 ;
        RECT 1435.995 1255.720 1436.510 1255.860 ;
        RECT 1436.190 1255.660 1436.510 1255.720 ;
        RECT 1436.190 1207.580 1436.510 1207.640 ;
        RECT 1435.995 1207.440 1436.510 1207.580 ;
        RECT 1436.190 1207.380 1436.510 1207.440 ;
        RECT 1436.190 1111.020 1436.510 1111.080 ;
        RECT 1437.110 1111.020 1437.430 1111.080 ;
        RECT 1436.190 1110.880 1437.430 1111.020 ;
        RECT 1436.190 1110.820 1436.510 1110.880 ;
        RECT 1437.110 1110.820 1437.430 1110.880 ;
        RECT 1436.190 917.900 1436.510 917.960 ;
        RECT 1437.110 917.900 1437.430 917.960 ;
        RECT 1436.190 917.760 1437.430 917.900 ;
        RECT 1436.190 917.700 1436.510 917.760 ;
        RECT 1437.110 917.700 1437.430 917.760 ;
        RECT 1436.190 796.860 1436.510 796.920 ;
        RECT 1437.110 796.860 1437.430 796.920 ;
        RECT 1436.190 796.720 1437.430 796.860 ;
        RECT 1436.190 796.660 1436.510 796.720 ;
        RECT 1437.110 796.660 1437.430 796.720 ;
        RECT 1435.730 386.480 1436.050 386.540 ;
        RECT 1436.190 386.480 1436.510 386.540 ;
        RECT 1435.730 386.340 1436.510 386.480 ;
        RECT 1435.730 386.280 1436.050 386.340 ;
        RECT 1436.190 386.280 1436.510 386.340 ;
        RECT 572.310 81.160 572.630 81.220 ;
        RECT 1436.190 81.160 1436.510 81.220 ;
        RECT 572.310 81.020 1436.510 81.160 ;
        RECT 572.310 80.960 572.630 81.020 ;
        RECT 1436.190 80.960 1436.510 81.020 ;
        RECT 567.710 14.860 568.030 14.920 ;
        RECT 572.310 14.860 572.630 14.920 ;
        RECT 567.710 14.720 572.630 14.860 ;
        RECT 567.710 14.660 568.030 14.720 ;
        RECT 572.310 14.660 572.630 14.720 ;
      LAYER via ;
        RECT 1435.760 1545.680 1436.020 1545.940 ;
        RECT 1436.220 1545.680 1436.480 1545.940 ;
        RECT 1436.220 1448.780 1436.480 1449.040 ;
        RECT 1436.220 1400.840 1436.480 1401.100 ;
        RECT 1436.220 1352.220 1436.480 1352.480 ;
        RECT 1436.220 1304.280 1436.480 1304.540 ;
        RECT 1436.220 1255.660 1436.480 1255.920 ;
        RECT 1436.220 1207.380 1436.480 1207.640 ;
        RECT 1436.220 1110.820 1436.480 1111.080 ;
        RECT 1437.140 1110.820 1437.400 1111.080 ;
        RECT 1436.220 917.700 1436.480 917.960 ;
        RECT 1437.140 917.700 1437.400 917.960 ;
        RECT 1436.220 796.660 1436.480 796.920 ;
        RECT 1437.140 796.660 1437.400 796.920 ;
        RECT 1435.760 386.280 1436.020 386.540 ;
        RECT 1436.220 386.280 1436.480 386.540 ;
        RECT 572.340 80.960 572.600 81.220 ;
        RECT 1436.220 80.960 1436.480 81.220 ;
        RECT 567.740 14.660 568.000 14.920 ;
        RECT 572.340 14.660 572.600 14.920 ;
      LAYER met2 ;
        RECT 1440.740 1700.410 1441.020 1702.400 ;
        RECT 1438.580 1700.270 1441.020 1700.410 ;
        RECT 1438.580 1689.530 1438.720 1700.270 ;
        RECT 1440.740 1700.000 1441.020 1700.270 ;
        RECT 1436.280 1689.390 1438.720 1689.530 ;
        RECT 1436.280 1618.130 1436.420 1689.390 ;
        RECT 1435.820 1617.990 1436.420 1618.130 ;
        RECT 1435.820 1545.970 1435.960 1617.990 ;
        RECT 1435.760 1545.650 1436.020 1545.970 ;
        RECT 1436.220 1545.650 1436.480 1545.970 ;
        RECT 1436.280 1449.070 1436.420 1545.650 ;
        RECT 1436.220 1448.750 1436.480 1449.070 ;
        RECT 1436.220 1400.810 1436.480 1401.130 ;
        RECT 1436.280 1352.510 1436.420 1400.810 ;
        RECT 1436.220 1352.190 1436.480 1352.510 ;
        RECT 1436.220 1304.250 1436.480 1304.570 ;
        RECT 1436.280 1255.950 1436.420 1304.250 ;
        RECT 1436.220 1255.630 1436.480 1255.950 ;
        RECT 1436.220 1207.350 1436.480 1207.670 ;
        RECT 1436.280 1159.245 1436.420 1207.350 ;
        RECT 1436.210 1158.875 1436.490 1159.245 ;
        RECT 1437.130 1158.875 1437.410 1159.245 ;
        RECT 1437.200 1111.110 1437.340 1158.875 ;
        RECT 1436.220 1110.790 1436.480 1111.110 ;
        RECT 1437.140 1110.790 1437.400 1111.110 ;
        RECT 1436.280 966.125 1436.420 1110.790 ;
        RECT 1436.210 965.755 1436.490 966.125 ;
        RECT 1437.130 965.755 1437.410 966.125 ;
        RECT 1437.200 917.990 1437.340 965.755 ;
        RECT 1436.220 917.670 1436.480 917.990 ;
        RECT 1437.140 917.670 1437.400 917.990 ;
        RECT 1436.280 796.950 1436.420 917.670 ;
        RECT 1436.220 796.630 1436.480 796.950 ;
        RECT 1437.140 796.630 1437.400 796.950 ;
        RECT 1437.200 773.005 1437.340 796.630 ;
        RECT 1436.210 772.635 1436.490 773.005 ;
        RECT 1437.130 772.635 1437.410 773.005 ;
        RECT 1436.280 700.810 1436.420 772.635 ;
        RECT 1436.280 700.670 1436.880 700.810 ;
        RECT 1436.740 699.450 1436.880 700.670 ;
        RECT 1436.280 699.310 1436.880 699.450 ;
        RECT 1436.280 400.080 1436.420 699.310 ;
        RECT 1435.820 399.940 1436.420 400.080 ;
        RECT 1435.820 386.570 1435.960 399.940 ;
        RECT 1435.760 386.250 1436.020 386.570 ;
        RECT 1436.220 386.250 1436.480 386.570 ;
        RECT 1436.280 218.010 1436.420 386.250 ;
        RECT 1436.280 217.870 1436.880 218.010 ;
        RECT 1436.740 216.650 1436.880 217.870 ;
        RECT 1436.280 216.510 1436.880 216.650 ;
        RECT 1436.280 81.250 1436.420 216.510 ;
        RECT 572.340 80.930 572.600 81.250 ;
        RECT 1436.220 80.930 1436.480 81.250 ;
        RECT 572.400 14.950 572.540 80.930 ;
        RECT 567.740 14.630 568.000 14.950 ;
        RECT 572.340 14.630 572.600 14.950 ;
        RECT 567.800 2.400 567.940 14.630 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1436.210 1158.920 1436.490 1159.200 ;
        RECT 1437.130 1158.920 1437.410 1159.200 ;
        RECT 1436.210 965.800 1436.490 966.080 ;
        RECT 1437.130 965.800 1437.410 966.080 ;
        RECT 1436.210 772.680 1436.490 772.960 ;
        RECT 1437.130 772.680 1437.410 772.960 ;
      LAYER met3 ;
        RECT 1436.185 1159.210 1436.515 1159.225 ;
        RECT 1437.105 1159.210 1437.435 1159.225 ;
        RECT 1436.185 1158.910 1437.435 1159.210 ;
        RECT 1436.185 1158.895 1436.515 1158.910 ;
        RECT 1437.105 1158.895 1437.435 1158.910 ;
        RECT 1436.185 966.090 1436.515 966.105 ;
        RECT 1437.105 966.090 1437.435 966.105 ;
        RECT 1436.185 965.790 1437.435 966.090 ;
        RECT 1436.185 965.775 1436.515 965.790 ;
        RECT 1437.105 965.775 1437.435 965.790 ;
        RECT 1436.185 772.970 1436.515 772.985 ;
        RECT 1437.105 772.970 1437.435 772.985 ;
        RECT 1436.185 772.670 1437.435 772.970 ;
        RECT 1436.185 772.655 1436.515 772.670 ;
        RECT 1437.105 772.655 1437.435 772.670 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1449.990 1688.000 1450.310 1688.060 ;
        RECT 1242.160 1687.860 1450.310 1688.000 ;
        RECT 1231.490 1687.660 1231.810 1687.720 ;
        RECT 1242.160 1687.660 1242.300 1687.860 ;
        RECT 1449.990 1687.800 1450.310 1687.860 ;
        RECT 1231.490 1687.520 1242.300 1687.660 ;
        RECT 1231.490 1687.460 1231.810 1687.520 ;
        RECT 586.110 70.620 586.430 70.680 ;
        RECT 1231.490 70.620 1231.810 70.680 ;
        RECT 586.110 70.480 1231.810 70.620 ;
        RECT 586.110 70.420 586.430 70.480 ;
        RECT 1231.490 70.420 1231.810 70.480 ;
      LAYER via ;
        RECT 1231.520 1687.460 1231.780 1687.720 ;
        RECT 1450.020 1687.800 1450.280 1688.060 ;
        RECT 586.140 70.420 586.400 70.680 ;
        RECT 1231.520 70.420 1231.780 70.680 ;
      LAYER met2 ;
        RECT 1449.940 1700.000 1450.220 1702.400 ;
        RECT 1450.080 1688.090 1450.220 1700.000 ;
        RECT 1450.020 1687.770 1450.280 1688.090 ;
        RECT 1231.520 1687.430 1231.780 1687.750 ;
        RECT 1231.580 70.710 1231.720 1687.430 ;
        RECT 586.140 70.390 586.400 70.710 ;
        RECT 1231.520 70.390 1231.780 70.710 ;
        RECT 586.200 17.410 586.340 70.390 ;
        RECT 585.740 17.270 586.340 17.410 ;
        RECT 585.740 2.400 585.880 17.270 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 96.210 65.520 96.530 65.580 ;
        RECT 1194.230 65.520 1194.550 65.580 ;
        RECT 96.210 65.380 1194.550 65.520 ;
        RECT 96.210 65.320 96.530 65.380 ;
        RECT 1194.230 65.320 1194.550 65.380 ;
        RECT 91.610 17.920 91.930 17.980 ;
        RECT 96.210 17.920 96.530 17.980 ;
        RECT 91.610 17.780 96.530 17.920 ;
        RECT 91.610 17.720 91.930 17.780 ;
        RECT 96.210 17.720 96.530 17.780 ;
      LAYER via ;
        RECT 96.240 65.320 96.500 65.580 ;
        RECT 1194.260 65.320 1194.520 65.580 ;
        RECT 91.640 17.720 91.900 17.980 ;
        RECT 96.240 17.720 96.500 17.980 ;
      LAYER met2 ;
        RECT 1195.560 1700.410 1195.840 1702.400 ;
        RECT 1194.320 1700.270 1195.840 1700.410 ;
        RECT 1194.320 65.610 1194.460 1700.270 ;
        RECT 1195.560 1700.000 1195.840 1700.270 ;
        RECT 96.240 65.290 96.500 65.610 ;
        RECT 1194.260 65.290 1194.520 65.610 ;
        RECT 96.300 18.010 96.440 65.290 ;
        RECT 91.640 17.690 91.900 18.010 ;
        RECT 96.240 17.690 96.500 18.010 ;
        RECT 91.700 2.400 91.840 17.690 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 81.500 607.130 81.560 ;
        RECT 1456.430 81.500 1456.750 81.560 ;
        RECT 606.810 81.360 1456.750 81.500 ;
        RECT 606.810 81.300 607.130 81.360 ;
        RECT 1456.430 81.300 1456.750 81.360 ;
        RECT 603.130 14.860 603.450 14.920 ;
        RECT 606.810 14.860 607.130 14.920 ;
        RECT 603.130 14.720 607.130 14.860 ;
        RECT 603.130 14.660 603.450 14.720 ;
        RECT 606.810 14.660 607.130 14.720 ;
      LAYER via ;
        RECT 606.840 81.300 607.100 81.560 ;
        RECT 1456.460 81.300 1456.720 81.560 ;
        RECT 603.160 14.660 603.420 14.920 ;
        RECT 606.840 14.660 607.100 14.920 ;
      LAYER met2 ;
        RECT 1459.140 1700.410 1459.420 1702.400 ;
        RECT 1456.520 1700.270 1459.420 1700.410 ;
        RECT 1456.520 81.590 1456.660 1700.270 ;
        RECT 1459.140 1700.000 1459.420 1700.270 ;
        RECT 606.840 81.270 607.100 81.590 ;
        RECT 1456.460 81.270 1456.720 81.590 ;
        RECT 606.900 14.950 607.040 81.270 ;
        RECT 603.160 14.630 603.420 14.950 ;
        RECT 606.840 14.630 607.100 14.950 ;
        RECT 603.220 2.400 603.360 14.630 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1463.865 1587.205 1464.035 1635.315 ;
        RECT 1463.865 1490.985 1464.035 1538.755 ;
        RECT 1463.405 1442.025 1463.575 1490.475 ;
        RECT 1464.785 1248.565 1464.955 1290.215 ;
        RECT 1463.865 904.145 1464.035 993.395 ;
        RECT 1463.865 710.685 1464.035 758.795 ;
        RECT 1463.865 517.905 1464.035 565.675 ;
        RECT 1463.405 469.285 1463.575 517.395 ;
        RECT 1463.865 227.885 1464.035 275.995 ;
        RECT 1463.865 179.605 1464.035 185.895 ;
      LAYER mcon ;
        RECT 1463.865 1635.145 1464.035 1635.315 ;
        RECT 1463.865 1538.585 1464.035 1538.755 ;
        RECT 1463.405 1490.305 1463.575 1490.475 ;
        RECT 1464.785 1290.045 1464.955 1290.215 ;
        RECT 1463.865 993.225 1464.035 993.395 ;
        RECT 1463.865 758.625 1464.035 758.795 ;
        RECT 1463.865 565.505 1464.035 565.675 ;
        RECT 1463.405 517.225 1463.575 517.395 ;
        RECT 1463.865 275.825 1464.035 275.995 ;
        RECT 1463.865 185.725 1464.035 185.895 ;
      LAYER met1 ;
        RECT 1463.790 1645.160 1464.110 1645.220 ;
        RECT 1466.090 1645.160 1466.410 1645.220 ;
        RECT 1463.790 1645.020 1466.410 1645.160 ;
        RECT 1463.790 1644.960 1464.110 1645.020 ;
        RECT 1466.090 1644.960 1466.410 1645.020 ;
        RECT 1463.790 1635.300 1464.110 1635.360 ;
        RECT 1463.595 1635.160 1464.110 1635.300 ;
        RECT 1463.790 1635.100 1464.110 1635.160 ;
        RECT 1463.790 1587.360 1464.110 1587.420 ;
        RECT 1463.595 1587.220 1464.110 1587.360 ;
        RECT 1463.790 1587.160 1464.110 1587.220 ;
        RECT 1463.790 1538.740 1464.110 1538.800 ;
        RECT 1463.595 1538.600 1464.110 1538.740 ;
        RECT 1463.790 1538.540 1464.110 1538.600 ;
        RECT 1463.790 1491.140 1464.110 1491.200 ;
        RECT 1463.595 1491.000 1464.110 1491.140 ;
        RECT 1463.790 1490.940 1464.110 1491.000 ;
        RECT 1463.345 1490.460 1463.635 1490.505 ;
        RECT 1463.790 1490.460 1464.110 1490.520 ;
        RECT 1463.345 1490.320 1464.110 1490.460 ;
        RECT 1463.345 1490.275 1463.635 1490.320 ;
        RECT 1463.790 1490.260 1464.110 1490.320 ;
        RECT 1463.330 1442.180 1463.650 1442.240 ;
        RECT 1463.135 1442.040 1463.650 1442.180 ;
        RECT 1463.330 1441.980 1463.650 1442.040 ;
        RECT 1463.330 1401.040 1463.650 1401.100 ;
        RECT 1463.790 1401.040 1464.110 1401.100 ;
        RECT 1463.330 1400.900 1464.110 1401.040 ;
        RECT 1463.330 1400.840 1463.650 1400.900 ;
        RECT 1463.790 1400.840 1464.110 1400.900 ;
        RECT 1463.790 1304.280 1464.110 1304.540 ;
        RECT 1463.880 1303.860 1464.020 1304.280 ;
        RECT 1463.790 1303.600 1464.110 1303.860 ;
        RECT 1464.250 1290.200 1464.570 1290.260 ;
        RECT 1464.725 1290.200 1465.015 1290.245 ;
        RECT 1464.250 1290.060 1465.015 1290.200 ;
        RECT 1464.250 1290.000 1464.570 1290.060 ;
        RECT 1464.725 1290.015 1465.015 1290.060 ;
        RECT 1464.250 1248.720 1464.570 1248.780 ;
        RECT 1464.725 1248.720 1465.015 1248.765 ;
        RECT 1464.250 1248.580 1465.015 1248.720 ;
        RECT 1464.250 1248.520 1464.570 1248.580 ;
        RECT 1464.725 1248.535 1465.015 1248.580 ;
        RECT 1463.790 1200.780 1464.110 1200.840 ;
        RECT 1464.250 1200.780 1464.570 1200.840 ;
        RECT 1463.790 1200.640 1464.570 1200.780 ;
        RECT 1463.790 1200.580 1464.110 1200.640 ;
        RECT 1464.250 1200.580 1464.570 1200.640 ;
        RECT 1463.790 1152.840 1464.110 1152.900 ;
        RECT 1464.250 1152.840 1464.570 1152.900 ;
        RECT 1463.790 1152.700 1464.570 1152.840 ;
        RECT 1463.790 1152.640 1464.110 1152.700 ;
        RECT 1464.250 1152.640 1464.570 1152.700 ;
        RECT 1463.790 1000.520 1464.110 1000.580 ;
        RECT 1464.250 1000.520 1464.570 1000.580 ;
        RECT 1463.790 1000.380 1464.570 1000.520 ;
        RECT 1463.790 1000.320 1464.110 1000.380 ;
        RECT 1464.250 1000.320 1464.570 1000.380 ;
        RECT 1463.805 993.380 1464.095 993.425 ;
        RECT 1464.250 993.380 1464.570 993.440 ;
        RECT 1463.805 993.240 1464.570 993.380 ;
        RECT 1463.805 993.195 1464.095 993.240 ;
        RECT 1464.250 993.180 1464.570 993.240 ;
        RECT 1463.790 904.300 1464.110 904.360 ;
        RECT 1463.595 904.160 1464.110 904.300 ;
        RECT 1463.790 904.100 1464.110 904.160 ;
        RECT 1463.790 856.160 1464.110 856.420 ;
        RECT 1463.880 855.740 1464.020 856.160 ;
        RECT 1463.790 855.480 1464.110 855.740 ;
        RECT 1463.790 758.780 1464.110 758.840 ;
        RECT 1463.595 758.640 1464.110 758.780 ;
        RECT 1463.790 758.580 1464.110 758.640 ;
        RECT 1463.790 710.840 1464.110 710.900 ;
        RECT 1463.595 710.700 1464.110 710.840 ;
        RECT 1463.790 710.640 1464.110 710.700 ;
        RECT 1463.790 565.660 1464.110 565.720 ;
        RECT 1463.595 565.520 1464.110 565.660 ;
        RECT 1463.790 565.460 1464.110 565.520 ;
        RECT 1463.790 518.060 1464.110 518.120 ;
        RECT 1463.595 517.920 1464.110 518.060 ;
        RECT 1463.790 517.860 1464.110 517.920 ;
        RECT 1463.345 517.380 1463.635 517.425 ;
        RECT 1463.790 517.380 1464.110 517.440 ;
        RECT 1463.345 517.240 1464.110 517.380 ;
        RECT 1463.345 517.195 1463.635 517.240 ;
        RECT 1463.790 517.180 1464.110 517.240 ;
        RECT 1463.330 469.440 1463.650 469.500 ;
        RECT 1463.135 469.300 1463.650 469.440 ;
        RECT 1463.330 469.240 1463.650 469.300 ;
        RECT 1463.790 345.140 1464.110 345.400 ;
        RECT 1463.880 344.720 1464.020 345.140 ;
        RECT 1463.790 344.460 1464.110 344.720 ;
        RECT 1462.410 324.260 1462.730 324.320 ;
        RECT 1463.790 324.260 1464.110 324.320 ;
        RECT 1462.410 324.120 1464.110 324.260 ;
        RECT 1462.410 324.060 1462.730 324.120 ;
        RECT 1463.790 324.060 1464.110 324.120 ;
        RECT 1463.790 275.980 1464.110 276.040 ;
        RECT 1463.595 275.840 1464.110 275.980 ;
        RECT 1463.790 275.780 1464.110 275.840 ;
        RECT 1463.805 228.040 1464.095 228.085 ;
        RECT 1464.710 228.040 1465.030 228.100 ;
        RECT 1463.805 227.900 1465.030 228.040 ;
        RECT 1463.805 227.855 1464.095 227.900 ;
        RECT 1464.710 227.840 1465.030 227.900 ;
        RECT 1463.805 185.880 1464.095 185.925 ;
        RECT 1464.710 185.880 1465.030 185.940 ;
        RECT 1463.805 185.740 1465.030 185.880 ;
        RECT 1463.805 185.695 1464.095 185.740 ;
        RECT 1464.710 185.680 1465.030 185.740 ;
        RECT 1463.790 179.760 1464.110 179.820 ;
        RECT 1463.595 179.620 1464.110 179.760 ;
        RECT 1463.790 179.560 1464.110 179.620 ;
        RECT 1463.790 144.740 1464.110 144.800 ;
        RECT 1464.250 144.740 1464.570 144.800 ;
        RECT 1463.790 144.600 1464.570 144.740 ;
        RECT 1463.790 144.540 1464.110 144.600 ;
        RECT 1464.250 144.540 1464.570 144.600 ;
        RECT 627.050 81.840 627.370 81.900 ;
        RECT 1463.790 81.840 1464.110 81.900 ;
        RECT 627.050 81.700 1464.110 81.840 ;
        RECT 627.050 81.640 627.370 81.700 ;
        RECT 1463.790 81.640 1464.110 81.700 ;
        RECT 621.070 20.980 621.390 21.040 ;
        RECT 627.050 20.980 627.370 21.040 ;
        RECT 621.070 20.840 627.370 20.980 ;
        RECT 621.070 20.780 621.390 20.840 ;
        RECT 627.050 20.780 627.370 20.840 ;
      LAYER via ;
        RECT 1463.820 1644.960 1464.080 1645.220 ;
        RECT 1466.120 1644.960 1466.380 1645.220 ;
        RECT 1463.820 1635.100 1464.080 1635.360 ;
        RECT 1463.820 1587.160 1464.080 1587.420 ;
        RECT 1463.820 1538.540 1464.080 1538.800 ;
        RECT 1463.820 1490.940 1464.080 1491.200 ;
        RECT 1463.820 1490.260 1464.080 1490.520 ;
        RECT 1463.360 1441.980 1463.620 1442.240 ;
        RECT 1463.360 1400.840 1463.620 1401.100 ;
        RECT 1463.820 1400.840 1464.080 1401.100 ;
        RECT 1463.820 1304.280 1464.080 1304.540 ;
        RECT 1463.820 1303.600 1464.080 1303.860 ;
        RECT 1464.280 1290.000 1464.540 1290.260 ;
        RECT 1464.280 1248.520 1464.540 1248.780 ;
        RECT 1463.820 1200.580 1464.080 1200.840 ;
        RECT 1464.280 1200.580 1464.540 1200.840 ;
        RECT 1463.820 1152.640 1464.080 1152.900 ;
        RECT 1464.280 1152.640 1464.540 1152.900 ;
        RECT 1463.820 1000.320 1464.080 1000.580 ;
        RECT 1464.280 1000.320 1464.540 1000.580 ;
        RECT 1464.280 993.180 1464.540 993.440 ;
        RECT 1463.820 904.100 1464.080 904.360 ;
        RECT 1463.820 856.160 1464.080 856.420 ;
        RECT 1463.820 855.480 1464.080 855.740 ;
        RECT 1463.820 758.580 1464.080 758.840 ;
        RECT 1463.820 710.640 1464.080 710.900 ;
        RECT 1463.820 565.460 1464.080 565.720 ;
        RECT 1463.820 517.860 1464.080 518.120 ;
        RECT 1463.820 517.180 1464.080 517.440 ;
        RECT 1463.360 469.240 1463.620 469.500 ;
        RECT 1463.820 345.140 1464.080 345.400 ;
        RECT 1463.820 344.460 1464.080 344.720 ;
        RECT 1462.440 324.060 1462.700 324.320 ;
        RECT 1463.820 324.060 1464.080 324.320 ;
        RECT 1463.820 275.780 1464.080 276.040 ;
        RECT 1464.740 227.840 1465.000 228.100 ;
        RECT 1464.740 185.680 1465.000 185.940 ;
        RECT 1463.820 179.560 1464.080 179.820 ;
        RECT 1463.820 144.540 1464.080 144.800 ;
        RECT 1464.280 144.540 1464.540 144.800 ;
        RECT 627.080 81.640 627.340 81.900 ;
        RECT 1463.820 81.640 1464.080 81.900 ;
        RECT 621.100 20.780 621.360 21.040 ;
        RECT 627.080 20.780 627.340 21.040 ;
      LAYER met2 ;
        RECT 1468.340 1700.410 1468.620 1702.400 ;
        RECT 1466.180 1700.270 1468.620 1700.410 ;
        RECT 1466.180 1645.250 1466.320 1700.270 ;
        RECT 1468.340 1700.000 1468.620 1700.270 ;
        RECT 1463.820 1644.930 1464.080 1645.250 ;
        RECT 1466.120 1644.930 1466.380 1645.250 ;
        RECT 1463.880 1635.390 1464.020 1644.930 ;
        RECT 1463.820 1635.070 1464.080 1635.390 ;
        RECT 1463.820 1587.130 1464.080 1587.450 ;
        RECT 1463.880 1538.830 1464.020 1587.130 ;
        RECT 1463.820 1538.510 1464.080 1538.830 ;
        RECT 1463.820 1490.910 1464.080 1491.230 ;
        RECT 1463.880 1490.550 1464.020 1490.910 ;
        RECT 1463.820 1490.230 1464.080 1490.550 ;
        RECT 1463.360 1441.950 1463.620 1442.270 ;
        RECT 1463.420 1401.130 1463.560 1441.950 ;
        RECT 1463.360 1400.810 1463.620 1401.130 ;
        RECT 1463.820 1400.810 1464.080 1401.130 ;
        RECT 1463.880 1304.570 1464.020 1400.810 ;
        RECT 1463.820 1304.250 1464.080 1304.570 ;
        RECT 1463.820 1303.570 1464.080 1303.890 ;
        RECT 1463.880 1297.170 1464.020 1303.570 ;
        RECT 1463.880 1297.030 1464.480 1297.170 ;
        RECT 1464.340 1290.290 1464.480 1297.030 ;
        RECT 1464.280 1289.970 1464.540 1290.290 ;
        RECT 1464.280 1248.490 1464.540 1248.810 ;
        RECT 1464.340 1200.870 1464.480 1248.490 ;
        RECT 1463.820 1200.550 1464.080 1200.870 ;
        RECT 1464.280 1200.550 1464.540 1200.870 ;
        RECT 1463.880 1177.490 1464.020 1200.550 ;
        RECT 1463.880 1177.350 1464.480 1177.490 ;
        RECT 1464.340 1152.930 1464.480 1177.350 ;
        RECT 1463.820 1152.610 1464.080 1152.930 ;
        RECT 1464.280 1152.610 1464.540 1152.930 ;
        RECT 1463.880 1000.610 1464.020 1152.610 ;
        RECT 1463.820 1000.290 1464.080 1000.610 ;
        RECT 1464.280 1000.290 1464.540 1000.610 ;
        RECT 1464.340 993.470 1464.480 1000.290 ;
        RECT 1464.280 993.150 1464.540 993.470 ;
        RECT 1463.820 904.070 1464.080 904.390 ;
        RECT 1463.880 856.450 1464.020 904.070 ;
        RECT 1463.820 856.130 1464.080 856.450 ;
        RECT 1463.820 855.450 1464.080 855.770 ;
        RECT 1463.880 758.870 1464.020 855.450 ;
        RECT 1463.820 758.550 1464.080 758.870 ;
        RECT 1463.820 710.610 1464.080 710.930 ;
        RECT 1463.880 565.750 1464.020 710.610 ;
        RECT 1463.820 565.430 1464.080 565.750 ;
        RECT 1463.820 517.830 1464.080 518.150 ;
        RECT 1463.880 517.470 1464.020 517.830 ;
        RECT 1463.820 517.150 1464.080 517.470 ;
        RECT 1463.360 469.210 1463.620 469.530 ;
        RECT 1463.420 426.770 1463.560 469.210 ;
        RECT 1463.420 426.630 1464.020 426.770 ;
        RECT 1463.880 345.430 1464.020 426.630 ;
        RECT 1463.820 345.110 1464.080 345.430 ;
        RECT 1463.820 344.430 1464.080 344.750 ;
        RECT 1463.880 324.350 1464.020 344.430 ;
        RECT 1462.440 324.030 1462.700 324.350 ;
        RECT 1463.820 324.030 1464.080 324.350 ;
        RECT 1462.500 276.605 1462.640 324.030 ;
        RECT 1462.430 276.235 1462.710 276.605 ;
        RECT 1463.810 276.235 1464.090 276.605 ;
        RECT 1463.880 276.070 1464.020 276.235 ;
        RECT 1463.820 275.750 1464.080 276.070 ;
        RECT 1464.740 227.810 1465.000 228.130 ;
        RECT 1464.800 185.970 1464.940 227.810 ;
        RECT 1464.740 185.650 1465.000 185.970 ;
        RECT 1463.820 179.530 1464.080 179.850 ;
        RECT 1463.880 169.050 1464.020 179.530 ;
        RECT 1463.880 168.910 1464.940 169.050 ;
        RECT 1464.800 158.170 1464.940 168.910 ;
        RECT 1464.340 158.030 1464.940 158.170 ;
        RECT 1464.340 144.830 1464.480 158.030 ;
        RECT 1463.820 144.510 1464.080 144.830 ;
        RECT 1464.280 144.510 1464.540 144.830 ;
        RECT 1463.880 81.930 1464.020 144.510 ;
        RECT 627.080 81.610 627.340 81.930 ;
        RECT 1463.820 81.610 1464.080 81.930 ;
        RECT 627.140 21.070 627.280 81.610 ;
        RECT 621.100 20.750 621.360 21.070 ;
        RECT 627.080 20.750 627.340 21.070 ;
        RECT 621.160 2.400 621.300 20.750 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 1462.430 276.280 1462.710 276.560 ;
        RECT 1463.810 276.280 1464.090 276.560 ;
      LAYER met3 ;
        RECT 1462.405 276.570 1462.735 276.585 ;
        RECT 1463.785 276.570 1464.115 276.585 ;
        RECT 1462.405 276.270 1464.115 276.570 ;
        RECT 1462.405 276.255 1462.735 276.270 ;
        RECT 1463.785 276.255 1464.115 276.270 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 72.320 117.230 72.380 ;
        RECT 1208.490 72.320 1208.810 72.380 ;
        RECT 116.910 72.180 1208.810 72.320 ;
        RECT 116.910 72.120 117.230 72.180 ;
        RECT 1208.490 72.120 1208.810 72.180 ;
      LAYER via ;
        RECT 116.940 72.120 117.200 72.380 ;
        RECT 1208.520 72.120 1208.780 72.380 ;
      LAYER met2 ;
        RECT 1207.980 1700.410 1208.260 1702.400 ;
        RECT 1207.980 1700.270 1208.720 1700.410 ;
        RECT 1207.980 1700.000 1208.260 1700.270 ;
        RECT 1208.580 72.410 1208.720 1700.270 ;
        RECT 116.940 72.090 117.200 72.410 ;
        RECT 1208.520 72.090 1208.780 72.410 ;
        RECT 117.000 17.410 117.140 72.090 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1215.005 1490.645 1215.175 1538.755 ;
        RECT 1215.925 1121.065 1216.095 1158.635 ;
        RECT 1215.465 1007.165 1215.635 1089.955 ;
        RECT 1215.465 807.245 1215.635 855.355 ;
        RECT 1215.465 620.925 1215.635 669.375 ;
        RECT 1215.925 483.565 1216.095 530.995 ;
        RECT 1215.005 276.165 1215.175 324.275 ;
        RECT 1215.005 179.605 1215.175 227.715 ;
      LAYER mcon ;
        RECT 1215.005 1538.585 1215.175 1538.755 ;
        RECT 1215.925 1158.465 1216.095 1158.635 ;
        RECT 1215.465 1089.785 1215.635 1089.955 ;
        RECT 1215.465 855.185 1215.635 855.355 ;
        RECT 1215.465 669.205 1215.635 669.375 ;
        RECT 1215.925 530.825 1216.095 530.995 ;
        RECT 1215.005 324.105 1215.175 324.275 ;
        RECT 1215.005 227.545 1215.175 227.715 ;
      LAYER met1 ;
        RECT 1214.945 1538.740 1215.235 1538.785 ;
        RECT 1215.390 1538.740 1215.710 1538.800 ;
        RECT 1214.945 1538.600 1215.710 1538.740 ;
        RECT 1214.945 1538.555 1215.235 1538.600 ;
        RECT 1215.390 1538.540 1215.710 1538.600 ;
        RECT 1214.930 1490.800 1215.250 1490.860 ;
        RECT 1214.735 1490.660 1215.250 1490.800 ;
        RECT 1214.930 1490.600 1215.250 1490.660 ;
        RECT 1214.930 1414.300 1215.250 1414.360 ;
        RECT 1215.850 1414.300 1216.170 1414.360 ;
        RECT 1214.930 1414.160 1216.170 1414.300 ;
        RECT 1214.930 1414.100 1215.250 1414.160 ;
        RECT 1215.850 1414.100 1216.170 1414.160 ;
        RECT 1214.010 1400.700 1214.330 1400.760 ;
        RECT 1215.850 1400.700 1216.170 1400.760 ;
        RECT 1214.010 1400.560 1216.170 1400.700 ;
        RECT 1214.010 1400.500 1214.330 1400.560 ;
        RECT 1215.850 1400.500 1216.170 1400.560 ;
        RECT 1215.850 1317.880 1216.170 1318.140 ;
        RECT 1215.940 1317.460 1216.080 1317.880 ;
        RECT 1215.850 1317.200 1216.170 1317.460 ;
        RECT 1214.010 1304.140 1214.330 1304.200 ;
        RECT 1215.850 1304.140 1216.170 1304.200 ;
        RECT 1214.010 1304.000 1216.170 1304.140 ;
        RECT 1214.010 1303.940 1214.330 1304.000 ;
        RECT 1215.850 1303.940 1216.170 1304.000 ;
        RECT 1214.930 1207.580 1215.250 1207.640 ;
        RECT 1215.850 1207.580 1216.170 1207.640 ;
        RECT 1214.930 1207.440 1216.170 1207.580 ;
        RECT 1214.930 1207.380 1215.250 1207.440 ;
        RECT 1215.850 1207.380 1216.170 1207.440 ;
        RECT 1214.930 1159.300 1215.250 1159.360 ;
        RECT 1215.390 1159.300 1215.710 1159.360 ;
        RECT 1214.930 1159.160 1215.710 1159.300 ;
        RECT 1214.930 1159.100 1215.250 1159.160 ;
        RECT 1215.390 1159.100 1215.710 1159.160 ;
        RECT 1215.850 1158.620 1216.170 1158.680 ;
        RECT 1215.655 1158.480 1216.170 1158.620 ;
        RECT 1215.850 1158.420 1216.170 1158.480 ;
        RECT 1215.865 1121.220 1216.155 1121.265 ;
        RECT 1216.770 1121.220 1217.090 1121.280 ;
        RECT 1215.865 1121.080 1217.090 1121.220 ;
        RECT 1215.865 1121.035 1216.155 1121.080 ;
        RECT 1216.770 1121.020 1217.090 1121.080 ;
        RECT 1215.390 1097.080 1215.710 1097.140 ;
        RECT 1216.770 1097.080 1217.090 1097.140 ;
        RECT 1215.390 1096.940 1217.090 1097.080 ;
        RECT 1215.390 1096.880 1215.710 1096.940 ;
        RECT 1216.770 1096.880 1217.090 1096.940 ;
        RECT 1215.390 1089.940 1215.710 1090.000 ;
        RECT 1215.195 1089.800 1215.710 1089.940 ;
        RECT 1215.390 1089.740 1215.710 1089.800 ;
        RECT 1215.390 1007.320 1215.710 1007.380 ;
        RECT 1215.195 1007.180 1215.710 1007.320 ;
        RECT 1215.390 1007.120 1215.710 1007.180 ;
        RECT 1215.850 980.260 1216.170 980.520 ;
        RECT 1215.940 979.840 1216.080 980.260 ;
        RECT 1215.850 979.580 1216.170 979.840 ;
        RECT 1215.850 903.960 1216.170 904.020 ;
        RECT 1216.770 903.960 1217.090 904.020 ;
        RECT 1215.850 903.820 1217.090 903.960 ;
        RECT 1215.850 903.760 1216.170 903.820 ;
        RECT 1216.770 903.760 1217.090 903.820 ;
        RECT 1215.390 855.340 1215.710 855.400 ;
        RECT 1215.195 855.200 1215.710 855.340 ;
        RECT 1215.390 855.140 1215.710 855.200 ;
        RECT 1215.405 807.400 1215.695 807.445 ;
        RECT 1215.850 807.400 1216.170 807.460 ;
        RECT 1215.405 807.260 1216.170 807.400 ;
        RECT 1215.405 807.215 1215.695 807.260 ;
        RECT 1215.850 807.200 1216.170 807.260 ;
        RECT 1215.850 787.140 1216.170 787.400 ;
        RECT 1215.940 786.720 1216.080 787.140 ;
        RECT 1215.850 786.460 1216.170 786.720 ;
        RECT 1215.390 669.360 1215.710 669.420 ;
        RECT 1215.195 669.220 1215.710 669.360 ;
        RECT 1215.390 669.160 1215.710 669.220 ;
        RECT 1215.405 621.080 1215.695 621.125 ;
        RECT 1216.310 621.080 1216.630 621.140 ;
        RECT 1215.405 620.940 1216.630 621.080 ;
        RECT 1215.405 620.895 1215.695 620.940 ;
        RECT 1216.310 620.880 1216.630 620.940 ;
        RECT 1215.390 545.060 1215.710 545.320 ;
        RECT 1215.480 544.920 1215.620 545.060 ;
        RECT 1215.850 544.920 1216.170 544.980 ;
        RECT 1215.480 544.780 1216.170 544.920 ;
        RECT 1215.850 544.720 1216.170 544.780 ;
        RECT 1215.850 530.980 1216.170 531.040 ;
        RECT 1215.655 530.840 1216.170 530.980 ;
        RECT 1215.850 530.780 1216.170 530.840 ;
        RECT 1215.850 483.720 1216.170 483.780 ;
        RECT 1215.655 483.580 1216.170 483.720 ;
        RECT 1215.850 483.520 1216.170 483.580 ;
        RECT 1215.390 483.040 1215.710 483.100 ;
        RECT 1215.850 483.040 1216.170 483.100 ;
        RECT 1215.390 482.900 1216.170 483.040 ;
        RECT 1215.390 482.840 1215.710 482.900 ;
        RECT 1215.850 482.840 1216.170 482.900 ;
        RECT 1215.390 434.420 1215.710 434.480 ;
        RECT 1216.310 434.420 1216.630 434.480 ;
        RECT 1215.390 434.280 1216.630 434.420 ;
        RECT 1215.390 434.220 1215.710 434.280 ;
        RECT 1216.310 434.220 1216.630 434.280 ;
        RECT 1215.390 351.940 1215.710 352.200 ;
        RECT 1215.480 351.460 1215.620 351.940 ;
        RECT 1215.850 351.460 1216.170 351.520 ;
        RECT 1215.480 351.320 1216.170 351.460 ;
        RECT 1215.850 351.260 1216.170 351.320 ;
        RECT 1214.945 324.260 1215.235 324.305 ;
        RECT 1215.850 324.260 1216.170 324.320 ;
        RECT 1214.945 324.120 1216.170 324.260 ;
        RECT 1214.945 324.075 1215.235 324.120 ;
        RECT 1215.850 324.060 1216.170 324.120 ;
        RECT 1214.930 276.320 1215.250 276.380 ;
        RECT 1214.735 276.180 1215.250 276.320 ;
        RECT 1214.930 276.120 1215.250 276.180 ;
        RECT 1215.850 234.500 1216.170 234.560 ;
        RECT 1216.310 234.500 1216.630 234.560 ;
        RECT 1215.850 234.360 1216.630 234.500 ;
        RECT 1215.850 234.300 1216.170 234.360 ;
        RECT 1216.310 234.300 1216.630 234.360 ;
        RECT 1214.945 227.700 1215.235 227.745 ;
        RECT 1216.310 227.700 1216.630 227.760 ;
        RECT 1214.945 227.560 1216.630 227.700 ;
        RECT 1214.945 227.515 1215.235 227.560 ;
        RECT 1216.310 227.500 1216.630 227.560 ;
        RECT 1214.930 179.760 1215.250 179.820 ;
        RECT 1214.735 179.620 1215.250 179.760 ;
        RECT 1214.930 179.560 1215.250 179.620 ;
        RECT 144.510 79.800 144.830 79.860 ;
        RECT 1215.390 79.800 1215.710 79.860 ;
        RECT 144.510 79.660 1215.710 79.800 ;
        RECT 144.510 79.600 144.830 79.660 ;
        RECT 1215.390 79.600 1215.710 79.660 ;
        RECT 139.450 15.880 139.770 15.940 ;
        RECT 144.510 15.880 144.830 15.940 ;
        RECT 139.450 15.740 144.830 15.880 ;
        RECT 139.450 15.680 139.770 15.740 ;
        RECT 144.510 15.680 144.830 15.740 ;
      LAYER via ;
        RECT 1215.420 1538.540 1215.680 1538.800 ;
        RECT 1214.960 1490.600 1215.220 1490.860 ;
        RECT 1214.960 1414.100 1215.220 1414.360 ;
        RECT 1215.880 1414.100 1216.140 1414.360 ;
        RECT 1214.040 1400.500 1214.300 1400.760 ;
        RECT 1215.880 1400.500 1216.140 1400.760 ;
        RECT 1215.880 1317.880 1216.140 1318.140 ;
        RECT 1215.880 1317.200 1216.140 1317.460 ;
        RECT 1214.040 1303.940 1214.300 1304.200 ;
        RECT 1215.880 1303.940 1216.140 1304.200 ;
        RECT 1214.960 1207.380 1215.220 1207.640 ;
        RECT 1215.880 1207.380 1216.140 1207.640 ;
        RECT 1214.960 1159.100 1215.220 1159.360 ;
        RECT 1215.420 1159.100 1215.680 1159.360 ;
        RECT 1215.880 1158.420 1216.140 1158.680 ;
        RECT 1216.800 1121.020 1217.060 1121.280 ;
        RECT 1215.420 1096.880 1215.680 1097.140 ;
        RECT 1216.800 1096.880 1217.060 1097.140 ;
        RECT 1215.420 1089.740 1215.680 1090.000 ;
        RECT 1215.420 1007.120 1215.680 1007.380 ;
        RECT 1215.880 980.260 1216.140 980.520 ;
        RECT 1215.880 979.580 1216.140 979.840 ;
        RECT 1215.880 903.760 1216.140 904.020 ;
        RECT 1216.800 903.760 1217.060 904.020 ;
        RECT 1215.420 855.140 1215.680 855.400 ;
        RECT 1215.880 807.200 1216.140 807.460 ;
        RECT 1215.880 787.140 1216.140 787.400 ;
        RECT 1215.880 786.460 1216.140 786.720 ;
        RECT 1215.420 669.160 1215.680 669.420 ;
        RECT 1216.340 620.880 1216.600 621.140 ;
        RECT 1215.420 545.060 1215.680 545.320 ;
        RECT 1215.880 544.720 1216.140 544.980 ;
        RECT 1215.880 530.780 1216.140 531.040 ;
        RECT 1215.880 483.520 1216.140 483.780 ;
        RECT 1215.420 482.840 1215.680 483.100 ;
        RECT 1215.880 482.840 1216.140 483.100 ;
        RECT 1215.420 434.220 1215.680 434.480 ;
        RECT 1216.340 434.220 1216.600 434.480 ;
        RECT 1215.420 351.940 1215.680 352.200 ;
        RECT 1215.880 351.260 1216.140 351.520 ;
        RECT 1215.880 324.060 1216.140 324.320 ;
        RECT 1214.960 276.120 1215.220 276.380 ;
        RECT 1215.880 234.300 1216.140 234.560 ;
        RECT 1216.340 234.300 1216.600 234.560 ;
        RECT 1216.340 227.500 1216.600 227.760 ;
        RECT 1214.960 179.560 1215.220 179.820 ;
        RECT 144.540 79.600 144.800 79.860 ;
        RECT 1215.420 79.600 1215.680 79.860 ;
        RECT 139.480 15.680 139.740 15.940 ;
        RECT 144.540 15.680 144.800 15.940 ;
      LAYER met2 ;
        RECT 1220.400 1701.090 1220.680 1702.400 ;
        RECT 1217.780 1700.950 1220.680 1701.090 ;
        RECT 1217.780 1636.605 1217.920 1700.950 ;
        RECT 1220.400 1700.000 1220.680 1700.950 ;
        RECT 1217.710 1636.235 1217.990 1636.605 ;
        RECT 1215.410 1635.555 1215.690 1635.925 ;
        RECT 1215.480 1538.830 1215.620 1635.555 ;
        RECT 1215.420 1538.510 1215.680 1538.830 ;
        RECT 1214.960 1490.570 1215.220 1490.890 ;
        RECT 1215.020 1414.390 1215.160 1490.570 ;
        RECT 1214.960 1414.070 1215.220 1414.390 ;
        RECT 1215.880 1414.070 1216.140 1414.390 ;
        RECT 1215.940 1400.790 1216.080 1414.070 ;
        RECT 1214.040 1400.470 1214.300 1400.790 ;
        RECT 1215.880 1400.470 1216.140 1400.790 ;
        RECT 1214.100 1353.045 1214.240 1400.470 ;
        RECT 1214.030 1352.675 1214.310 1353.045 ;
        RECT 1215.870 1351.995 1216.150 1352.365 ;
        RECT 1215.940 1318.170 1216.080 1351.995 ;
        RECT 1215.880 1317.850 1216.140 1318.170 ;
        RECT 1215.880 1317.170 1216.140 1317.490 ;
        RECT 1215.940 1304.230 1216.080 1317.170 ;
        RECT 1214.040 1303.910 1214.300 1304.230 ;
        RECT 1215.880 1303.910 1216.140 1304.230 ;
        RECT 1214.100 1256.485 1214.240 1303.910 ;
        RECT 1214.030 1256.115 1214.310 1256.485 ;
        RECT 1214.950 1255.435 1215.230 1255.805 ;
        RECT 1215.020 1207.670 1215.160 1255.435 ;
        RECT 1214.960 1207.525 1215.220 1207.670 ;
        RECT 1215.880 1207.525 1216.140 1207.670 ;
        RECT 1214.950 1207.155 1215.230 1207.525 ;
        RECT 1215.870 1207.155 1216.150 1207.525 ;
        RECT 1215.020 1159.390 1215.160 1207.155 ;
        RECT 1214.960 1159.070 1215.220 1159.390 ;
        RECT 1215.420 1159.130 1215.680 1159.390 ;
        RECT 1215.420 1159.070 1216.080 1159.130 ;
        RECT 1215.480 1158.990 1216.080 1159.070 ;
        RECT 1215.940 1158.710 1216.080 1158.990 ;
        RECT 1215.880 1158.390 1216.140 1158.710 ;
        RECT 1216.800 1120.990 1217.060 1121.310 ;
        RECT 1216.860 1097.170 1217.000 1120.990 ;
        RECT 1215.420 1096.850 1215.680 1097.170 ;
        RECT 1216.800 1096.850 1217.060 1097.170 ;
        RECT 1215.480 1090.030 1215.620 1096.850 ;
        RECT 1215.420 1089.710 1215.680 1090.030 ;
        RECT 1215.420 1007.090 1215.680 1007.410 ;
        RECT 1215.480 1000.690 1215.620 1007.090 ;
        RECT 1215.480 1000.550 1216.080 1000.690 ;
        RECT 1215.940 980.550 1216.080 1000.550 ;
        RECT 1215.880 980.230 1216.140 980.550 ;
        RECT 1215.880 979.550 1216.140 979.870 ;
        RECT 1215.940 904.050 1216.080 979.550 ;
        RECT 1215.880 903.730 1216.140 904.050 ;
        RECT 1216.800 903.730 1217.060 904.050 ;
        RECT 1216.860 855.965 1217.000 903.730 ;
        RECT 1215.870 855.850 1216.150 855.965 ;
        RECT 1215.480 855.710 1216.150 855.850 ;
        RECT 1215.480 855.430 1215.620 855.710 ;
        RECT 1215.870 855.595 1216.150 855.710 ;
        RECT 1216.790 855.595 1217.070 855.965 ;
        RECT 1215.420 855.110 1215.680 855.430 ;
        RECT 1215.880 807.170 1216.140 807.490 ;
        RECT 1215.940 787.430 1216.080 807.170 ;
        RECT 1215.880 787.110 1216.140 787.430 ;
        RECT 1215.880 786.430 1216.140 786.750 ;
        RECT 1215.940 676.330 1216.080 786.430 ;
        RECT 1215.480 676.190 1216.080 676.330 ;
        RECT 1215.480 669.450 1215.620 676.190 ;
        RECT 1215.420 669.130 1215.680 669.450 ;
        RECT 1216.340 620.850 1216.600 621.170 ;
        RECT 1216.400 596.090 1216.540 620.850 ;
        RECT 1215.480 595.950 1216.540 596.090 ;
        RECT 1215.480 545.350 1215.620 595.950 ;
        RECT 1215.420 545.030 1215.680 545.350 ;
        RECT 1215.880 544.690 1216.140 545.010 ;
        RECT 1215.940 531.070 1216.080 544.690 ;
        RECT 1215.880 530.750 1216.140 531.070 ;
        RECT 1215.880 483.490 1216.140 483.810 ;
        RECT 1215.940 483.130 1216.080 483.490 ;
        RECT 1215.420 482.810 1215.680 483.130 ;
        RECT 1215.880 482.810 1216.140 483.130 ;
        RECT 1215.480 434.510 1215.620 482.810 ;
        RECT 1215.420 434.190 1215.680 434.510 ;
        RECT 1216.340 434.190 1216.600 434.510 ;
        RECT 1216.400 387.445 1216.540 434.190 ;
        RECT 1216.330 387.075 1216.610 387.445 ;
        RECT 1215.410 379.595 1215.690 379.965 ;
        RECT 1215.480 352.230 1215.620 379.595 ;
        RECT 1215.420 351.910 1215.680 352.230 ;
        RECT 1215.880 351.230 1216.140 351.550 ;
        RECT 1215.940 324.350 1216.080 351.230 ;
        RECT 1215.880 324.030 1216.140 324.350 ;
        RECT 1214.960 276.090 1215.220 276.410 ;
        RECT 1215.020 254.730 1215.160 276.090 ;
        RECT 1215.020 254.590 1216.080 254.730 ;
        RECT 1215.940 234.590 1216.080 254.590 ;
        RECT 1215.880 234.270 1216.140 234.590 ;
        RECT 1216.340 234.270 1216.600 234.590 ;
        RECT 1216.400 227.790 1216.540 234.270 ;
        RECT 1216.340 227.470 1216.600 227.790 ;
        RECT 1214.960 179.530 1215.220 179.850 ;
        RECT 1215.020 158.170 1215.160 179.530 ;
        RECT 1215.020 158.030 1215.620 158.170 ;
        RECT 1215.480 79.890 1215.620 158.030 ;
        RECT 144.540 79.570 144.800 79.890 ;
        RECT 1215.420 79.570 1215.680 79.890 ;
        RECT 144.600 15.970 144.740 79.570 ;
        RECT 139.480 15.650 139.740 15.970 ;
        RECT 144.540 15.650 144.800 15.970 ;
        RECT 139.540 2.400 139.680 15.650 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 1217.710 1636.280 1217.990 1636.560 ;
        RECT 1215.410 1635.600 1215.690 1635.880 ;
        RECT 1214.030 1352.720 1214.310 1353.000 ;
        RECT 1215.870 1352.040 1216.150 1352.320 ;
        RECT 1214.030 1256.160 1214.310 1256.440 ;
        RECT 1214.950 1255.480 1215.230 1255.760 ;
        RECT 1214.950 1207.200 1215.230 1207.480 ;
        RECT 1215.870 1207.200 1216.150 1207.480 ;
        RECT 1215.870 855.640 1216.150 855.920 ;
        RECT 1216.790 855.640 1217.070 855.920 ;
        RECT 1216.330 387.120 1216.610 387.400 ;
        RECT 1215.410 379.640 1215.690 379.920 ;
      LAYER met3 ;
        RECT 1217.685 1636.570 1218.015 1636.585 ;
        RECT 1214.710 1636.270 1218.015 1636.570 ;
        RECT 1214.710 1635.890 1215.010 1636.270 ;
        RECT 1217.685 1636.255 1218.015 1636.270 ;
        RECT 1215.385 1635.890 1215.715 1635.905 ;
        RECT 1214.710 1635.590 1215.715 1635.890 ;
        RECT 1215.385 1635.575 1215.715 1635.590 ;
        RECT 1214.005 1353.010 1214.335 1353.025 ;
        RECT 1214.005 1352.710 1215.010 1353.010 ;
        RECT 1214.005 1352.695 1214.335 1352.710 ;
        RECT 1214.710 1352.330 1215.010 1352.710 ;
        RECT 1215.845 1352.330 1216.175 1352.345 ;
        RECT 1214.710 1352.030 1216.175 1352.330 ;
        RECT 1215.845 1352.015 1216.175 1352.030 ;
        RECT 1214.005 1256.450 1214.335 1256.465 ;
        RECT 1214.005 1256.150 1215.010 1256.450 ;
        RECT 1214.005 1256.135 1214.335 1256.150 ;
        RECT 1214.710 1255.785 1215.010 1256.150 ;
        RECT 1214.710 1255.470 1215.255 1255.785 ;
        RECT 1214.925 1255.455 1215.255 1255.470 ;
        RECT 1214.925 1207.490 1215.255 1207.505 ;
        RECT 1215.845 1207.490 1216.175 1207.505 ;
        RECT 1214.925 1207.190 1216.175 1207.490 ;
        RECT 1214.925 1207.175 1215.255 1207.190 ;
        RECT 1215.845 1207.175 1216.175 1207.190 ;
        RECT 1215.845 855.930 1216.175 855.945 ;
        RECT 1216.765 855.930 1217.095 855.945 ;
        RECT 1215.845 855.630 1217.095 855.930 ;
        RECT 1215.845 855.615 1216.175 855.630 ;
        RECT 1216.765 855.615 1217.095 855.630 ;
        RECT 1215.590 387.410 1215.970 387.420 ;
        RECT 1216.305 387.410 1216.635 387.425 ;
        RECT 1215.590 387.110 1216.635 387.410 ;
        RECT 1215.590 387.100 1215.970 387.110 ;
        RECT 1216.305 387.095 1216.635 387.110 ;
        RECT 1215.385 379.940 1215.715 379.945 ;
        RECT 1215.385 379.930 1215.970 379.940 ;
        RECT 1215.385 379.630 1216.170 379.930 ;
        RECT 1215.385 379.620 1215.970 379.630 ;
        RECT 1215.385 379.615 1215.715 379.620 ;
      LAYER via3 ;
        RECT 1215.620 387.100 1215.940 387.420 ;
        RECT 1215.620 379.620 1215.940 379.940 ;
      LAYER met4 ;
        RECT 1215.615 387.095 1215.945 387.425 ;
        RECT 1215.630 379.945 1215.930 387.095 ;
        RECT 1215.615 379.615 1215.945 379.945 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 79.460 158.630 79.520 ;
        RECT 1228.730 79.460 1229.050 79.520 ;
        RECT 158.310 79.320 1229.050 79.460 ;
        RECT 158.310 79.260 158.630 79.320 ;
        RECT 1228.730 79.260 1229.050 79.320 ;
      LAYER via ;
        RECT 158.340 79.260 158.600 79.520 ;
        RECT 1228.760 79.260 1229.020 79.520 ;
      LAYER met2 ;
        RECT 1229.600 1700.410 1229.880 1702.400 ;
        RECT 1228.820 1700.270 1229.880 1700.410 ;
        RECT 1228.820 79.550 1228.960 1700.270 ;
        RECT 1229.600 1700.000 1229.880 1700.270 ;
        RECT 158.340 79.230 158.600 79.550 ;
        RECT 1228.760 79.230 1229.020 79.550 ;
        RECT 158.400 3.130 158.540 79.230 ;
        RECT 157.480 2.990 158.540 3.130 ;
        RECT 157.480 2.400 157.620 2.990 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 230.990 1689.020 231.310 1689.080 ;
        RECT 1238.390 1689.020 1238.710 1689.080 ;
        RECT 230.990 1688.880 1238.710 1689.020 ;
        RECT 230.990 1688.820 231.310 1688.880 ;
        RECT 1238.390 1688.820 1238.710 1688.880 ;
        RECT 174.870 19.960 175.190 20.020 ;
        RECT 230.990 19.960 231.310 20.020 ;
        RECT 174.870 19.820 231.310 19.960 ;
        RECT 174.870 19.760 175.190 19.820 ;
        RECT 230.990 19.760 231.310 19.820 ;
      LAYER via ;
        RECT 231.020 1688.820 231.280 1689.080 ;
        RECT 1238.420 1688.820 1238.680 1689.080 ;
        RECT 174.900 19.760 175.160 20.020 ;
        RECT 231.020 19.760 231.280 20.020 ;
      LAYER met2 ;
        RECT 1238.340 1700.000 1238.620 1702.400 ;
        RECT 1238.480 1689.110 1238.620 1700.000 ;
        RECT 231.020 1688.790 231.280 1689.110 ;
        RECT 1238.420 1688.790 1238.680 1689.110 ;
        RECT 231.080 20.050 231.220 1688.790 ;
        RECT 174.900 19.730 175.160 20.050 ;
        RECT 231.020 19.730 231.280 20.050 ;
        RECT 174.960 2.400 175.100 19.730 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.070 1688.680 1242.390 1688.740 ;
        RECT 1247.590 1688.680 1247.910 1688.740 ;
        RECT 1242.070 1688.540 1247.910 1688.680 ;
        RECT 1242.070 1688.480 1242.390 1688.540 ;
        RECT 1247.590 1688.480 1247.910 1688.540 ;
        RECT 192.810 18.940 193.130 19.000 ;
        RECT 1242.070 18.940 1242.390 19.000 ;
        RECT 192.810 18.800 1242.390 18.940 ;
        RECT 192.810 18.740 193.130 18.800 ;
        RECT 1242.070 18.740 1242.390 18.800 ;
      LAYER via ;
        RECT 1242.100 1688.480 1242.360 1688.740 ;
        RECT 1247.620 1688.480 1247.880 1688.740 ;
        RECT 192.840 18.740 193.100 19.000 ;
        RECT 1242.100 18.740 1242.360 19.000 ;
      LAYER met2 ;
        RECT 1247.540 1700.000 1247.820 1702.400 ;
        RECT 1247.680 1688.770 1247.820 1700.000 ;
        RECT 1242.100 1688.450 1242.360 1688.770 ;
        RECT 1247.620 1688.450 1247.880 1688.770 ;
        RECT 1242.160 19.030 1242.300 1688.450 ;
        RECT 192.840 18.710 193.100 19.030 ;
        RECT 1242.100 18.710 1242.360 19.030 ;
        RECT 192.900 2.400 193.040 18.710 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 251.690 1689.360 252.010 1689.420 ;
        RECT 1256.790 1689.360 1257.110 1689.420 ;
        RECT 251.690 1689.220 1257.110 1689.360 ;
        RECT 251.690 1689.160 252.010 1689.220 ;
        RECT 1256.790 1689.160 1257.110 1689.220 ;
        RECT 210.750 20.640 211.070 20.700 ;
        RECT 251.690 20.640 252.010 20.700 ;
        RECT 210.750 20.500 252.010 20.640 ;
        RECT 210.750 20.440 211.070 20.500 ;
        RECT 251.690 20.440 252.010 20.500 ;
      LAYER via ;
        RECT 251.720 1689.160 251.980 1689.420 ;
        RECT 1256.820 1689.160 1257.080 1689.420 ;
        RECT 210.780 20.440 211.040 20.700 ;
        RECT 251.720 20.440 251.980 20.700 ;
      LAYER met2 ;
        RECT 1256.740 1700.000 1257.020 1702.400 ;
        RECT 1256.880 1689.450 1257.020 1700.000 ;
        RECT 251.720 1689.130 251.980 1689.450 ;
        RECT 1256.820 1689.130 1257.080 1689.450 ;
        RECT 251.780 20.730 251.920 1689.130 ;
        RECT 210.780 20.410 211.040 20.730 ;
        RECT 251.720 20.410 251.980 20.730 ;
        RECT 210.840 2.400 210.980 20.410 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1259.090 1672.020 1259.410 1672.080 ;
        RECT 1265.990 1672.020 1266.310 1672.080 ;
        RECT 1259.090 1671.880 1266.310 1672.020 ;
        RECT 1259.090 1671.820 1259.410 1671.880 ;
        RECT 1265.990 1671.820 1266.310 1671.880 ;
        RECT 228.690 19.620 229.010 19.680 ;
        RECT 1259.090 19.620 1259.410 19.680 ;
        RECT 228.690 19.480 1259.410 19.620 ;
        RECT 228.690 19.420 229.010 19.480 ;
        RECT 1259.090 19.420 1259.410 19.480 ;
      LAYER via ;
        RECT 1259.120 1671.820 1259.380 1672.080 ;
        RECT 1266.020 1671.820 1266.280 1672.080 ;
        RECT 228.720 19.420 228.980 19.680 ;
        RECT 1259.120 19.420 1259.380 19.680 ;
      LAYER met2 ;
        RECT 1265.940 1700.000 1266.220 1702.400 ;
        RECT 1266.080 1672.110 1266.220 1700.000 ;
        RECT 1259.120 1671.790 1259.380 1672.110 ;
        RECT 1266.020 1671.790 1266.280 1672.110 ;
        RECT 1259.180 19.710 1259.320 1671.790 ;
        RECT 228.720 19.390 228.980 19.710 ;
        RECT 1259.120 19.390 1259.380 19.710 ;
        RECT 228.780 2.400 228.920 19.390 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1140.870 1687.660 1141.190 1687.720 ;
        RECT 1174.450 1687.660 1174.770 1687.720 ;
        RECT 1140.870 1687.520 1174.770 1687.660 ;
        RECT 1140.870 1687.460 1141.190 1687.520 ;
        RECT 1174.450 1687.460 1174.770 1687.520 ;
        RECT 79.190 1686.980 79.510 1687.040 ;
        RECT 1140.870 1686.980 1141.190 1687.040 ;
        RECT 79.190 1686.840 1141.190 1686.980 ;
        RECT 79.190 1686.780 79.510 1686.840 ;
        RECT 1140.870 1686.780 1141.190 1686.840 ;
        RECT 50.210 15.200 50.530 15.260 ;
        RECT 79.190 15.200 79.510 15.260 ;
        RECT 50.210 15.060 79.510 15.200 ;
        RECT 50.210 15.000 50.530 15.060 ;
        RECT 79.190 15.000 79.510 15.060 ;
      LAYER via ;
        RECT 1140.900 1687.460 1141.160 1687.720 ;
        RECT 1174.480 1687.460 1174.740 1687.720 ;
        RECT 79.220 1686.780 79.480 1687.040 ;
        RECT 1140.900 1686.780 1141.160 1687.040 ;
        RECT 50.240 15.000 50.500 15.260 ;
        RECT 79.220 15.000 79.480 15.260 ;
      LAYER met2 ;
        RECT 1174.400 1700.000 1174.680 1702.400 ;
        RECT 1174.540 1687.750 1174.680 1700.000 ;
        RECT 1140.900 1687.430 1141.160 1687.750 ;
        RECT 1174.480 1687.430 1174.740 1687.750 ;
        RECT 1140.960 1687.070 1141.100 1687.430 ;
        RECT 79.220 1686.750 79.480 1687.070 ;
        RECT 1140.900 1686.750 1141.160 1687.070 ;
        RECT 79.280 15.290 79.420 1686.750 ;
        RECT 50.240 14.970 50.500 15.290 ;
        RECT 79.220 14.970 79.480 15.290 ;
        RECT 50.300 2.400 50.440 14.970 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1265.990 1671.340 1266.310 1671.400 ;
        RECT 1278.410 1671.340 1278.730 1671.400 ;
        RECT 1265.990 1671.200 1278.730 1671.340 ;
        RECT 1265.990 1671.140 1266.310 1671.200 ;
        RECT 1278.410 1671.140 1278.730 1671.200 ;
        RECT 252.610 20.300 252.930 20.360 ;
        RECT 1265.990 20.300 1266.310 20.360 ;
        RECT 252.610 20.160 1266.310 20.300 ;
        RECT 252.610 20.100 252.930 20.160 ;
        RECT 1265.990 20.100 1266.310 20.160 ;
      LAYER via ;
        RECT 1266.020 1671.140 1266.280 1671.400 ;
        RECT 1278.440 1671.140 1278.700 1671.400 ;
        RECT 252.640 20.100 252.900 20.360 ;
        RECT 1266.020 20.100 1266.280 20.360 ;
      LAYER met2 ;
        RECT 1278.360 1700.000 1278.640 1702.400 ;
        RECT 1278.500 1671.430 1278.640 1700.000 ;
        RECT 1266.020 1671.110 1266.280 1671.430 ;
        RECT 1278.440 1671.110 1278.700 1671.430 ;
        RECT 1266.080 20.390 1266.220 1671.110 ;
        RECT 252.640 20.070 252.900 20.390 ;
        RECT 1266.020 20.070 1266.280 20.390 ;
        RECT 252.700 2.400 252.840 20.070 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 286.190 1689.700 286.510 1689.760 ;
        RECT 1287.610 1689.700 1287.930 1689.760 ;
        RECT 286.190 1689.560 1287.930 1689.700 ;
        RECT 286.190 1689.500 286.510 1689.560 ;
        RECT 1287.610 1689.500 1287.930 1689.560 ;
        RECT 270.090 16.560 270.410 16.620 ;
        RECT 286.190 16.560 286.510 16.620 ;
        RECT 270.090 16.420 286.510 16.560 ;
        RECT 270.090 16.360 270.410 16.420 ;
        RECT 286.190 16.360 286.510 16.420 ;
      LAYER via ;
        RECT 286.220 1689.500 286.480 1689.760 ;
        RECT 1287.640 1689.500 1287.900 1689.760 ;
        RECT 270.120 16.360 270.380 16.620 ;
        RECT 286.220 16.360 286.480 16.620 ;
      LAYER met2 ;
        RECT 1287.560 1700.000 1287.840 1702.400 ;
        RECT 1287.700 1689.790 1287.840 1700.000 ;
        RECT 286.220 1689.470 286.480 1689.790 ;
        RECT 1287.640 1689.470 1287.900 1689.790 ;
        RECT 286.280 16.650 286.420 1689.470 ;
        RECT 270.120 16.330 270.380 16.650 ;
        RECT 286.220 16.330 286.480 16.650 ;
        RECT 270.180 2.400 270.320 16.330 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1279.790 1686.640 1280.110 1686.700 ;
        RECT 1296.810 1686.640 1297.130 1686.700 ;
        RECT 1279.790 1686.500 1297.130 1686.640 ;
        RECT 1279.790 1686.440 1280.110 1686.500 ;
        RECT 1296.810 1686.440 1297.130 1686.500 ;
        RECT 288.030 20.640 288.350 20.700 ;
        RECT 1279.790 20.640 1280.110 20.700 ;
        RECT 288.030 20.500 1280.110 20.640 ;
        RECT 288.030 20.440 288.350 20.500 ;
        RECT 1279.790 20.440 1280.110 20.500 ;
      LAYER via ;
        RECT 1279.820 1686.440 1280.080 1686.700 ;
        RECT 1296.840 1686.440 1297.100 1686.700 ;
        RECT 288.060 20.440 288.320 20.700 ;
        RECT 1279.820 20.440 1280.080 20.700 ;
      LAYER met2 ;
        RECT 1296.760 1700.000 1297.040 1702.400 ;
        RECT 1296.900 1686.730 1297.040 1700.000 ;
        RECT 1279.820 1686.410 1280.080 1686.730 ;
        RECT 1296.840 1686.410 1297.100 1686.730 ;
        RECT 1279.880 20.730 1280.020 1686.410 ;
        RECT 288.060 20.410 288.320 20.730 ;
        RECT 1279.820 20.410 1280.080 20.730 ;
        RECT 288.120 2.400 288.260 20.410 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 334.490 1690.040 334.810 1690.100 ;
        RECT 1306.010 1690.040 1306.330 1690.100 ;
        RECT 334.490 1689.900 1306.330 1690.040 ;
        RECT 334.490 1689.840 334.810 1689.900 ;
        RECT 1306.010 1689.840 1306.330 1689.900 ;
        RECT 305.970 15.880 306.290 15.940 ;
        RECT 334.490 15.880 334.810 15.940 ;
        RECT 305.970 15.740 334.810 15.880 ;
        RECT 305.970 15.680 306.290 15.740 ;
        RECT 334.490 15.680 334.810 15.740 ;
      LAYER via ;
        RECT 334.520 1689.840 334.780 1690.100 ;
        RECT 1306.040 1689.840 1306.300 1690.100 ;
        RECT 306.000 15.680 306.260 15.940 ;
        RECT 334.520 15.680 334.780 15.940 ;
      LAYER met2 ;
        RECT 1305.960 1700.000 1306.240 1702.400 ;
        RECT 1306.100 1690.130 1306.240 1700.000 ;
        RECT 334.520 1689.810 334.780 1690.130 ;
        RECT 1306.040 1689.810 1306.300 1690.130 ;
        RECT 334.580 15.970 334.720 1689.810 ;
        RECT 306.000 15.650 306.260 15.970 ;
        RECT 334.520 15.650 334.780 15.970 ;
        RECT 306.060 2.400 306.200 15.650 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1286.690 1686.980 1287.010 1687.040 ;
        RECT 1315.210 1686.980 1315.530 1687.040 ;
        RECT 1286.690 1686.840 1315.530 1686.980 ;
        RECT 1286.690 1686.780 1287.010 1686.840 ;
        RECT 1315.210 1686.780 1315.530 1686.840 ;
        RECT 1286.690 16.900 1287.010 16.960 ;
        RECT 358.960 16.760 1287.010 16.900 ;
        RECT 323.910 16.220 324.230 16.280 ;
        RECT 358.960 16.220 359.100 16.760 ;
        RECT 1286.690 16.700 1287.010 16.760 ;
        RECT 323.910 16.080 359.100 16.220 ;
        RECT 323.910 16.020 324.230 16.080 ;
      LAYER via ;
        RECT 1286.720 1686.780 1286.980 1687.040 ;
        RECT 1315.240 1686.780 1315.500 1687.040 ;
        RECT 323.940 16.020 324.200 16.280 ;
        RECT 1286.720 16.700 1286.980 16.960 ;
      LAYER met2 ;
        RECT 1315.160 1700.000 1315.440 1702.400 ;
        RECT 1315.300 1687.070 1315.440 1700.000 ;
        RECT 1286.720 1686.750 1286.980 1687.070 ;
        RECT 1315.240 1686.750 1315.500 1687.070 ;
        RECT 1286.780 16.990 1286.920 1686.750 ;
        RECT 1286.720 16.670 1286.980 16.990 ;
        RECT 323.940 15.990 324.200 16.310 ;
        RECT 324.000 2.400 324.140 15.990 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 355.190 1690.380 355.510 1690.440 ;
        RECT 1324.410 1690.380 1324.730 1690.440 ;
        RECT 355.190 1690.240 1324.730 1690.380 ;
        RECT 355.190 1690.180 355.510 1690.240 ;
        RECT 1324.410 1690.180 1324.730 1690.240 ;
        RECT 341.390 15.200 341.710 15.260 ;
        RECT 355.190 15.200 355.510 15.260 ;
        RECT 341.390 15.060 355.510 15.200 ;
        RECT 341.390 15.000 341.710 15.060 ;
        RECT 355.190 15.000 355.510 15.060 ;
      LAYER via ;
        RECT 355.220 1690.180 355.480 1690.440 ;
        RECT 1324.440 1690.180 1324.700 1690.440 ;
        RECT 341.420 15.000 341.680 15.260 ;
        RECT 355.220 15.000 355.480 15.260 ;
      LAYER met2 ;
        RECT 1324.360 1700.000 1324.640 1702.400 ;
        RECT 1324.500 1690.470 1324.640 1700.000 ;
        RECT 355.220 1690.150 355.480 1690.470 ;
        RECT 1324.440 1690.150 1324.700 1690.470 ;
        RECT 355.280 15.290 355.420 1690.150 ;
        RECT 341.420 14.970 341.680 15.290 ;
        RECT 355.220 14.970 355.480 15.290 ;
        RECT 341.480 2.400 341.620 14.970 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1293.590 1688.680 1293.910 1688.740 ;
        RECT 1333.610 1688.680 1333.930 1688.740 ;
        RECT 1293.590 1688.540 1333.930 1688.680 ;
        RECT 1293.590 1688.480 1293.910 1688.540 ;
        RECT 1333.610 1688.480 1333.930 1688.540 ;
        RECT 359.330 16.560 359.650 16.620 ;
        RECT 1293.590 16.560 1293.910 16.620 ;
        RECT 359.330 16.420 1293.910 16.560 ;
        RECT 359.330 16.360 359.650 16.420 ;
        RECT 1293.590 16.360 1293.910 16.420 ;
      LAYER via ;
        RECT 1293.620 1688.480 1293.880 1688.740 ;
        RECT 1333.640 1688.480 1333.900 1688.740 ;
        RECT 359.360 16.360 359.620 16.620 ;
        RECT 1293.620 16.360 1293.880 16.620 ;
      LAYER met2 ;
        RECT 1333.560 1700.000 1333.840 1702.400 ;
        RECT 1333.700 1688.770 1333.840 1700.000 ;
        RECT 1293.620 1688.450 1293.880 1688.770 ;
        RECT 1333.640 1688.450 1333.900 1688.770 ;
        RECT 1293.680 16.650 1293.820 1688.450 ;
        RECT 359.360 16.330 359.620 16.650 ;
        RECT 1293.620 16.330 1293.880 16.650 ;
        RECT 359.420 2.400 359.560 16.330 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 534.590 1683.920 534.910 1683.980 ;
        RECT 1342.810 1683.920 1343.130 1683.980 ;
        RECT 534.590 1683.780 1335.220 1683.920 ;
        RECT 534.590 1683.720 534.910 1683.780 ;
        RECT 1335.080 1683.580 1335.220 1683.780 ;
        RECT 1338.300 1683.780 1343.130 1683.920 ;
        RECT 1338.300 1683.580 1338.440 1683.780 ;
        RECT 1342.810 1683.720 1343.130 1683.780 ;
        RECT 1335.080 1683.440 1338.440 1683.580 ;
        RECT 534.590 14.860 534.910 14.920 ;
        RECT 502.020 14.720 534.910 14.860 ;
        RECT 377.270 14.520 377.590 14.580 ;
        RECT 502.020 14.520 502.160 14.720 ;
        RECT 534.590 14.660 534.910 14.720 ;
        RECT 377.270 14.380 502.160 14.520 ;
        RECT 377.270 14.320 377.590 14.380 ;
      LAYER via ;
        RECT 534.620 1683.720 534.880 1683.980 ;
        RECT 1342.840 1683.720 1343.100 1683.980 ;
        RECT 377.300 14.320 377.560 14.580 ;
        RECT 534.620 14.660 534.880 14.920 ;
      LAYER met2 ;
        RECT 1342.760 1700.000 1343.040 1702.400 ;
        RECT 1342.900 1684.010 1343.040 1700.000 ;
        RECT 534.620 1683.690 534.880 1684.010 ;
        RECT 1342.840 1683.690 1343.100 1684.010 ;
        RECT 534.680 14.950 534.820 1683.690 ;
        RECT 534.620 14.630 534.880 14.950 ;
        RECT 377.300 14.290 377.560 14.610 ;
        RECT 377.360 2.400 377.500 14.290 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 414.605 14.705 414.775 15.895 ;
      LAYER mcon ;
        RECT 414.605 15.725 414.775 15.895 ;
      LAYER met1 ;
        RECT 1307.390 1687.320 1307.710 1687.380 ;
        RECT 1307.390 1687.180 1320.960 1687.320 ;
        RECT 1307.390 1687.120 1307.710 1687.180 ;
        RECT 1320.820 1686.640 1320.960 1687.180 ;
        RECT 1352.010 1686.640 1352.330 1686.700 ;
        RECT 1320.820 1686.500 1352.330 1686.640 ;
        RECT 1352.010 1686.440 1352.330 1686.500 ;
        RECT 1307.390 16.220 1307.710 16.280 ;
        RECT 448.660 16.080 1307.710 16.220 ;
        RECT 414.545 15.880 414.835 15.925 ;
        RECT 448.660 15.880 448.800 16.080 ;
        RECT 1307.390 16.020 1307.710 16.080 ;
        RECT 414.545 15.740 448.800 15.880 ;
        RECT 414.545 15.695 414.835 15.740 ;
        RECT 395.210 14.860 395.530 14.920 ;
        RECT 414.545 14.860 414.835 14.905 ;
        RECT 395.210 14.720 414.835 14.860 ;
        RECT 395.210 14.660 395.530 14.720 ;
        RECT 414.545 14.675 414.835 14.720 ;
      LAYER via ;
        RECT 1307.420 1687.120 1307.680 1687.380 ;
        RECT 1352.040 1686.440 1352.300 1686.700 ;
        RECT 1307.420 16.020 1307.680 16.280 ;
        RECT 395.240 14.660 395.500 14.920 ;
      LAYER met2 ;
        RECT 1351.960 1700.000 1352.240 1702.400 ;
        RECT 1307.420 1687.090 1307.680 1687.410 ;
        RECT 1307.480 16.310 1307.620 1687.090 ;
        RECT 1352.100 1686.730 1352.240 1700.000 ;
        RECT 1352.040 1686.410 1352.300 1686.730 ;
        RECT 1307.420 15.990 1307.680 16.310 ;
        RECT 395.240 14.630 395.500 14.950 ;
        RECT 395.300 2.400 395.440 14.630 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 424.190 1686.300 424.510 1686.360 ;
        RECT 1361.210 1686.300 1361.530 1686.360 ;
        RECT 424.190 1686.160 1361.530 1686.300 ;
        RECT 424.190 1686.100 424.510 1686.160 ;
        RECT 1361.210 1686.100 1361.530 1686.160 ;
        RECT 424.190 16.220 424.510 16.280 ;
        RECT 414.160 16.080 424.510 16.220 ;
        RECT 413.150 15.880 413.470 15.940 ;
        RECT 414.160 15.880 414.300 16.080 ;
        RECT 424.190 16.020 424.510 16.080 ;
        RECT 413.150 15.740 414.300 15.880 ;
        RECT 413.150 15.680 413.470 15.740 ;
      LAYER via ;
        RECT 424.220 1686.100 424.480 1686.360 ;
        RECT 1361.240 1686.100 1361.500 1686.360 ;
        RECT 413.180 15.680 413.440 15.940 ;
        RECT 424.220 16.020 424.480 16.280 ;
      LAYER met2 ;
        RECT 1361.160 1700.000 1361.440 1702.400 ;
        RECT 1361.300 1686.390 1361.440 1700.000 ;
        RECT 424.220 1686.070 424.480 1686.390 ;
        RECT 1361.240 1686.070 1361.500 1686.390 ;
        RECT 424.280 16.310 424.420 1686.070 ;
        RECT 424.220 15.990 424.480 16.310 ;
        RECT 413.180 15.650 413.440 15.970 ;
        RECT 413.240 2.400 413.380 15.650 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1181.425 1448.485 1181.595 1490.475 ;
        RECT 1181.425 1200.965 1181.595 1221.535 ;
        RECT 1181.425 1152.685 1181.595 1200.455 ;
        RECT 1181.425 1014.305 1181.595 1028.075 ;
        RECT 1181.425 945.285 1181.595 993.395 ;
        RECT 1181.885 807.245 1182.055 896.835 ;
        RECT 1182.345 662.405 1182.515 710.515 ;
        RECT 1181.885 565.845 1182.055 613.955 ;
        RECT 1181.425 379.525 1181.595 427.635 ;
        RECT 1181.425 338.045 1181.595 351.815 ;
        RECT 1181.885 235.025 1182.055 331.075 ;
      LAYER mcon ;
        RECT 1181.425 1490.305 1181.595 1490.475 ;
        RECT 1181.425 1221.365 1181.595 1221.535 ;
        RECT 1181.425 1200.285 1181.595 1200.455 ;
        RECT 1181.425 1027.905 1181.595 1028.075 ;
        RECT 1181.425 993.225 1181.595 993.395 ;
        RECT 1181.885 896.665 1182.055 896.835 ;
        RECT 1182.345 710.345 1182.515 710.515 ;
        RECT 1181.885 613.785 1182.055 613.955 ;
        RECT 1181.425 427.465 1181.595 427.635 ;
        RECT 1181.425 351.645 1181.595 351.815 ;
        RECT 1181.885 330.905 1182.055 331.075 ;
      LAYER met1 ;
        RECT 1181.350 1635.640 1181.670 1635.700 ;
        RECT 1184.570 1635.640 1184.890 1635.700 ;
        RECT 1181.350 1635.500 1184.890 1635.640 ;
        RECT 1181.350 1635.440 1181.670 1635.500 ;
        RECT 1184.570 1635.440 1184.890 1635.500 ;
        RECT 1181.350 1545.540 1181.670 1545.600 ;
        RECT 1181.810 1545.540 1182.130 1545.600 ;
        RECT 1181.350 1545.400 1182.130 1545.540 ;
        RECT 1181.350 1545.340 1181.670 1545.400 ;
        RECT 1181.810 1545.340 1182.130 1545.400 ;
        RECT 1181.350 1490.460 1181.670 1490.520 ;
        RECT 1181.155 1490.320 1181.670 1490.460 ;
        RECT 1181.350 1490.260 1181.670 1490.320 ;
        RECT 1181.365 1448.640 1181.655 1448.685 ;
        RECT 1182.270 1448.640 1182.590 1448.700 ;
        RECT 1181.365 1448.500 1182.590 1448.640 ;
        RECT 1181.365 1448.455 1181.655 1448.500 ;
        RECT 1182.270 1448.440 1182.590 1448.500 ;
        RECT 1181.810 1393.900 1182.130 1393.960 ;
        RECT 1183.190 1393.900 1183.510 1393.960 ;
        RECT 1181.810 1393.760 1183.510 1393.900 ;
        RECT 1181.810 1393.700 1182.130 1393.760 ;
        RECT 1183.190 1393.700 1183.510 1393.760 ;
        RECT 1181.810 1352.760 1182.130 1352.820 ;
        RECT 1181.440 1352.620 1182.130 1352.760 ;
        RECT 1181.440 1352.480 1181.580 1352.620 ;
        RECT 1181.810 1352.560 1182.130 1352.620 ;
        RECT 1181.350 1352.220 1181.670 1352.480 ;
        RECT 1181.350 1318.080 1181.670 1318.140 ;
        RECT 1181.350 1317.940 1182.040 1318.080 ;
        RECT 1181.350 1317.880 1181.670 1317.940 ;
        RECT 1181.900 1317.800 1182.040 1317.940 ;
        RECT 1181.810 1317.540 1182.130 1317.800 ;
        RECT 1181.810 1269.460 1182.130 1269.520 ;
        RECT 1181.440 1269.320 1182.130 1269.460 ;
        RECT 1181.440 1268.840 1181.580 1269.320 ;
        RECT 1181.810 1269.260 1182.130 1269.320 ;
        RECT 1181.350 1268.580 1181.670 1268.840 ;
        RECT 1181.350 1221.520 1181.670 1221.580 ;
        RECT 1181.155 1221.380 1181.670 1221.520 ;
        RECT 1181.350 1221.320 1181.670 1221.380 ;
        RECT 1181.350 1201.120 1181.670 1201.180 ;
        RECT 1181.155 1200.980 1181.670 1201.120 ;
        RECT 1181.350 1200.920 1181.670 1200.980 ;
        RECT 1181.350 1200.440 1181.670 1200.500 ;
        RECT 1181.155 1200.300 1181.670 1200.440 ;
        RECT 1181.350 1200.240 1181.670 1200.300 ;
        RECT 1181.350 1152.840 1181.670 1152.900 ;
        RECT 1181.155 1152.700 1181.670 1152.840 ;
        RECT 1181.350 1152.640 1181.670 1152.700 ;
        RECT 1181.350 1104.220 1181.670 1104.280 ;
        RECT 1182.270 1104.220 1182.590 1104.280 ;
        RECT 1181.350 1104.080 1182.590 1104.220 ;
        RECT 1181.350 1104.020 1181.670 1104.080 ;
        RECT 1182.270 1104.020 1182.590 1104.080 ;
        RECT 1181.810 1080.080 1182.130 1080.140 ;
        RECT 1182.730 1080.080 1183.050 1080.140 ;
        RECT 1181.810 1079.940 1183.050 1080.080 ;
        RECT 1181.810 1079.880 1182.130 1079.940 ;
        RECT 1182.730 1079.880 1183.050 1079.940 ;
        RECT 1181.350 1028.060 1181.670 1028.120 ;
        RECT 1181.155 1027.920 1181.670 1028.060 ;
        RECT 1181.350 1027.860 1181.670 1027.920 ;
        RECT 1181.350 1014.460 1181.670 1014.520 ;
        RECT 1181.155 1014.320 1181.670 1014.460 ;
        RECT 1181.350 1014.260 1181.670 1014.320 ;
        RECT 1181.350 993.380 1181.670 993.440 ;
        RECT 1181.155 993.240 1181.670 993.380 ;
        RECT 1181.350 993.180 1181.670 993.240 ;
        RECT 1181.365 945.440 1181.655 945.485 ;
        RECT 1181.810 945.440 1182.130 945.500 ;
        RECT 1181.365 945.300 1182.130 945.440 ;
        RECT 1181.365 945.255 1181.655 945.300 ;
        RECT 1181.810 945.240 1182.130 945.300 ;
        RECT 1181.810 896.820 1182.130 896.880 ;
        RECT 1181.615 896.680 1182.130 896.820 ;
        RECT 1181.810 896.620 1182.130 896.680 ;
        RECT 1181.810 807.400 1182.130 807.460 ;
        RECT 1181.615 807.260 1182.130 807.400 ;
        RECT 1181.810 807.200 1182.130 807.260 ;
        RECT 1181.350 765.920 1181.670 765.980 ;
        RECT 1181.810 765.920 1182.130 765.980 ;
        RECT 1181.350 765.780 1182.130 765.920 ;
        RECT 1181.350 765.720 1181.670 765.780 ;
        RECT 1181.810 765.720 1182.130 765.780 ;
        RECT 1181.350 717.640 1181.670 717.700 ;
        RECT 1182.270 717.640 1182.590 717.700 ;
        RECT 1181.350 717.500 1182.590 717.640 ;
        RECT 1181.350 717.440 1181.670 717.500 ;
        RECT 1182.270 717.440 1182.590 717.500 ;
        RECT 1182.270 710.500 1182.590 710.560 ;
        RECT 1182.075 710.360 1182.590 710.500 ;
        RECT 1182.270 710.300 1182.590 710.360 ;
        RECT 1182.270 662.560 1182.590 662.620 ;
        RECT 1182.075 662.420 1182.590 662.560 ;
        RECT 1182.270 662.360 1182.590 662.420 ;
        RECT 1181.810 621.420 1182.130 621.480 ;
        RECT 1182.270 621.420 1182.590 621.480 ;
        RECT 1181.810 621.280 1182.590 621.420 ;
        RECT 1181.810 621.220 1182.130 621.280 ;
        RECT 1182.270 621.220 1182.590 621.280 ;
        RECT 1181.810 613.940 1182.130 614.000 ;
        RECT 1181.615 613.800 1182.130 613.940 ;
        RECT 1181.810 613.740 1182.130 613.800 ;
        RECT 1181.825 566.000 1182.115 566.045 ;
        RECT 1182.270 566.000 1182.590 566.060 ;
        RECT 1181.825 565.860 1182.590 566.000 ;
        RECT 1181.825 565.815 1182.115 565.860 ;
        RECT 1182.270 565.800 1182.590 565.860 ;
        RECT 1181.350 530.980 1181.670 531.040 ;
        RECT 1182.730 530.980 1183.050 531.040 ;
        RECT 1181.350 530.840 1183.050 530.980 ;
        RECT 1181.350 530.780 1181.670 530.840 ;
        RECT 1182.730 530.780 1183.050 530.840 ;
        RECT 1181.350 427.620 1181.670 427.680 ;
        RECT 1181.155 427.480 1181.670 427.620 ;
        RECT 1181.350 427.420 1181.670 427.480 ;
        RECT 1181.350 379.680 1181.670 379.740 ;
        RECT 1181.155 379.540 1181.670 379.680 ;
        RECT 1181.350 379.480 1181.670 379.540 ;
        RECT 1181.350 351.800 1181.670 351.860 ;
        RECT 1181.155 351.660 1181.670 351.800 ;
        RECT 1181.350 351.600 1181.670 351.660 ;
        RECT 1181.350 338.200 1181.670 338.260 ;
        RECT 1181.155 338.060 1181.670 338.200 ;
        RECT 1181.350 338.000 1181.670 338.060 ;
        RECT 1181.350 331.060 1181.670 331.120 ;
        RECT 1181.825 331.060 1182.115 331.105 ;
        RECT 1181.350 330.920 1182.115 331.060 ;
        RECT 1181.350 330.860 1181.670 330.920 ;
        RECT 1181.825 330.875 1182.115 330.920 ;
        RECT 1181.350 235.180 1181.670 235.240 ;
        RECT 1181.825 235.180 1182.115 235.225 ;
        RECT 1181.350 235.040 1182.115 235.180 ;
        RECT 1181.350 234.980 1181.670 235.040 ;
        RECT 1181.825 234.995 1182.115 235.040 ;
        RECT 1181.350 234.500 1181.670 234.560 ;
        RECT 1182.270 234.500 1182.590 234.560 ;
        RECT 1181.350 234.360 1182.590 234.500 ;
        RECT 1181.350 234.300 1181.670 234.360 ;
        RECT 1182.270 234.300 1182.590 234.360 ;
        RECT 1181.350 145.080 1181.670 145.140 ;
        RECT 1181.810 145.080 1182.130 145.140 ;
        RECT 1181.350 144.940 1182.130 145.080 ;
        RECT 1181.350 144.880 1181.670 144.940 ;
        RECT 1181.810 144.880 1182.130 144.940 ;
        RECT 1181.350 96.600 1181.670 96.860 ;
        RECT 1181.440 96.120 1181.580 96.600 ;
        RECT 1181.810 96.120 1182.130 96.180 ;
        RECT 1181.440 95.980 1182.130 96.120 ;
        RECT 1181.810 95.920 1182.130 95.980 ;
        RECT 74.130 17.580 74.450 17.640 ;
        RECT 1181.810 17.580 1182.130 17.640 ;
        RECT 74.130 17.440 1182.130 17.580 ;
        RECT 74.130 17.380 74.450 17.440 ;
        RECT 1181.810 17.380 1182.130 17.440 ;
      LAYER via ;
        RECT 1181.380 1635.440 1181.640 1635.700 ;
        RECT 1184.600 1635.440 1184.860 1635.700 ;
        RECT 1181.380 1545.340 1181.640 1545.600 ;
        RECT 1181.840 1545.340 1182.100 1545.600 ;
        RECT 1181.380 1490.260 1181.640 1490.520 ;
        RECT 1182.300 1448.440 1182.560 1448.700 ;
        RECT 1181.840 1393.700 1182.100 1393.960 ;
        RECT 1183.220 1393.700 1183.480 1393.960 ;
        RECT 1181.840 1352.560 1182.100 1352.820 ;
        RECT 1181.380 1352.220 1181.640 1352.480 ;
        RECT 1181.380 1317.880 1181.640 1318.140 ;
        RECT 1181.840 1317.540 1182.100 1317.800 ;
        RECT 1181.840 1269.260 1182.100 1269.520 ;
        RECT 1181.380 1268.580 1181.640 1268.840 ;
        RECT 1181.380 1221.320 1181.640 1221.580 ;
        RECT 1181.380 1200.920 1181.640 1201.180 ;
        RECT 1181.380 1200.240 1181.640 1200.500 ;
        RECT 1181.380 1152.640 1181.640 1152.900 ;
        RECT 1181.380 1104.020 1181.640 1104.280 ;
        RECT 1182.300 1104.020 1182.560 1104.280 ;
        RECT 1181.840 1079.880 1182.100 1080.140 ;
        RECT 1182.760 1079.880 1183.020 1080.140 ;
        RECT 1181.380 1027.860 1181.640 1028.120 ;
        RECT 1181.380 1014.260 1181.640 1014.520 ;
        RECT 1181.380 993.180 1181.640 993.440 ;
        RECT 1181.840 945.240 1182.100 945.500 ;
        RECT 1181.840 896.620 1182.100 896.880 ;
        RECT 1181.840 807.200 1182.100 807.460 ;
        RECT 1181.380 765.720 1181.640 765.980 ;
        RECT 1181.840 765.720 1182.100 765.980 ;
        RECT 1181.380 717.440 1181.640 717.700 ;
        RECT 1182.300 717.440 1182.560 717.700 ;
        RECT 1182.300 710.300 1182.560 710.560 ;
        RECT 1182.300 662.360 1182.560 662.620 ;
        RECT 1181.840 621.220 1182.100 621.480 ;
        RECT 1182.300 621.220 1182.560 621.480 ;
        RECT 1181.840 613.740 1182.100 614.000 ;
        RECT 1182.300 565.800 1182.560 566.060 ;
        RECT 1181.380 530.780 1181.640 531.040 ;
        RECT 1182.760 530.780 1183.020 531.040 ;
        RECT 1181.380 427.420 1181.640 427.680 ;
        RECT 1181.380 379.480 1181.640 379.740 ;
        RECT 1181.380 351.600 1181.640 351.860 ;
        RECT 1181.380 338.000 1181.640 338.260 ;
        RECT 1181.380 330.860 1181.640 331.120 ;
        RECT 1181.380 234.980 1181.640 235.240 ;
        RECT 1181.380 234.300 1181.640 234.560 ;
        RECT 1182.300 234.300 1182.560 234.560 ;
        RECT 1181.380 144.880 1181.640 145.140 ;
        RECT 1181.840 144.880 1182.100 145.140 ;
        RECT 1181.380 96.600 1181.640 96.860 ;
        RECT 1181.840 95.920 1182.100 96.180 ;
        RECT 74.160 17.380 74.420 17.640 ;
        RECT 1181.840 17.380 1182.100 17.640 ;
      LAYER met2 ;
        RECT 1186.360 1700.410 1186.640 1702.400 ;
        RECT 1184.660 1700.270 1186.640 1700.410 ;
        RECT 1184.660 1635.730 1184.800 1700.270 ;
        RECT 1186.360 1700.000 1186.640 1700.270 ;
        RECT 1181.380 1635.410 1181.640 1635.730 ;
        RECT 1184.600 1635.410 1184.860 1635.730 ;
        RECT 1181.440 1607.250 1181.580 1635.410 ;
        RECT 1181.440 1607.110 1182.040 1607.250 ;
        RECT 1181.900 1545.630 1182.040 1607.110 ;
        RECT 1181.380 1545.310 1181.640 1545.630 ;
        RECT 1181.840 1545.310 1182.100 1545.630 ;
        RECT 1181.440 1490.550 1181.580 1545.310 ;
        RECT 1181.380 1490.230 1181.640 1490.550 ;
        RECT 1182.300 1448.410 1182.560 1448.730 ;
        RECT 1182.360 1442.125 1182.500 1448.410 ;
        RECT 1182.290 1441.755 1182.570 1442.125 ;
        RECT 1183.210 1441.755 1183.490 1442.125 ;
        RECT 1181.900 1393.990 1182.040 1394.145 ;
        RECT 1183.280 1393.990 1183.420 1441.755 ;
        RECT 1181.840 1393.730 1182.100 1393.990 ;
        RECT 1181.440 1393.670 1182.100 1393.730 ;
        RECT 1183.220 1393.670 1183.480 1393.990 ;
        RECT 1181.440 1393.590 1182.040 1393.670 ;
        RECT 1181.440 1386.930 1181.580 1393.590 ;
        RECT 1181.440 1386.790 1182.040 1386.930 ;
        RECT 1181.900 1352.850 1182.040 1386.790 ;
        RECT 1181.840 1352.530 1182.100 1352.850 ;
        RECT 1181.380 1352.190 1181.640 1352.510 ;
        RECT 1181.440 1318.170 1181.580 1352.190 ;
        RECT 1181.380 1317.850 1181.640 1318.170 ;
        RECT 1181.840 1317.510 1182.100 1317.830 ;
        RECT 1181.900 1269.550 1182.040 1317.510 ;
        RECT 1181.840 1269.230 1182.100 1269.550 ;
        RECT 1181.380 1268.550 1181.640 1268.870 ;
        RECT 1181.440 1221.610 1181.580 1268.550 ;
        RECT 1181.380 1221.290 1181.640 1221.610 ;
        RECT 1181.380 1200.890 1181.640 1201.210 ;
        RECT 1181.440 1200.530 1181.580 1200.890 ;
        RECT 1181.380 1200.210 1181.640 1200.530 ;
        RECT 1181.380 1152.610 1181.640 1152.930 ;
        RECT 1181.440 1152.445 1181.580 1152.610 ;
        RECT 1181.370 1152.075 1181.650 1152.445 ;
        RECT 1182.290 1152.075 1182.570 1152.445 ;
        RECT 1181.440 1104.310 1181.580 1104.465 ;
        RECT 1182.360 1104.310 1182.500 1152.075 ;
        RECT 1181.380 1104.050 1181.640 1104.310 ;
        RECT 1181.380 1103.990 1182.040 1104.050 ;
        RECT 1182.300 1103.990 1182.560 1104.310 ;
        RECT 1181.440 1103.910 1182.040 1103.990 ;
        RECT 1181.900 1080.170 1182.040 1103.910 ;
        RECT 1181.840 1079.850 1182.100 1080.170 ;
        RECT 1182.760 1079.850 1183.020 1080.170 ;
        RECT 1182.820 1055.885 1182.960 1079.850 ;
        RECT 1181.370 1055.515 1181.650 1055.885 ;
        RECT 1182.750 1055.515 1183.030 1055.885 ;
        RECT 1181.440 1028.150 1181.580 1055.515 ;
        RECT 1181.380 1027.830 1181.640 1028.150 ;
        RECT 1181.380 1014.230 1181.640 1014.550 ;
        RECT 1181.440 993.470 1181.580 1014.230 ;
        RECT 1181.380 993.150 1181.640 993.470 ;
        RECT 1181.840 945.210 1182.100 945.530 ;
        RECT 1181.900 896.910 1182.040 945.210 ;
        RECT 1181.840 896.590 1182.100 896.910 ;
        RECT 1181.840 807.170 1182.100 807.490 ;
        RECT 1181.900 766.010 1182.040 807.170 ;
        RECT 1181.380 765.690 1181.640 766.010 ;
        RECT 1181.840 765.690 1182.100 766.010 ;
        RECT 1181.440 717.730 1181.580 765.690 ;
        RECT 1181.380 717.410 1181.640 717.730 ;
        RECT 1182.300 717.410 1182.560 717.730 ;
        RECT 1182.360 710.590 1182.500 717.410 ;
        RECT 1182.300 710.270 1182.560 710.590 ;
        RECT 1182.300 662.330 1182.560 662.650 ;
        RECT 1182.360 621.510 1182.500 662.330 ;
        RECT 1181.840 621.190 1182.100 621.510 ;
        RECT 1182.300 621.190 1182.560 621.510 ;
        RECT 1181.900 614.030 1182.040 621.190 ;
        RECT 1181.840 613.710 1182.100 614.030 ;
        RECT 1182.300 565.770 1182.560 566.090 ;
        RECT 1182.360 531.605 1182.500 565.770 ;
        RECT 1181.370 531.235 1181.650 531.605 ;
        RECT 1182.290 531.235 1182.570 531.605 ;
        RECT 1181.440 531.070 1181.580 531.235 ;
        RECT 1181.380 530.750 1181.640 531.070 ;
        RECT 1182.760 530.750 1183.020 531.070 ;
        RECT 1182.820 483.325 1182.960 530.750 ;
        RECT 1181.830 482.955 1182.110 483.325 ;
        RECT 1182.750 482.955 1183.030 483.325 ;
        RECT 1181.900 435.725 1182.040 482.955 ;
        RECT 1181.830 435.355 1182.110 435.725 ;
        RECT 1181.370 434.675 1181.650 435.045 ;
        RECT 1181.440 427.710 1181.580 434.675 ;
        RECT 1181.380 427.390 1181.640 427.710 ;
        RECT 1181.380 379.450 1181.640 379.770 ;
        RECT 1181.440 351.890 1181.580 379.450 ;
        RECT 1181.380 351.570 1181.640 351.890 ;
        RECT 1181.380 337.970 1181.640 338.290 ;
        RECT 1181.440 331.150 1181.580 337.970 ;
        RECT 1181.380 330.830 1181.640 331.150 ;
        RECT 1181.380 234.950 1181.640 235.270 ;
        RECT 1181.440 234.590 1181.580 234.950 ;
        RECT 1181.380 234.270 1181.640 234.590 ;
        RECT 1182.300 234.270 1182.560 234.590 ;
        RECT 1182.360 206.450 1182.500 234.270 ;
        RECT 1181.900 206.310 1182.500 206.450 ;
        RECT 1181.900 145.170 1182.040 206.310 ;
        RECT 1181.380 144.850 1181.640 145.170 ;
        RECT 1181.840 144.850 1182.100 145.170 ;
        RECT 1181.440 96.890 1181.580 144.850 ;
        RECT 1181.380 96.570 1181.640 96.890 ;
        RECT 1181.840 95.890 1182.100 96.210 ;
        RECT 1181.900 17.670 1182.040 95.890 ;
        RECT 74.160 17.350 74.420 17.670 ;
        RECT 1181.840 17.350 1182.100 17.670 ;
        RECT 74.220 2.400 74.360 17.350 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 1182.290 1441.800 1182.570 1442.080 ;
        RECT 1183.210 1441.800 1183.490 1442.080 ;
        RECT 1181.370 1152.120 1181.650 1152.400 ;
        RECT 1182.290 1152.120 1182.570 1152.400 ;
        RECT 1181.370 1055.560 1181.650 1055.840 ;
        RECT 1182.750 1055.560 1183.030 1055.840 ;
        RECT 1181.370 531.280 1181.650 531.560 ;
        RECT 1182.290 531.280 1182.570 531.560 ;
        RECT 1181.830 483.000 1182.110 483.280 ;
        RECT 1182.750 483.000 1183.030 483.280 ;
        RECT 1181.830 435.400 1182.110 435.680 ;
        RECT 1181.370 434.720 1181.650 435.000 ;
      LAYER met3 ;
        RECT 1182.265 1442.090 1182.595 1442.105 ;
        RECT 1183.185 1442.090 1183.515 1442.105 ;
        RECT 1182.265 1441.790 1183.515 1442.090 ;
        RECT 1182.265 1441.775 1182.595 1441.790 ;
        RECT 1183.185 1441.775 1183.515 1441.790 ;
        RECT 1181.345 1152.410 1181.675 1152.425 ;
        RECT 1182.265 1152.410 1182.595 1152.425 ;
        RECT 1181.345 1152.110 1182.595 1152.410 ;
        RECT 1181.345 1152.095 1181.675 1152.110 ;
        RECT 1182.265 1152.095 1182.595 1152.110 ;
        RECT 1181.345 1055.850 1181.675 1055.865 ;
        RECT 1182.725 1055.850 1183.055 1055.865 ;
        RECT 1181.345 1055.550 1183.055 1055.850 ;
        RECT 1181.345 1055.535 1181.675 1055.550 ;
        RECT 1182.725 1055.535 1183.055 1055.550 ;
        RECT 1181.345 531.570 1181.675 531.585 ;
        RECT 1182.265 531.570 1182.595 531.585 ;
        RECT 1181.345 531.270 1182.595 531.570 ;
        RECT 1181.345 531.255 1181.675 531.270 ;
        RECT 1182.265 531.255 1182.595 531.270 ;
        RECT 1181.805 483.290 1182.135 483.305 ;
        RECT 1182.725 483.290 1183.055 483.305 ;
        RECT 1181.805 482.990 1183.055 483.290 ;
        RECT 1181.805 482.975 1182.135 482.990 ;
        RECT 1182.725 482.975 1183.055 482.990 ;
        RECT 1181.805 435.690 1182.135 435.705 ;
        RECT 1180.670 435.390 1182.135 435.690 ;
        RECT 1180.670 435.010 1180.970 435.390 ;
        RECT 1181.805 435.375 1182.135 435.390 ;
        RECT 1181.345 435.010 1181.675 435.025 ;
        RECT 1180.670 434.710 1181.675 435.010 ;
        RECT 1181.345 434.695 1181.675 434.710 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 493.265 14.025 493.435 14.875 ;
      LAYER mcon ;
        RECT 493.265 14.705 493.435 14.875 ;
      LAYER met1 ;
        RECT 527.690 1684.260 528.010 1684.320 ;
        RECT 1370.410 1684.260 1370.730 1684.320 ;
        RECT 527.690 1684.120 1370.730 1684.260 ;
        RECT 527.690 1684.060 528.010 1684.120 ;
        RECT 1370.410 1684.060 1370.730 1684.120 ;
        RECT 430.630 14.860 430.950 14.920 ;
        RECT 493.205 14.860 493.495 14.905 ;
        RECT 430.630 14.720 493.495 14.860 ;
        RECT 430.630 14.660 430.950 14.720 ;
        RECT 493.205 14.675 493.495 14.720 ;
        RECT 493.205 14.180 493.495 14.225 ;
        RECT 527.690 14.180 528.010 14.240 ;
        RECT 493.205 14.040 528.010 14.180 ;
        RECT 493.205 13.995 493.495 14.040 ;
        RECT 527.690 13.980 528.010 14.040 ;
      LAYER via ;
        RECT 527.720 1684.060 527.980 1684.320 ;
        RECT 1370.440 1684.060 1370.700 1684.320 ;
        RECT 430.660 14.660 430.920 14.920 ;
        RECT 527.720 13.980 527.980 14.240 ;
      LAYER met2 ;
        RECT 1370.360 1700.000 1370.640 1702.400 ;
        RECT 1370.500 1684.350 1370.640 1700.000 ;
        RECT 527.720 1684.030 527.980 1684.350 ;
        RECT 1370.440 1684.030 1370.700 1684.350 ;
        RECT 430.660 14.630 430.920 14.950 ;
        RECT 430.720 2.400 430.860 14.630 ;
        RECT 527.780 14.270 527.920 1684.030 ;
        RECT 527.720 13.950 527.980 14.270 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1337.365 1686.825 1337.535 1687.675 ;
      LAYER mcon ;
        RECT 1337.365 1687.505 1337.535 1687.675 ;
      LAYER met1 ;
        RECT 1314.290 1687.660 1314.610 1687.720 ;
        RECT 1337.305 1687.660 1337.595 1687.705 ;
        RECT 1314.290 1687.520 1337.595 1687.660 ;
        RECT 1314.290 1687.460 1314.610 1687.520 ;
        RECT 1337.305 1687.475 1337.595 1687.520 ;
        RECT 1337.305 1686.980 1337.595 1687.025 ;
        RECT 1379.610 1686.980 1379.930 1687.040 ;
        RECT 1337.305 1686.840 1379.930 1686.980 ;
        RECT 1337.305 1686.795 1337.595 1686.840 ;
        RECT 1379.610 1686.780 1379.930 1686.840 ;
        RECT 449.030 15.880 449.350 15.940 ;
        RECT 1314.290 15.880 1314.610 15.940 ;
        RECT 449.030 15.740 1314.610 15.880 ;
        RECT 449.030 15.680 449.350 15.740 ;
        RECT 1314.290 15.680 1314.610 15.740 ;
      LAYER via ;
        RECT 1314.320 1687.460 1314.580 1687.720 ;
        RECT 1379.640 1686.780 1379.900 1687.040 ;
        RECT 449.060 15.680 449.320 15.940 ;
        RECT 1314.320 15.680 1314.580 15.940 ;
      LAYER met2 ;
        RECT 1379.560 1700.000 1379.840 1702.400 ;
        RECT 1314.320 1687.430 1314.580 1687.750 ;
        RECT 1314.380 15.970 1314.520 1687.430 ;
        RECT 1379.700 1687.070 1379.840 1700.000 ;
        RECT 1379.640 1686.750 1379.900 1687.070 ;
        RECT 449.060 15.650 449.320 15.970 ;
        RECT 1314.320 15.650 1314.580 15.970 ;
        RECT 449.120 7.890 449.260 15.650 ;
        RECT 448.660 7.750 449.260 7.890 ;
        RECT 448.660 2.400 448.800 7.750 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 486.290 1685.960 486.610 1686.020 ;
        RECT 1388.810 1685.960 1389.130 1686.020 ;
        RECT 486.290 1685.820 1389.130 1685.960 ;
        RECT 486.290 1685.760 486.610 1685.820 ;
        RECT 1388.810 1685.760 1389.130 1685.820 ;
        RECT 486.290 15.540 486.610 15.600 ;
        RECT 483.160 15.400 486.610 15.540 ;
        RECT 466.510 15.200 466.830 15.260 ;
        RECT 483.160 15.200 483.300 15.400 ;
        RECT 486.290 15.340 486.610 15.400 ;
        RECT 466.510 15.060 483.300 15.200 ;
        RECT 466.510 15.000 466.830 15.060 ;
      LAYER via ;
        RECT 486.320 1685.760 486.580 1686.020 ;
        RECT 1388.840 1685.760 1389.100 1686.020 ;
        RECT 466.540 15.000 466.800 15.260 ;
        RECT 486.320 15.340 486.580 15.600 ;
      LAYER met2 ;
        RECT 1388.760 1700.000 1389.040 1702.400 ;
        RECT 1388.900 1686.050 1389.040 1700.000 ;
        RECT 486.320 1685.730 486.580 1686.050 ;
        RECT 1388.840 1685.730 1389.100 1686.050 ;
        RECT 486.380 15.630 486.520 1685.730 ;
        RECT 486.320 15.310 486.580 15.630 ;
        RECT 466.540 14.970 466.800 15.290 ;
        RECT 466.600 2.400 466.740 14.970 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1321.190 1687.320 1321.510 1687.380 ;
        RECT 1398.010 1687.320 1398.330 1687.380 ;
        RECT 1321.190 1687.180 1398.330 1687.320 ;
        RECT 1321.190 1687.120 1321.510 1687.180 ;
        RECT 1398.010 1687.120 1398.330 1687.180 ;
        RECT 1321.190 15.540 1321.510 15.600 ;
        RECT 559.060 15.400 1321.510 15.540 ;
        RECT 484.450 15.200 484.770 15.260 ;
        RECT 559.060 15.200 559.200 15.400 ;
        RECT 1321.190 15.340 1321.510 15.400 ;
        RECT 484.450 15.060 493.880 15.200 ;
        RECT 484.450 15.000 484.770 15.060 ;
        RECT 493.740 14.860 493.880 15.060 ;
        RECT 496.960 15.060 559.200 15.200 ;
        RECT 496.960 14.860 497.100 15.060 ;
        RECT 493.740 14.720 497.100 14.860 ;
      LAYER via ;
        RECT 1321.220 1687.120 1321.480 1687.380 ;
        RECT 1398.040 1687.120 1398.300 1687.380 ;
        RECT 484.480 15.000 484.740 15.260 ;
        RECT 1321.220 15.340 1321.480 15.600 ;
      LAYER met2 ;
        RECT 1397.960 1700.000 1398.240 1702.400 ;
        RECT 1398.100 1687.410 1398.240 1700.000 ;
        RECT 1321.220 1687.090 1321.480 1687.410 ;
        RECT 1398.040 1687.090 1398.300 1687.410 ;
        RECT 1321.280 15.630 1321.420 1687.090 ;
        RECT 1321.220 15.310 1321.480 15.630 ;
        RECT 484.480 14.970 484.740 15.290 ;
        RECT 484.540 2.400 484.680 14.970 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1321.650 1688.340 1321.970 1688.400 ;
        RECT 1407.210 1688.340 1407.530 1688.400 ;
        RECT 1321.650 1688.200 1407.530 1688.340 ;
        RECT 1321.650 1688.140 1321.970 1688.200 ;
        RECT 1407.210 1688.140 1407.530 1688.200 ;
        RECT 1321.650 15.200 1321.970 15.260 ;
        RECT 559.520 15.060 1321.970 15.200 ;
        RECT 502.390 14.520 502.710 14.580 ;
        RECT 559.520 14.520 559.660 15.060 ;
        RECT 1321.650 15.000 1321.970 15.060 ;
        RECT 502.390 14.380 559.660 14.520 ;
        RECT 502.390 14.320 502.710 14.380 ;
      LAYER via ;
        RECT 1321.680 1688.140 1321.940 1688.400 ;
        RECT 1407.240 1688.140 1407.500 1688.400 ;
        RECT 502.420 14.320 502.680 14.580 ;
        RECT 1321.680 15.000 1321.940 15.260 ;
      LAYER met2 ;
        RECT 1407.160 1700.000 1407.440 1702.400 ;
        RECT 1407.300 1688.430 1407.440 1700.000 ;
        RECT 1321.680 1688.110 1321.940 1688.430 ;
        RECT 1407.240 1688.110 1407.500 1688.430 ;
        RECT 1321.740 15.290 1321.880 1688.110 ;
        RECT 1321.680 14.970 1321.940 15.290 ;
        RECT 502.420 14.290 502.680 14.610 ;
        RECT 502.480 2.400 502.620 14.290 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 1685.620 524.330 1685.680 ;
        RECT 1415.950 1685.620 1416.270 1685.680 ;
        RECT 524.010 1685.480 1416.270 1685.620 ;
        RECT 524.010 1685.420 524.330 1685.480 ;
        RECT 1415.950 1685.420 1416.270 1685.480 ;
        RECT 519.870 15.540 520.190 15.600 ;
        RECT 524.010 15.540 524.330 15.600 ;
        RECT 519.870 15.400 524.330 15.540 ;
        RECT 519.870 15.340 520.190 15.400 ;
        RECT 524.010 15.340 524.330 15.400 ;
      LAYER via ;
        RECT 524.040 1685.420 524.300 1685.680 ;
        RECT 1415.980 1685.420 1416.240 1685.680 ;
        RECT 519.900 15.340 520.160 15.600 ;
        RECT 524.040 15.340 524.300 15.600 ;
      LAYER met2 ;
        RECT 1415.900 1700.000 1416.180 1702.400 ;
        RECT 1416.040 1685.710 1416.180 1700.000 ;
        RECT 524.040 1685.390 524.300 1685.710 ;
        RECT 1415.980 1685.390 1416.240 1685.710 ;
        RECT 524.100 15.630 524.240 1685.390 ;
        RECT 519.900 15.310 520.160 15.630 ;
        RECT 524.040 15.310 524.300 15.630 ;
        RECT 519.960 2.400 520.100 15.310 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1337.825 1642.285 1337.995 1687.675 ;
        RECT 1335.525 1538.925 1335.695 1545.895 ;
        RECT 1335.065 1400.885 1335.235 1490.475 ;
        RECT 1335.065 1297.185 1335.235 1318.095 ;
        RECT 1335.525 1104.065 1335.695 1124.975 ;
        RECT 1335.065 1048.985 1335.235 1097.095 ;
        RECT 1335.065 765.765 1335.235 787.355 ;
        RECT 1335.065 524.705 1335.235 572.475 ;
        RECT 1335.065 476.085 1335.235 524.195 ;
        RECT 1335.065 179.605 1335.235 227.715 ;
      LAYER mcon ;
        RECT 1337.825 1687.505 1337.995 1687.675 ;
        RECT 1335.525 1545.725 1335.695 1545.895 ;
        RECT 1335.065 1490.305 1335.235 1490.475 ;
        RECT 1335.065 1317.925 1335.235 1318.095 ;
        RECT 1335.525 1124.805 1335.695 1124.975 ;
        RECT 1335.065 1096.925 1335.235 1097.095 ;
        RECT 1335.065 787.185 1335.235 787.355 ;
        RECT 1335.065 572.305 1335.235 572.475 ;
        RECT 1335.065 524.025 1335.235 524.195 ;
        RECT 1335.065 227.545 1335.235 227.715 ;
      LAYER met1 ;
        RECT 1337.765 1687.660 1338.055 1687.705 ;
        RECT 1425.150 1687.660 1425.470 1687.720 ;
        RECT 1337.765 1687.520 1425.470 1687.660 ;
        RECT 1337.765 1687.475 1338.055 1687.520 ;
        RECT 1425.150 1687.460 1425.470 1687.520 ;
        RECT 1335.450 1642.440 1335.770 1642.500 ;
        RECT 1337.765 1642.440 1338.055 1642.485 ;
        RECT 1335.450 1642.300 1338.055 1642.440 ;
        RECT 1335.450 1642.240 1335.770 1642.300 ;
        RECT 1337.765 1642.255 1338.055 1642.300 ;
        RECT 1335.450 1545.880 1335.770 1545.940 ;
        RECT 1335.255 1545.740 1335.770 1545.880 ;
        RECT 1335.450 1545.680 1335.770 1545.740 ;
        RECT 1335.450 1539.080 1335.770 1539.140 ;
        RECT 1335.255 1538.940 1335.770 1539.080 ;
        RECT 1335.450 1538.880 1335.770 1538.940 ;
        RECT 1335.005 1490.460 1335.295 1490.505 ;
        RECT 1335.450 1490.460 1335.770 1490.520 ;
        RECT 1335.005 1490.320 1335.770 1490.460 ;
        RECT 1335.005 1490.275 1335.295 1490.320 ;
        RECT 1335.450 1490.260 1335.770 1490.320 ;
        RECT 1334.990 1401.040 1335.310 1401.100 ;
        RECT 1334.795 1400.900 1335.310 1401.040 ;
        RECT 1334.990 1400.840 1335.310 1400.900 ;
        RECT 1334.990 1352.760 1335.310 1352.820 ;
        RECT 1335.450 1352.760 1335.770 1352.820 ;
        RECT 1334.990 1352.620 1335.770 1352.760 ;
        RECT 1334.990 1352.560 1335.310 1352.620 ;
        RECT 1335.450 1352.560 1335.770 1352.620 ;
        RECT 1334.990 1318.080 1335.310 1318.140 ;
        RECT 1334.795 1317.940 1335.310 1318.080 ;
        RECT 1334.990 1317.880 1335.310 1317.940 ;
        RECT 1334.990 1297.340 1335.310 1297.400 ;
        RECT 1334.795 1297.200 1335.310 1297.340 ;
        RECT 1334.990 1297.140 1335.310 1297.200 ;
        RECT 1335.450 1124.960 1335.770 1125.020 ;
        RECT 1335.255 1124.820 1335.770 1124.960 ;
        RECT 1335.450 1124.760 1335.770 1124.820 ;
        RECT 1335.450 1104.220 1335.770 1104.280 ;
        RECT 1335.255 1104.080 1335.770 1104.220 ;
        RECT 1335.450 1104.020 1335.770 1104.080 ;
        RECT 1335.005 1097.080 1335.295 1097.125 ;
        RECT 1335.450 1097.080 1335.770 1097.140 ;
        RECT 1335.005 1096.940 1335.770 1097.080 ;
        RECT 1335.005 1096.895 1335.295 1096.940 ;
        RECT 1335.450 1096.880 1335.770 1096.940 ;
        RECT 1334.990 1049.140 1335.310 1049.200 ;
        RECT 1334.795 1049.000 1335.310 1049.140 ;
        RECT 1334.990 1048.940 1335.310 1049.000 ;
        RECT 1334.990 966.180 1335.310 966.240 ;
        RECT 1335.450 966.180 1335.770 966.240 ;
        RECT 1334.990 966.040 1335.770 966.180 ;
        RECT 1334.990 965.980 1335.310 966.040 ;
        RECT 1335.450 965.980 1335.770 966.040 ;
        RECT 1335.450 932.180 1335.770 932.240 ;
        RECT 1335.080 932.040 1335.770 932.180 ;
        RECT 1335.080 931.560 1335.220 932.040 ;
        RECT 1335.450 931.980 1335.770 932.040 ;
        RECT 1334.990 931.300 1335.310 931.560 ;
        RECT 1334.990 787.340 1335.310 787.400 ;
        RECT 1334.795 787.200 1335.310 787.340 ;
        RECT 1334.990 787.140 1335.310 787.200 ;
        RECT 1334.990 765.920 1335.310 765.980 ;
        RECT 1334.795 765.780 1335.310 765.920 ;
        RECT 1334.990 765.720 1335.310 765.780 ;
        RECT 1334.990 717.980 1335.310 718.040 ;
        RECT 1335.450 717.980 1335.770 718.040 ;
        RECT 1334.990 717.840 1335.770 717.980 ;
        RECT 1334.990 717.780 1335.310 717.840 ;
        RECT 1335.450 717.780 1335.770 717.840 ;
        RECT 1334.990 627.880 1335.310 627.940 ;
        RECT 1336.370 627.880 1336.690 627.940 ;
        RECT 1334.990 627.740 1336.690 627.880 ;
        RECT 1334.990 627.680 1335.310 627.740 ;
        RECT 1336.370 627.680 1336.690 627.740 ;
        RECT 1335.005 572.460 1335.295 572.505 ;
        RECT 1335.450 572.460 1335.770 572.520 ;
        RECT 1335.005 572.320 1335.770 572.460 ;
        RECT 1335.005 572.275 1335.295 572.320 ;
        RECT 1335.450 572.260 1335.770 572.320 ;
        RECT 1334.990 524.860 1335.310 524.920 ;
        RECT 1334.795 524.720 1335.310 524.860 ;
        RECT 1334.990 524.660 1335.310 524.720 ;
        RECT 1334.990 524.180 1335.310 524.240 ;
        RECT 1334.795 524.040 1335.310 524.180 ;
        RECT 1334.990 523.980 1335.310 524.040 ;
        RECT 1335.005 476.240 1335.295 476.285 ;
        RECT 1335.450 476.240 1335.770 476.300 ;
        RECT 1335.005 476.100 1335.770 476.240 ;
        RECT 1335.005 476.055 1335.295 476.100 ;
        RECT 1335.450 476.040 1335.770 476.100 ;
        RECT 1335.450 372.880 1335.770 372.940 ;
        RECT 1336.370 372.880 1336.690 372.940 ;
        RECT 1335.450 372.740 1336.690 372.880 ;
        RECT 1335.450 372.680 1335.770 372.740 ;
        RECT 1336.370 372.680 1336.690 372.740 ;
        RECT 1336.370 338.540 1336.690 338.600 ;
        RECT 1336.000 338.400 1336.690 338.540 ;
        RECT 1336.000 337.920 1336.140 338.400 ;
        RECT 1336.370 338.340 1336.690 338.400 ;
        RECT 1335.910 337.660 1336.230 337.920 ;
        RECT 1335.450 289.920 1335.770 289.980 ;
        RECT 1335.910 289.920 1336.230 289.980 ;
        RECT 1335.450 289.780 1336.230 289.920 ;
        RECT 1335.450 289.720 1335.770 289.780 ;
        RECT 1335.910 289.720 1336.230 289.780 ;
        RECT 1334.990 234.500 1335.310 234.560 ;
        RECT 1335.910 234.500 1336.230 234.560 ;
        RECT 1334.990 234.360 1336.230 234.500 ;
        RECT 1334.990 234.300 1335.310 234.360 ;
        RECT 1335.910 234.300 1336.230 234.360 ;
        RECT 1335.005 227.700 1335.295 227.745 ;
        RECT 1335.910 227.700 1336.230 227.760 ;
        RECT 1335.005 227.560 1336.230 227.700 ;
        RECT 1335.005 227.515 1335.295 227.560 ;
        RECT 1335.910 227.500 1336.230 227.560 ;
        RECT 1334.990 179.760 1335.310 179.820 ;
        RECT 1334.795 179.620 1335.310 179.760 ;
        RECT 1334.990 179.560 1335.310 179.620 ;
        RECT 1334.990 137.940 1335.310 138.000 ;
        RECT 1335.450 137.940 1335.770 138.000 ;
        RECT 1334.990 137.800 1335.770 137.940 ;
        RECT 1334.990 137.740 1335.310 137.800 ;
        RECT 1335.450 137.740 1335.770 137.800 ;
        RECT 1334.530 14.860 1334.850 14.920 ;
        RECT 607.820 14.720 1334.850 14.860 ;
        RECT 537.810 14.180 538.130 14.240 ;
        RECT 607.820 14.180 607.960 14.720 ;
        RECT 1334.530 14.660 1334.850 14.720 ;
        RECT 537.810 14.040 607.960 14.180 ;
        RECT 537.810 13.980 538.130 14.040 ;
      LAYER via ;
        RECT 1425.180 1687.460 1425.440 1687.720 ;
        RECT 1335.480 1642.240 1335.740 1642.500 ;
        RECT 1335.480 1545.680 1335.740 1545.940 ;
        RECT 1335.480 1538.880 1335.740 1539.140 ;
        RECT 1335.480 1490.260 1335.740 1490.520 ;
        RECT 1335.020 1400.840 1335.280 1401.100 ;
        RECT 1335.020 1352.560 1335.280 1352.820 ;
        RECT 1335.480 1352.560 1335.740 1352.820 ;
        RECT 1335.020 1317.880 1335.280 1318.140 ;
        RECT 1335.020 1297.140 1335.280 1297.400 ;
        RECT 1335.480 1124.760 1335.740 1125.020 ;
        RECT 1335.480 1104.020 1335.740 1104.280 ;
        RECT 1335.480 1096.880 1335.740 1097.140 ;
        RECT 1335.020 1048.940 1335.280 1049.200 ;
        RECT 1335.020 965.980 1335.280 966.240 ;
        RECT 1335.480 965.980 1335.740 966.240 ;
        RECT 1335.480 931.980 1335.740 932.240 ;
        RECT 1335.020 931.300 1335.280 931.560 ;
        RECT 1335.020 787.140 1335.280 787.400 ;
        RECT 1335.020 765.720 1335.280 765.980 ;
        RECT 1335.020 717.780 1335.280 718.040 ;
        RECT 1335.480 717.780 1335.740 718.040 ;
        RECT 1335.020 627.680 1335.280 627.940 ;
        RECT 1336.400 627.680 1336.660 627.940 ;
        RECT 1335.480 572.260 1335.740 572.520 ;
        RECT 1335.020 524.660 1335.280 524.920 ;
        RECT 1335.020 523.980 1335.280 524.240 ;
        RECT 1335.480 476.040 1335.740 476.300 ;
        RECT 1335.480 372.680 1335.740 372.940 ;
        RECT 1336.400 372.680 1336.660 372.940 ;
        RECT 1336.400 338.340 1336.660 338.600 ;
        RECT 1335.940 337.660 1336.200 337.920 ;
        RECT 1335.480 289.720 1335.740 289.980 ;
        RECT 1335.940 289.720 1336.200 289.980 ;
        RECT 1335.020 234.300 1335.280 234.560 ;
        RECT 1335.940 234.300 1336.200 234.560 ;
        RECT 1335.940 227.500 1336.200 227.760 ;
        RECT 1335.020 179.560 1335.280 179.820 ;
        RECT 1335.020 137.740 1335.280 138.000 ;
        RECT 1335.480 137.740 1335.740 138.000 ;
        RECT 537.840 13.980 538.100 14.240 ;
        RECT 1334.560 14.660 1334.820 14.920 ;
      LAYER met2 ;
        RECT 1425.100 1700.000 1425.380 1702.400 ;
        RECT 1425.240 1687.750 1425.380 1700.000 ;
        RECT 1425.180 1687.430 1425.440 1687.750 ;
        RECT 1335.480 1642.210 1335.740 1642.530 ;
        RECT 1335.540 1545.970 1335.680 1642.210 ;
        RECT 1335.480 1545.650 1335.740 1545.970 ;
        RECT 1335.480 1538.850 1335.740 1539.170 ;
        RECT 1335.540 1490.550 1335.680 1538.850 ;
        RECT 1335.480 1490.230 1335.740 1490.550 ;
        RECT 1335.020 1400.810 1335.280 1401.130 ;
        RECT 1335.080 1352.850 1335.220 1400.810 ;
        RECT 1335.020 1352.530 1335.280 1352.850 ;
        RECT 1335.480 1352.530 1335.740 1352.850 ;
        RECT 1335.540 1345.450 1335.680 1352.530 ;
        RECT 1335.080 1345.310 1335.680 1345.450 ;
        RECT 1335.080 1318.170 1335.220 1345.310 ;
        RECT 1335.020 1317.850 1335.280 1318.170 ;
        RECT 1335.020 1297.110 1335.280 1297.430 ;
        RECT 1335.080 1272.690 1335.220 1297.110 ;
        RECT 1334.160 1272.550 1335.220 1272.690 ;
        RECT 1334.160 1190.410 1334.300 1272.550 ;
        RECT 1334.160 1190.270 1335.680 1190.410 ;
        RECT 1335.540 1125.050 1335.680 1190.270 ;
        RECT 1335.480 1124.730 1335.740 1125.050 ;
        RECT 1335.480 1103.990 1335.740 1104.310 ;
        RECT 1335.540 1097.170 1335.680 1103.990 ;
        RECT 1335.480 1096.850 1335.740 1097.170 ;
        RECT 1335.020 1048.910 1335.280 1049.230 ;
        RECT 1335.080 1014.290 1335.220 1048.910 ;
        RECT 1335.080 1014.150 1335.680 1014.290 ;
        RECT 1335.540 1013.610 1335.680 1014.150 ;
        RECT 1335.080 1013.470 1335.680 1013.610 ;
        RECT 1335.080 966.270 1335.220 1013.470 ;
        RECT 1335.020 965.950 1335.280 966.270 ;
        RECT 1335.480 965.950 1335.740 966.270 ;
        RECT 1335.540 932.270 1335.680 965.950 ;
        RECT 1335.480 931.950 1335.740 932.270 ;
        RECT 1335.020 931.270 1335.280 931.590 ;
        RECT 1335.080 917.845 1335.220 931.270 ;
        RECT 1335.010 917.475 1335.290 917.845 ;
        RECT 1335.930 917.475 1336.210 917.845 ;
        RECT 1336.000 869.620 1336.140 917.475 ;
        RECT 1335.540 869.480 1336.140 869.620 ;
        RECT 1335.540 821.170 1335.680 869.480 ;
        RECT 1335.080 821.030 1335.680 821.170 ;
        RECT 1335.080 787.430 1335.220 821.030 ;
        RECT 1335.020 787.110 1335.280 787.430 ;
        RECT 1335.020 765.690 1335.280 766.010 ;
        RECT 1335.080 718.070 1335.220 765.690 ;
        RECT 1335.020 717.750 1335.280 718.070 ;
        RECT 1335.480 717.750 1335.740 718.070 ;
        RECT 1335.540 669.530 1335.680 717.750 ;
        RECT 1335.080 669.390 1335.680 669.530 ;
        RECT 1335.080 627.970 1335.220 669.390 ;
        RECT 1335.020 627.650 1335.280 627.970 ;
        RECT 1336.400 627.650 1336.660 627.970 ;
        RECT 1336.460 579.885 1336.600 627.650 ;
        RECT 1335.470 579.515 1335.750 579.885 ;
        RECT 1336.390 579.515 1336.670 579.885 ;
        RECT 1335.540 572.550 1335.680 579.515 ;
        RECT 1335.480 572.230 1335.740 572.550 ;
        RECT 1335.020 524.630 1335.280 524.950 ;
        RECT 1335.080 524.270 1335.220 524.630 ;
        RECT 1335.020 523.950 1335.280 524.270 ;
        RECT 1335.480 476.010 1335.740 476.330 ;
        RECT 1335.540 428.130 1335.680 476.010 ;
        RECT 1335.080 427.990 1335.680 428.130 ;
        RECT 1335.080 396.850 1335.220 427.990 ;
        RECT 1335.080 396.710 1335.680 396.850 ;
        RECT 1335.540 372.970 1335.680 396.710 ;
        RECT 1335.480 372.650 1335.740 372.970 ;
        RECT 1336.400 372.650 1336.660 372.970 ;
        RECT 1336.460 338.630 1336.600 372.650 ;
        RECT 1336.400 338.310 1336.660 338.630 ;
        RECT 1335.940 337.630 1336.200 337.950 ;
        RECT 1336.000 290.010 1336.140 337.630 ;
        RECT 1335.480 289.690 1335.740 290.010 ;
        RECT 1335.940 289.690 1336.200 290.010 ;
        RECT 1335.540 235.010 1335.680 289.690 ;
        RECT 1335.080 234.870 1335.680 235.010 ;
        RECT 1335.080 234.590 1335.220 234.870 ;
        RECT 1335.020 234.270 1335.280 234.590 ;
        RECT 1335.940 234.270 1336.200 234.590 ;
        RECT 1336.000 227.790 1336.140 234.270 ;
        RECT 1335.940 227.470 1336.200 227.790 ;
        RECT 1335.020 179.530 1335.280 179.850 ;
        RECT 1335.080 138.030 1335.220 179.530 ;
        RECT 1335.020 137.710 1335.280 138.030 ;
        RECT 1335.480 137.710 1335.740 138.030 ;
        RECT 1335.540 48.010 1335.680 137.710 ;
        RECT 1334.620 47.870 1335.680 48.010 ;
        RECT 1334.620 14.950 1334.760 47.870 ;
        RECT 1334.560 14.630 1334.820 14.950 ;
        RECT 537.840 13.950 538.100 14.270 ;
        RECT 537.900 2.400 538.040 13.950 ;
        RECT 537.690 -4.800 538.250 2.400 ;
      LAYER via2 ;
        RECT 1335.010 917.520 1335.290 917.800 ;
        RECT 1335.930 917.520 1336.210 917.800 ;
        RECT 1335.470 579.560 1335.750 579.840 ;
        RECT 1336.390 579.560 1336.670 579.840 ;
      LAYER met3 ;
        RECT 1334.985 917.810 1335.315 917.825 ;
        RECT 1335.905 917.810 1336.235 917.825 ;
        RECT 1334.985 917.510 1336.235 917.810 ;
        RECT 1334.985 917.495 1335.315 917.510 ;
        RECT 1335.905 917.495 1336.235 917.510 ;
        RECT 1335.445 579.850 1335.775 579.865 ;
        RECT 1336.365 579.850 1336.695 579.865 ;
        RECT 1335.445 579.550 1336.695 579.850 ;
        RECT 1335.445 579.535 1335.775 579.550 ;
        RECT 1336.365 579.535 1336.695 579.550 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 558.510 1685.280 558.830 1685.340 ;
        RECT 1434.350 1685.280 1434.670 1685.340 ;
        RECT 558.510 1685.140 1434.670 1685.280 ;
        RECT 558.510 1685.080 558.830 1685.140 ;
        RECT 1434.350 1685.080 1434.670 1685.140 ;
        RECT 555.750 15.540 556.070 15.600 ;
        RECT 558.510 15.540 558.830 15.600 ;
        RECT 555.750 15.400 558.830 15.540 ;
        RECT 555.750 15.340 556.070 15.400 ;
        RECT 558.510 15.340 558.830 15.400 ;
      LAYER via ;
        RECT 558.540 1685.080 558.800 1685.340 ;
        RECT 1434.380 1685.080 1434.640 1685.340 ;
        RECT 555.780 15.340 556.040 15.600 ;
        RECT 558.540 15.340 558.800 15.600 ;
      LAYER met2 ;
        RECT 1434.300 1700.000 1434.580 1702.400 ;
        RECT 1434.440 1685.370 1434.580 1700.000 ;
        RECT 558.540 1685.050 558.800 1685.370 ;
        RECT 1434.380 1685.050 1434.640 1685.370 ;
        RECT 558.600 15.630 558.740 1685.050 ;
        RECT 555.780 15.310 556.040 15.630 ;
        RECT 558.540 15.310 558.800 15.630 ;
        RECT 555.840 2.400 555.980 15.310 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 607.345 14.365 608.435 14.535 ;
      LAYER mcon ;
        RECT 608.265 14.365 608.435 14.535 ;
      LAYER met1 ;
        RECT 1341.890 1689.360 1342.210 1689.420 ;
        RECT 1443.550 1689.360 1443.870 1689.420 ;
        RECT 1341.890 1689.220 1443.870 1689.360 ;
        RECT 1341.890 1689.160 1342.210 1689.220 ;
        RECT 1443.550 1689.160 1443.870 1689.220 ;
        RECT 573.690 14.520 574.010 14.580 ;
        RECT 607.285 14.520 607.575 14.565 ;
        RECT 573.690 14.380 607.575 14.520 ;
        RECT 573.690 14.320 574.010 14.380 ;
        RECT 607.285 14.335 607.575 14.380 ;
        RECT 608.205 14.520 608.495 14.565 ;
        RECT 1341.890 14.520 1342.210 14.580 ;
        RECT 608.205 14.380 1342.210 14.520 ;
        RECT 608.205 14.335 608.495 14.380 ;
        RECT 1341.890 14.320 1342.210 14.380 ;
      LAYER via ;
        RECT 1341.920 1689.160 1342.180 1689.420 ;
        RECT 1443.580 1689.160 1443.840 1689.420 ;
        RECT 573.720 14.320 573.980 14.580 ;
        RECT 1341.920 14.320 1342.180 14.580 ;
      LAYER met2 ;
        RECT 1443.500 1700.000 1443.780 1702.400 ;
        RECT 1443.640 1689.450 1443.780 1700.000 ;
        RECT 1341.920 1689.130 1342.180 1689.450 ;
        RECT 1443.580 1689.130 1443.840 1689.450 ;
        RECT 1341.980 14.610 1342.120 1689.130 ;
        RECT 573.720 14.290 573.980 14.610 ;
        RECT 1341.920 14.290 1342.180 14.610 ;
        RECT 573.780 2.400 573.920 14.290 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 1684.940 593.330 1685.000 ;
        RECT 1452.750 1684.940 1453.070 1685.000 ;
        RECT 593.010 1684.800 1453.070 1684.940 ;
        RECT 593.010 1684.740 593.330 1684.800 ;
        RECT 1452.750 1684.740 1453.070 1684.800 ;
      LAYER via ;
        RECT 593.040 1684.740 593.300 1685.000 ;
        RECT 1452.780 1684.740 1453.040 1685.000 ;
      LAYER met2 ;
        RECT 1452.700 1700.000 1452.980 1702.400 ;
        RECT 1452.840 1685.030 1452.980 1700.000 ;
        RECT 593.040 1684.710 593.300 1685.030 ;
        RECT 1452.780 1684.710 1453.040 1685.030 ;
        RECT 593.100 16.730 593.240 1684.710 ;
        RECT 591.260 16.590 593.240 16.730 ;
        RECT 591.260 2.400 591.400 16.590 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 120.590 1687.320 120.910 1687.380 ;
        RECT 120.590 1687.180 1186.180 1687.320 ;
        RECT 120.590 1687.120 120.910 1687.180 ;
        RECT 1186.040 1686.980 1186.180 1687.180 ;
        RECT 1198.830 1686.980 1199.150 1687.040 ;
        RECT 1186.040 1686.840 1199.150 1686.980 ;
        RECT 1198.830 1686.780 1199.150 1686.840 ;
        RECT 97.590 17.920 97.910 17.980 ;
        RECT 120.590 17.920 120.910 17.980 ;
        RECT 97.590 17.780 120.910 17.920 ;
        RECT 97.590 17.720 97.910 17.780 ;
        RECT 120.590 17.720 120.910 17.780 ;
      LAYER via ;
        RECT 120.620 1687.120 120.880 1687.380 ;
        RECT 1198.860 1686.780 1199.120 1687.040 ;
        RECT 97.620 17.720 97.880 17.980 ;
        RECT 120.620 17.720 120.880 17.980 ;
      LAYER met2 ;
        RECT 1198.780 1700.000 1199.060 1702.400 ;
        RECT 120.620 1687.090 120.880 1687.410 ;
        RECT 120.680 18.010 120.820 1687.090 ;
        RECT 1198.920 1687.070 1199.060 1700.000 ;
        RECT 1198.860 1686.750 1199.120 1687.070 ;
        RECT 97.620 17.690 97.880 18.010 ;
        RECT 120.620 17.690 120.880 18.010 ;
        RECT 97.680 2.400 97.820 17.690 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1348.790 1689.020 1349.110 1689.080 ;
        RECT 1461.950 1689.020 1462.270 1689.080 ;
        RECT 1348.790 1688.880 1462.270 1689.020 ;
        RECT 1348.790 1688.820 1349.110 1688.880 ;
        RECT 1461.950 1688.820 1462.270 1688.880 ;
        RECT 609.110 14.180 609.430 14.240 ;
        RECT 1348.790 14.180 1349.110 14.240 ;
        RECT 609.110 14.040 1349.110 14.180 ;
        RECT 609.110 13.980 609.430 14.040 ;
        RECT 1348.790 13.980 1349.110 14.040 ;
      LAYER via ;
        RECT 1348.820 1688.820 1349.080 1689.080 ;
        RECT 1461.980 1688.820 1462.240 1689.080 ;
        RECT 609.140 13.980 609.400 14.240 ;
        RECT 1348.820 13.980 1349.080 14.240 ;
      LAYER met2 ;
        RECT 1461.900 1700.000 1462.180 1702.400 ;
        RECT 1462.040 1689.110 1462.180 1700.000 ;
        RECT 1348.820 1688.790 1349.080 1689.110 ;
        RECT 1461.980 1688.790 1462.240 1689.110 ;
        RECT 1348.880 14.270 1349.020 1688.790 ;
        RECT 609.140 13.950 609.400 14.270 ;
        RECT 1348.820 13.950 1349.080 14.270 ;
        RECT 609.200 2.400 609.340 13.950 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 1684.600 627.830 1684.660 ;
        RECT 1471.150 1684.600 1471.470 1684.660 ;
        RECT 627.510 1684.460 1471.470 1684.600 ;
        RECT 627.510 1684.400 627.830 1684.460 ;
        RECT 1471.150 1684.400 1471.470 1684.460 ;
      LAYER via ;
        RECT 627.540 1684.400 627.800 1684.660 ;
        RECT 1471.180 1684.400 1471.440 1684.660 ;
      LAYER met2 ;
        RECT 1471.100 1700.000 1471.380 1702.400 ;
        RECT 1471.240 1684.690 1471.380 1700.000 ;
        RECT 627.540 1684.370 627.800 1684.690 ;
        RECT 1471.180 1684.370 1471.440 1684.690 ;
        RECT 627.600 17.410 627.740 1684.370 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1207.570 1678.140 1207.890 1678.200 ;
        RECT 1209.870 1678.140 1210.190 1678.200 ;
        RECT 1207.570 1678.000 1210.190 1678.140 ;
        RECT 1207.570 1677.940 1207.890 1678.000 ;
        RECT 1209.870 1677.940 1210.190 1678.000 ;
        RECT 121.510 17.920 121.830 17.980 ;
        RECT 1207.570 17.920 1207.890 17.980 ;
        RECT 121.510 17.780 1207.890 17.920 ;
        RECT 121.510 17.720 121.830 17.780 ;
        RECT 1207.570 17.720 1207.890 17.780 ;
      LAYER via ;
        RECT 1207.600 1677.940 1207.860 1678.200 ;
        RECT 1209.900 1677.940 1210.160 1678.200 ;
        RECT 121.540 17.720 121.800 17.980 ;
        RECT 1207.600 17.720 1207.860 17.980 ;
      LAYER met2 ;
        RECT 1211.200 1700.410 1211.480 1702.400 ;
        RECT 1209.960 1700.270 1211.480 1700.410 ;
        RECT 1209.960 1678.230 1210.100 1700.270 ;
        RECT 1211.200 1700.000 1211.480 1700.270 ;
        RECT 1207.600 1677.910 1207.860 1678.230 ;
        RECT 1209.900 1677.910 1210.160 1678.230 ;
        RECT 1207.660 18.010 1207.800 1677.910 ;
        RECT 121.540 17.690 121.800 18.010 ;
        RECT 1207.600 17.690 1207.860 18.010 ;
        RECT 121.600 2.400 121.740 17.690 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1197.065 1687.505 1197.235 1688.355 ;
      LAYER mcon ;
        RECT 1197.065 1688.185 1197.235 1688.355 ;
      LAYER met1 ;
        RECT 161.990 1688.340 162.310 1688.400 ;
        RECT 1197.005 1688.340 1197.295 1688.385 ;
        RECT 161.990 1688.200 1197.295 1688.340 ;
        RECT 161.990 1688.140 162.310 1688.200 ;
        RECT 1197.005 1688.155 1197.295 1688.200 ;
        RECT 1197.005 1687.660 1197.295 1687.705 ;
        RECT 1223.210 1687.660 1223.530 1687.720 ;
        RECT 1197.005 1687.520 1223.530 1687.660 ;
        RECT 1197.005 1687.475 1197.295 1687.520 ;
        RECT 1223.210 1687.460 1223.530 1687.520 ;
        RECT 145.430 15.880 145.750 15.940 ;
        RECT 161.990 15.880 162.310 15.940 ;
        RECT 145.430 15.740 162.310 15.880 ;
        RECT 145.430 15.680 145.750 15.740 ;
        RECT 161.990 15.680 162.310 15.740 ;
      LAYER via ;
        RECT 162.020 1688.140 162.280 1688.400 ;
        RECT 1223.240 1687.460 1223.500 1687.720 ;
        RECT 145.460 15.680 145.720 15.940 ;
        RECT 162.020 15.680 162.280 15.940 ;
      LAYER met2 ;
        RECT 1223.160 1700.000 1223.440 1702.400 ;
        RECT 162.020 1688.110 162.280 1688.430 ;
        RECT 162.080 15.970 162.220 1688.110 ;
        RECT 1223.300 1687.750 1223.440 1700.000 ;
        RECT 1223.240 1687.430 1223.500 1687.750 ;
        RECT 145.460 15.650 145.720 15.970 ;
        RECT 162.020 15.650 162.280 15.970 ;
        RECT 145.520 2.400 145.660 15.650 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1228.270 1677.800 1228.590 1677.860 ;
        RECT 1232.410 1677.800 1232.730 1677.860 ;
        RECT 1228.270 1677.660 1232.730 1677.800 ;
        RECT 1228.270 1677.600 1228.590 1677.660 ;
        RECT 1232.410 1677.600 1232.730 1677.660 ;
        RECT 163.370 18.600 163.690 18.660 ;
        RECT 1228.270 18.600 1228.590 18.660 ;
        RECT 163.370 18.460 1228.590 18.600 ;
        RECT 163.370 18.400 163.690 18.460 ;
        RECT 1228.270 18.400 1228.590 18.460 ;
      LAYER via ;
        RECT 1228.300 1677.600 1228.560 1677.860 ;
        RECT 1232.440 1677.600 1232.700 1677.860 ;
        RECT 163.400 18.400 163.660 18.660 ;
        RECT 1228.300 18.400 1228.560 18.660 ;
      LAYER met2 ;
        RECT 1232.360 1700.000 1232.640 1702.400 ;
        RECT 1232.500 1677.890 1232.640 1700.000 ;
        RECT 1228.300 1677.570 1228.560 1677.890 ;
        RECT 1232.440 1677.570 1232.700 1677.890 ;
        RECT 1228.360 18.690 1228.500 1677.570 ;
        RECT 163.400 18.370 163.660 18.690 ;
        RECT 1228.300 18.370 1228.560 18.690 ;
        RECT 163.460 2.400 163.600 18.370 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1173.145 1688.525 1175.155 1688.695 ;
        RECT 1174.985 1687.505 1175.155 1688.525 ;
      LAYER met1 ;
        RECT 196.490 1688.680 196.810 1688.740 ;
        RECT 1173.085 1688.680 1173.375 1688.725 ;
        RECT 196.490 1688.540 1173.375 1688.680 ;
        RECT 196.490 1688.480 196.810 1688.540 ;
        RECT 1173.085 1688.495 1173.375 1688.540 ;
        RECT 1241.610 1688.000 1241.930 1688.060 ;
        RECT 1187.880 1687.860 1241.930 1688.000 ;
        RECT 1174.925 1687.660 1175.215 1687.705 ;
        RECT 1187.880 1687.660 1188.020 1687.860 ;
        RECT 1241.610 1687.800 1241.930 1687.860 ;
        RECT 1174.925 1687.520 1188.020 1687.660 ;
        RECT 1174.925 1687.475 1175.215 1687.520 ;
        RECT 180.850 16.900 181.170 16.960 ;
        RECT 196.490 16.900 196.810 16.960 ;
        RECT 180.850 16.760 196.810 16.900 ;
        RECT 180.850 16.700 181.170 16.760 ;
        RECT 196.490 16.700 196.810 16.760 ;
      LAYER via ;
        RECT 196.520 1688.480 196.780 1688.740 ;
        RECT 1241.640 1687.800 1241.900 1688.060 ;
        RECT 180.880 16.700 181.140 16.960 ;
        RECT 196.520 16.700 196.780 16.960 ;
      LAYER met2 ;
        RECT 1241.560 1700.000 1241.840 1702.400 ;
        RECT 196.520 1688.450 196.780 1688.770 ;
        RECT 196.580 16.990 196.720 1688.450 ;
        RECT 1241.700 1688.090 1241.840 1700.000 ;
        RECT 1241.640 1687.770 1241.900 1688.090 ;
        RECT 180.880 16.670 181.140 16.990 ;
        RECT 196.520 16.670 196.780 16.990 ;
        RECT 180.940 2.400 181.080 16.670 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 198.790 19.280 199.110 19.340 ;
        RECT 1248.970 19.280 1249.290 19.340 ;
        RECT 198.790 19.140 1249.290 19.280 ;
        RECT 198.790 19.080 199.110 19.140 ;
        RECT 1248.970 19.080 1249.290 19.140 ;
      LAYER via ;
        RECT 198.820 19.080 199.080 19.340 ;
        RECT 1249.000 19.080 1249.260 19.340 ;
      LAYER met2 ;
        RECT 1250.760 1700.410 1251.040 1702.400 ;
        RECT 1249.060 1700.270 1251.040 1700.410 ;
        RECT 1249.060 19.370 1249.200 1700.270 ;
        RECT 1250.760 1700.000 1251.040 1700.270 ;
        RECT 198.820 19.050 199.080 19.370 ;
        RECT 1249.000 19.050 1249.260 19.370 ;
        RECT 198.880 2.400 199.020 19.050 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 306.890 1686.640 307.210 1686.700 ;
        RECT 1260.010 1686.640 1260.330 1686.700 ;
        RECT 306.890 1686.500 1260.330 1686.640 ;
        RECT 306.890 1686.440 307.210 1686.500 ;
        RECT 1260.010 1686.440 1260.330 1686.500 ;
        RECT 251.780 16.760 291.480 16.900 ;
        RECT 216.730 16.220 217.050 16.280 ;
        RECT 251.780 16.220 251.920 16.760 ;
        RECT 291.340 16.560 291.480 16.760 ;
        RECT 306.890 16.560 307.210 16.620 ;
        RECT 291.340 16.420 307.210 16.560 ;
        RECT 306.890 16.360 307.210 16.420 ;
        RECT 216.730 16.080 251.920 16.220 ;
        RECT 216.730 16.020 217.050 16.080 ;
      LAYER via ;
        RECT 306.920 1686.440 307.180 1686.700 ;
        RECT 1260.040 1686.440 1260.300 1686.700 ;
        RECT 216.760 16.020 217.020 16.280 ;
        RECT 306.920 16.360 307.180 16.620 ;
      LAYER met2 ;
        RECT 1259.960 1700.000 1260.240 1702.400 ;
        RECT 1260.100 1686.730 1260.240 1700.000 ;
        RECT 306.920 1686.410 307.180 1686.730 ;
        RECT 1260.040 1686.410 1260.300 1686.730 ;
        RECT 306.980 16.650 307.120 1686.410 ;
        RECT 306.920 16.330 307.180 16.650 ;
        RECT 216.760 15.990 217.020 16.310 ;
        RECT 216.820 2.400 216.960 15.990 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1263.765 1304.325 1263.935 1352.435 ;
        RECT 1263.765 1207.425 1263.935 1255.875 ;
        RECT 1264.225 862.665 1264.395 910.775 ;
        RECT 1263.765 483.225 1263.935 530.995 ;
        RECT 1263.765 386.325 1263.935 434.435 ;
        RECT 1263.765 144.925 1263.935 186.915 ;
        RECT 1264.225 89.845 1264.395 137.955 ;
      LAYER mcon ;
        RECT 1263.765 1352.265 1263.935 1352.435 ;
        RECT 1263.765 1255.705 1263.935 1255.875 ;
        RECT 1264.225 910.605 1264.395 910.775 ;
        RECT 1263.765 530.825 1263.935 530.995 ;
        RECT 1263.765 434.265 1263.935 434.435 ;
        RECT 1263.765 186.745 1263.935 186.915 ;
        RECT 1264.225 137.785 1264.395 137.955 ;
      LAYER met1 ;
        RECT 1262.770 1681.540 1263.090 1681.600 ;
        RECT 1269.210 1681.540 1269.530 1681.600 ;
        RECT 1262.770 1681.400 1269.530 1681.540 ;
        RECT 1262.770 1681.340 1263.090 1681.400 ;
        RECT 1269.210 1681.340 1269.530 1681.400 ;
        RECT 1262.770 1545.880 1263.090 1545.940 ;
        RECT 1263.690 1545.880 1264.010 1545.940 ;
        RECT 1262.770 1545.740 1264.010 1545.880 ;
        RECT 1262.770 1545.680 1263.090 1545.740 ;
        RECT 1263.690 1545.680 1264.010 1545.740 ;
        RECT 1263.690 1352.420 1264.010 1352.480 ;
        RECT 1263.495 1352.280 1264.010 1352.420 ;
        RECT 1263.690 1352.220 1264.010 1352.280 ;
        RECT 1263.690 1304.480 1264.010 1304.540 ;
        RECT 1263.495 1304.340 1264.010 1304.480 ;
        RECT 1263.690 1304.280 1264.010 1304.340 ;
        RECT 1263.690 1255.860 1264.010 1255.920 ;
        RECT 1263.495 1255.720 1264.010 1255.860 ;
        RECT 1263.690 1255.660 1264.010 1255.720 ;
        RECT 1263.690 1207.580 1264.010 1207.640 ;
        RECT 1263.495 1207.440 1264.010 1207.580 ;
        RECT 1263.690 1207.380 1264.010 1207.440 ;
        RECT 1263.690 1111.020 1264.010 1111.080 ;
        RECT 1264.610 1111.020 1264.930 1111.080 ;
        RECT 1263.690 1110.880 1264.930 1111.020 ;
        RECT 1263.690 1110.820 1264.010 1110.880 ;
        RECT 1264.610 1110.820 1264.930 1110.880 ;
        RECT 1263.690 1062.740 1264.010 1062.800 ;
        RECT 1264.150 1062.740 1264.470 1062.800 ;
        RECT 1263.690 1062.600 1264.470 1062.740 ;
        RECT 1263.690 1062.540 1264.010 1062.600 ;
        RECT 1264.150 1062.540 1264.470 1062.600 ;
        RECT 1262.310 1014.460 1262.630 1014.520 ;
        RECT 1262.770 1014.460 1263.090 1014.520 ;
        RECT 1262.310 1014.320 1263.090 1014.460 ;
        RECT 1262.310 1014.260 1262.630 1014.320 ;
        RECT 1262.770 1014.260 1263.090 1014.320 ;
        RECT 1262.770 966.180 1263.090 966.240 ;
        RECT 1263.690 966.180 1264.010 966.240 ;
        RECT 1262.770 966.040 1264.010 966.180 ;
        RECT 1262.770 965.980 1263.090 966.040 ;
        RECT 1263.690 965.980 1264.010 966.040 ;
        RECT 1263.690 917.700 1264.010 917.960 ;
        RECT 1263.780 917.220 1263.920 917.700 ;
        RECT 1264.150 917.220 1264.470 917.280 ;
        RECT 1263.780 917.080 1264.470 917.220 ;
        RECT 1264.150 917.020 1264.470 917.080 ;
        RECT 1264.150 910.760 1264.470 910.820 ;
        RECT 1263.955 910.620 1264.470 910.760 ;
        RECT 1264.150 910.560 1264.470 910.620 ;
        RECT 1264.150 862.820 1264.470 862.880 ;
        RECT 1263.955 862.680 1264.470 862.820 ;
        RECT 1264.150 862.620 1264.470 862.680 ;
        RECT 1262.770 821.000 1263.090 821.060 ;
        RECT 1264.150 821.000 1264.470 821.060 ;
        RECT 1262.770 820.860 1264.470 821.000 ;
        RECT 1262.770 820.800 1263.090 820.860 ;
        RECT 1264.150 820.800 1264.470 820.860 ;
        RECT 1262.770 727.840 1263.090 727.900 ;
        RECT 1263.690 727.840 1264.010 727.900 ;
        RECT 1262.770 727.700 1264.010 727.840 ;
        RECT 1262.770 727.640 1263.090 727.700 ;
        RECT 1263.690 727.640 1264.010 727.700 ;
        RECT 1263.690 627.880 1264.010 627.940 ;
        RECT 1264.610 627.880 1264.930 627.940 ;
        RECT 1263.690 627.740 1264.930 627.880 ;
        RECT 1263.690 627.680 1264.010 627.740 ;
        RECT 1264.610 627.680 1264.930 627.740 ;
        RECT 1263.690 530.980 1264.010 531.040 ;
        RECT 1263.495 530.840 1264.010 530.980 ;
        RECT 1263.690 530.780 1264.010 530.840 ;
        RECT 1263.690 483.380 1264.010 483.440 ;
        RECT 1263.495 483.240 1264.010 483.380 ;
        RECT 1263.690 483.180 1264.010 483.240 ;
        RECT 1263.690 434.420 1264.010 434.480 ;
        RECT 1263.495 434.280 1264.010 434.420 ;
        RECT 1263.690 434.220 1264.010 434.280 ;
        RECT 1263.690 386.480 1264.010 386.540 ;
        RECT 1263.495 386.340 1264.010 386.480 ;
        RECT 1263.690 386.280 1264.010 386.340 ;
        RECT 1263.690 186.900 1264.010 186.960 ;
        RECT 1263.495 186.760 1264.010 186.900 ;
        RECT 1263.690 186.700 1264.010 186.760 ;
        RECT 1263.705 145.080 1263.995 145.125 ;
        RECT 1264.150 145.080 1264.470 145.140 ;
        RECT 1263.705 144.940 1264.470 145.080 ;
        RECT 1263.705 144.895 1263.995 144.940 ;
        RECT 1264.150 144.880 1264.470 144.940 ;
        RECT 1264.150 137.940 1264.470 138.000 ;
        RECT 1263.955 137.800 1264.470 137.940 ;
        RECT 1264.150 137.740 1264.470 137.800 ;
        RECT 1264.150 90.000 1264.470 90.060 ;
        RECT 1263.955 89.860 1264.470 90.000 ;
        RECT 1264.150 89.800 1264.470 89.860 ;
        RECT 234.670 19.960 234.990 20.020 ;
        RECT 1263.690 19.960 1264.010 20.020 ;
        RECT 234.670 19.820 1264.010 19.960 ;
        RECT 234.670 19.760 234.990 19.820 ;
        RECT 1263.690 19.760 1264.010 19.820 ;
      LAYER via ;
        RECT 1262.800 1681.340 1263.060 1681.600 ;
        RECT 1269.240 1681.340 1269.500 1681.600 ;
        RECT 1262.800 1545.680 1263.060 1545.940 ;
        RECT 1263.720 1545.680 1263.980 1545.940 ;
        RECT 1263.720 1352.220 1263.980 1352.480 ;
        RECT 1263.720 1304.280 1263.980 1304.540 ;
        RECT 1263.720 1255.660 1263.980 1255.920 ;
        RECT 1263.720 1207.380 1263.980 1207.640 ;
        RECT 1263.720 1110.820 1263.980 1111.080 ;
        RECT 1264.640 1110.820 1264.900 1111.080 ;
        RECT 1263.720 1062.540 1263.980 1062.800 ;
        RECT 1264.180 1062.540 1264.440 1062.800 ;
        RECT 1262.340 1014.260 1262.600 1014.520 ;
        RECT 1262.800 1014.260 1263.060 1014.520 ;
        RECT 1262.800 965.980 1263.060 966.240 ;
        RECT 1263.720 965.980 1263.980 966.240 ;
        RECT 1263.720 917.700 1263.980 917.960 ;
        RECT 1264.180 917.020 1264.440 917.280 ;
        RECT 1264.180 910.560 1264.440 910.820 ;
        RECT 1264.180 862.620 1264.440 862.880 ;
        RECT 1262.800 820.800 1263.060 821.060 ;
        RECT 1264.180 820.800 1264.440 821.060 ;
        RECT 1262.800 727.640 1263.060 727.900 ;
        RECT 1263.720 727.640 1263.980 727.900 ;
        RECT 1263.720 627.680 1263.980 627.940 ;
        RECT 1264.640 627.680 1264.900 627.940 ;
        RECT 1263.720 530.780 1263.980 531.040 ;
        RECT 1263.720 483.180 1263.980 483.440 ;
        RECT 1263.720 434.220 1263.980 434.480 ;
        RECT 1263.720 386.280 1263.980 386.540 ;
        RECT 1263.720 186.700 1263.980 186.960 ;
        RECT 1264.180 144.880 1264.440 145.140 ;
        RECT 1264.180 137.740 1264.440 138.000 ;
        RECT 1264.180 89.800 1264.440 90.060 ;
        RECT 234.700 19.760 234.960 20.020 ;
        RECT 1263.720 19.760 1263.980 20.020 ;
      LAYER met2 ;
        RECT 1269.160 1700.000 1269.440 1702.400 ;
        RECT 1269.300 1681.630 1269.440 1700.000 ;
        RECT 1262.800 1681.310 1263.060 1681.630 ;
        RECT 1269.240 1681.310 1269.500 1681.630 ;
        RECT 1262.860 1545.970 1263.000 1681.310 ;
        RECT 1262.800 1545.650 1263.060 1545.970 ;
        RECT 1263.720 1545.650 1263.980 1545.970 ;
        RECT 1263.780 1352.510 1263.920 1545.650 ;
        RECT 1263.720 1352.190 1263.980 1352.510 ;
        RECT 1263.720 1304.250 1263.980 1304.570 ;
        RECT 1263.780 1255.950 1263.920 1304.250 ;
        RECT 1263.720 1255.630 1263.980 1255.950 ;
        RECT 1263.780 1207.670 1263.920 1207.825 ;
        RECT 1263.720 1207.410 1263.980 1207.670 ;
        RECT 1263.720 1207.350 1264.380 1207.410 ;
        RECT 1263.780 1207.270 1264.380 1207.350 ;
        RECT 1264.240 1159.810 1264.380 1207.270 ;
        RECT 1263.780 1159.670 1264.380 1159.810 ;
        RECT 1263.780 1159.245 1263.920 1159.670 ;
        RECT 1263.710 1158.875 1263.990 1159.245 ;
        RECT 1264.630 1158.875 1264.910 1159.245 ;
        RECT 1263.780 1111.110 1263.920 1111.265 ;
        RECT 1264.700 1111.110 1264.840 1158.875 ;
        RECT 1263.720 1110.850 1263.980 1111.110 ;
        RECT 1263.720 1110.790 1264.380 1110.850 ;
        RECT 1264.640 1110.790 1264.900 1111.110 ;
        RECT 1263.780 1110.710 1264.380 1110.790 ;
        RECT 1264.240 1062.830 1264.380 1110.710 ;
        RECT 1263.720 1062.685 1263.980 1062.830 ;
        RECT 1262.330 1062.315 1262.610 1062.685 ;
        RECT 1263.710 1062.315 1263.990 1062.685 ;
        RECT 1264.180 1062.510 1264.440 1062.830 ;
        RECT 1262.400 1014.550 1262.540 1062.315 ;
        RECT 1262.340 1014.230 1262.600 1014.550 ;
        RECT 1262.800 1014.230 1263.060 1014.550 ;
        RECT 1262.860 966.270 1263.000 1014.230 ;
        RECT 1262.800 965.950 1263.060 966.270 ;
        RECT 1263.720 965.950 1263.980 966.270 ;
        RECT 1263.780 917.990 1263.920 965.950 ;
        RECT 1263.720 917.670 1263.980 917.990 ;
        RECT 1264.180 916.990 1264.440 917.310 ;
        RECT 1264.240 910.850 1264.380 916.990 ;
        RECT 1264.180 910.530 1264.440 910.850 ;
        RECT 1264.180 862.590 1264.440 862.910 ;
        RECT 1264.240 821.090 1264.380 862.590 ;
        RECT 1262.800 820.770 1263.060 821.090 ;
        RECT 1264.180 820.770 1264.440 821.090 ;
        RECT 1262.860 773.005 1263.000 820.770 ;
        RECT 1262.790 772.635 1263.070 773.005 ;
        RECT 1263.710 772.635 1263.990 773.005 ;
        RECT 1263.780 727.930 1263.920 772.635 ;
        RECT 1262.800 727.610 1263.060 727.930 ;
        RECT 1263.720 727.610 1263.980 727.930 ;
        RECT 1262.860 676.445 1263.000 727.610 ;
        RECT 1262.790 676.075 1263.070 676.445 ;
        RECT 1263.710 676.075 1263.990 676.445 ;
        RECT 1263.780 627.970 1263.920 676.075 ;
        RECT 1263.720 627.650 1263.980 627.970 ;
        RECT 1264.640 627.650 1264.900 627.970 ;
        RECT 1264.700 579.885 1264.840 627.650 ;
        RECT 1263.710 579.515 1263.990 579.885 ;
        RECT 1264.630 579.515 1264.910 579.885 ;
        RECT 1263.780 531.070 1263.920 579.515 ;
        RECT 1263.720 530.750 1263.980 531.070 ;
        RECT 1263.720 483.150 1263.980 483.470 ;
        RECT 1263.780 434.510 1263.920 483.150 ;
        RECT 1263.720 434.190 1263.980 434.510 ;
        RECT 1263.720 386.250 1263.980 386.570 ;
        RECT 1263.780 186.990 1263.920 386.250 ;
        RECT 1263.720 186.670 1263.980 186.990 ;
        RECT 1264.180 144.850 1264.440 145.170 ;
        RECT 1264.240 138.030 1264.380 144.850 ;
        RECT 1264.180 137.710 1264.440 138.030 ;
        RECT 1264.180 89.770 1264.440 90.090 ;
        RECT 1264.240 62.290 1264.380 89.770 ;
        RECT 1263.780 62.150 1264.380 62.290 ;
        RECT 1263.780 20.050 1263.920 62.150 ;
        RECT 234.700 19.730 234.960 20.050 ;
        RECT 1263.720 19.730 1263.980 20.050 ;
        RECT 234.760 2.400 234.900 19.730 ;
        RECT 234.550 -4.800 235.110 2.400 ;
      LAYER via2 ;
        RECT 1263.710 1158.920 1263.990 1159.200 ;
        RECT 1264.630 1158.920 1264.910 1159.200 ;
        RECT 1262.330 1062.360 1262.610 1062.640 ;
        RECT 1263.710 1062.360 1263.990 1062.640 ;
        RECT 1262.790 772.680 1263.070 772.960 ;
        RECT 1263.710 772.680 1263.990 772.960 ;
        RECT 1262.790 676.120 1263.070 676.400 ;
        RECT 1263.710 676.120 1263.990 676.400 ;
        RECT 1263.710 579.560 1263.990 579.840 ;
        RECT 1264.630 579.560 1264.910 579.840 ;
      LAYER met3 ;
        RECT 1263.685 1159.210 1264.015 1159.225 ;
        RECT 1264.605 1159.210 1264.935 1159.225 ;
        RECT 1263.685 1158.910 1264.935 1159.210 ;
        RECT 1263.685 1158.895 1264.015 1158.910 ;
        RECT 1264.605 1158.895 1264.935 1158.910 ;
        RECT 1262.305 1062.650 1262.635 1062.665 ;
        RECT 1263.685 1062.650 1264.015 1062.665 ;
        RECT 1262.305 1062.350 1264.015 1062.650 ;
        RECT 1262.305 1062.335 1262.635 1062.350 ;
        RECT 1263.685 1062.335 1264.015 1062.350 ;
        RECT 1262.765 772.970 1263.095 772.985 ;
        RECT 1263.685 772.970 1264.015 772.985 ;
        RECT 1262.765 772.670 1264.015 772.970 ;
        RECT 1262.765 772.655 1263.095 772.670 ;
        RECT 1263.685 772.655 1264.015 772.670 ;
        RECT 1262.765 676.410 1263.095 676.425 ;
        RECT 1263.685 676.410 1264.015 676.425 ;
        RECT 1262.765 676.110 1264.015 676.410 ;
        RECT 1262.765 676.095 1263.095 676.110 ;
        RECT 1263.685 676.095 1264.015 676.110 ;
        RECT 1263.685 579.850 1264.015 579.865 ;
        RECT 1264.605 579.850 1264.935 579.865 ;
        RECT 1263.685 579.550 1264.935 579.850 ;
        RECT 1263.685 579.535 1264.015 579.550 ;
        RECT 1264.605 579.535 1264.935 579.550 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1140.485 1686.995 1140.655 1687.675 ;
        RECT 1140.485 1686.825 1141.575 1686.995 ;
      LAYER mcon ;
        RECT 1140.485 1687.505 1140.655 1687.675 ;
        RECT 1141.405 1686.825 1141.575 1686.995 ;
      LAYER met1 ;
        RECT 86.090 1687.660 86.410 1687.720 ;
        RECT 1140.425 1687.660 1140.715 1687.705 ;
        RECT 86.090 1687.520 1140.715 1687.660 ;
        RECT 86.090 1687.460 86.410 1687.520 ;
        RECT 1140.425 1687.475 1140.715 1687.520 ;
        RECT 1141.345 1686.980 1141.635 1687.025 ;
        RECT 1177.210 1686.980 1177.530 1687.040 ;
        RECT 1141.345 1686.840 1177.530 1686.980 ;
        RECT 1141.345 1686.795 1141.635 1686.840 ;
        RECT 1177.210 1686.780 1177.530 1686.840 ;
        RECT 56.190 16.560 56.510 16.620 ;
        RECT 86.090 16.560 86.410 16.620 ;
        RECT 56.190 16.420 86.410 16.560 ;
        RECT 56.190 16.360 56.510 16.420 ;
        RECT 86.090 16.360 86.410 16.420 ;
      LAYER via ;
        RECT 86.120 1687.460 86.380 1687.720 ;
        RECT 1177.240 1686.780 1177.500 1687.040 ;
        RECT 56.220 16.360 56.480 16.620 ;
        RECT 86.120 16.360 86.380 16.620 ;
      LAYER met2 ;
        RECT 1177.160 1700.000 1177.440 1702.400 ;
        RECT 86.120 1687.430 86.380 1687.750 ;
        RECT 86.180 16.650 86.320 1687.430 ;
        RECT 1177.300 1687.070 1177.440 1700.000 ;
        RECT 1177.240 1686.750 1177.500 1687.070 ;
        RECT 56.220 16.330 56.480 16.650 ;
        RECT 86.120 16.330 86.380 16.650 ;
        RECT 56.280 2.400 56.420 16.330 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 80.110 17.240 80.430 17.300 ;
        RECT 1187.790 17.240 1188.110 17.300 ;
        RECT 80.110 17.100 1188.110 17.240 ;
        RECT 80.110 17.040 80.430 17.100 ;
        RECT 1187.790 17.040 1188.110 17.100 ;
      LAYER via ;
        RECT 80.140 17.040 80.400 17.300 ;
        RECT 1187.820 17.040 1188.080 17.300 ;
      LAYER met2 ;
        RECT 1189.580 1700.410 1189.860 1702.400 ;
        RECT 1187.880 1700.270 1189.860 1700.410 ;
        RECT 1187.880 17.330 1188.020 1700.270 ;
        RECT 1189.580 1700.000 1189.860 1700.270 ;
        RECT 80.140 17.010 80.400 17.330 ;
        RECT 1187.820 17.010 1188.080 17.330 ;
        RECT 80.200 2.400 80.340 17.010 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1187.405 1687.845 1187.575 1688.695 ;
      LAYER mcon ;
        RECT 1187.405 1688.525 1187.575 1688.695 ;
      LAYER met1 ;
        RECT 1187.345 1688.680 1187.635 1688.725 ;
        RECT 1202.050 1688.680 1202.370 1688.740 ;
        RECT 1187.345 1688.540 1202.370 1688.680 ;
        RECT 1187.345 1688.495 1187.635 1688.540 ;
        RECT 1202.050 1688.480 1202.370 1688.540 ;
        RECT 141.290 1688.000 141.610 1688.060 ;
        RECT 1187.345 1688.000 1187.635 1688.045 ;
        RECT 141.290 1687.860 1187.635 1688.000 ;
        RECT 141.290 1687.800 141.610 1687.860 ;
        RECT 1187.345 1687.815 1187.635 1687.860 ;
        RECT 103.570 16.560 103.890 16.620 ;
        RECT 141.290 16.560 141.610 16.620 ;
        RECT 103.570 16.420 141.610 16.560 ;
        RECT 103.570 16.360 103.890 16.420 ;
        RECT 141.290 16.360 141.610 16.420 ;
      LAYER via ;
        RECT 1202.080 1688.480 1202.340 1688.740 ;
        RECT 141.320 1687.800 141.580 1688.060 ;
        RECT 103.600 16.360 103.860 16.620 ;
        RECT 141.320 16.360 141.580 16.620 ;
      LAYER met2 ;
        RECT 1202.000 1700.000 1202.280 1702.400 ;
        RECT 1202.140 1688.770 1202.280 1700.000 ;
        RECT 1202.080 1688.450 1202.340 1688.770 ;
        RECT 141.320 1687.770 141.580 1688.090 ;
        RECT 141.380 16.650 141.520 1687.770 ;
        RECT 103.600 16.330 103.860 16.650 ;
        RECT 141.320 16.330 141.580 16.650 ;
        RECT 103.660 2.400 103.800 16.330 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1209.025 1449.165 1209.195 1497.275 ;
        RECT 1209.025 1352.605 1209.195 1400.715 ;
        RECT 1209.025 1256.045 1209.195 1304.155 ;
        RECT 1209.025 386.325 1209.195 434.775 ;
        RECT 1191.085 17.425 1191.255 18.275 ;
      LAYER mcon ;
        RECT 1209.025 1497.105 1209.195 1497.275 ;
        RECT 1209.025 1400.545 1209.195 1400.715 ;
        RECT 1209.025 1303.985 1209.195 1304.155 ;
        RECT 1209.025 434.605 1209.195 434.775 ;
        RECT 1191.085 18.105 1191.255 18.275 ;
      LAYER met1 ;
        RECT 1208.950 1642.440 1209.270 1642.500 ;
        RECT 1212.170 1642.440 1212.490 1642.500 ;
        RECT 1208.950 1642.300 1212.490 1642.440 ;
        RECT 1208.950 1642.240 1209.270 1642.300 ;
        RECT 1212.170 1642.240 1212.490 1642.300 ;
        RECT 1208.950 1497.260 1209.270 1497.320 ;
        RECT 1208.755 1497.120 1209.270 1497.260 ;
        RECT 1208.950 1497.060 1209.270 1497.120 ;
        RECT 1208.950 1449.320 1209.270 1449.380 ;
        RECT 1208.755 1449.180 1209.270 1449.320 ;
        RECT 1208.950 1449.120 1209.270 1449.180 ;
        RECT 1208.950 1400.700 1209.270 1400.760 ;
        RECT 1208.755 1400.560 1209.270 1400.700 ;
        RECT 1208.950 1400.500 1209.270 1400.560 ;
        RECT 1208.950 1352.760 1209.270 1352.820 ;
        RECT 1208.755 1352.620 1209.270 1352.760 ;
        RECT 1208.950 1352.560 1209.270 1352.620 ;
        RECT 1208.950 1304.140 1209.270 1304.200 ;
        RECT 1208.755 1304.000 1209.270 1304.140 ;
        RECT 1208.950 1303.940 1209.270 1304.000 ;
        RECT 1208.950 1256.200 1209.270 1256.260 ;
        RECT 1208.755 1256.060 1209.270 1256.200 ;
        RECT 1208.950 1256.000 1209.270 1256.060 ;
        RECT 1208.950 869.620 1209.270 869.680 ;
        RECT 1209.870 869.620 1210.190 869.680 ;
        RECT 1208.950 869.480 1210.190 869.620 ;
        RECT 1208.950 869.420 1209.270 869.480 ;
        RECT 1209.870 869.420 1210.190 869.480 ;
        RECT 1208.950 627.880 1209.270 627.940 ;
        RECT 1209.870 627.880 1210.190 627.940 ;
        RECT 1208.950 627.740 1210.190 627.880 ;
        RECT 1208.950 627.680 1209.270 627.740 ;
        RECT 1209.870 627.680 1210.190 627.740 ;
        RECT 1208.950 531.320 1209.270 531.380 ;
        RECT 1209.870 531.320 1210.190 531.380 ;
        RECT 1208.950 531.180 1210.190 531.320 ;
        RECT 1208.950 531.120 1209.270 531.180 ;
        RECT 1209.870 531.120 1210.190 531.180 ;
        RECT 1208.950 434.760 1209.270 434.820 ;
        RECT 1208.755 434.620 1209.270 434.760 ;
        RECT 1208.950 434.560 1209.270 434.620 ;
        RECT 1208.950 386.480 1209.270 386.540 ;
        RECT 1208.755 386.340 1209.270 386.480 ;
        RECT 1208.950 386.280 1209.270 386.340 ;
        RECT 127.490 18.260 127.810 18.320 ;
        RECT 1191.025 18.260 1191.315 18.305 ;
        RECT 127.490 18.120 1191.315 18.260 ;
        RECT 127.490 18.060 127.810 18.120 ;
        RECT 1191.025 18.075 1191.315 18.120 ;
        RECT 1191.025 17.580 1191.315 17.625 ;
        RECT 1208.950 17.580 1209.270 17.640 ;
        RECT 1191.025 17.440 1209.270 17.580 ;
        RECT 1191.025 17.395 1191.315 17.440 ;
        RECT 1208.950 17.380 1209.270 17.440 ;
      LAYER via ;
        RECT 1208.980 1642.240 1209.240 1642.500 ;
        RECT 1212.200 1642.240 1212.460 1642.500 ;
        RECT 1208.980 1497.060 1209.240 1497.320 ;
        RECT 1208.980 1449.120 1209.240 1449.380 ;
        RECT 1208.980 1400.500 1209.240 1400.760 ;
        RECT 1208.980 1352.560 1209.240 1352.820 ;
        RECT 1208.980 1303.940 1209.240 1304.200 ;
        RECT 1208.980 1256.000 1209.240 1256.260 ;
        RECT 1208.980 869.420 1209.240 869.680 ;
        RECT 1209.900 869.420 1210.160 869.680 ;
        RECT 1208.980 627.680 1209.240 627.940 ;
        RECT 1209.900 627.680 1210.160 627.940 ;
        RECT 1208.980 531.120 1209.240 531.380 ;
        RECT 1209.900 531.120 1210.160 531.380 ;
        RECT 1208.980 434.560 1209.240 434.820 ;
        RECT 1208.980 386.280 1209.240 386.540 ;
        RECT 127.520 18.060 127.780 18.320 ;
        RECT 1208.980 17.380 1209.240 17.640 ;
      LAYER met2 ;
        RECT 1213.960 1700.410 1214.240 1702.400 ;
        RECT 1212.260 1700.270 1214.240 1700.410 ;
        RECT 1212.260 1642.530 1212.400 1700.270 ;
        RECT 1213.960 1700.000 1214.240 1700.270 ;
        RECT 1208.980 1642.210 1209.240 1642.530 ;
        RECT 1212.200 1642.210 1212.460 1642.530 ;
        RECT 1209.040 1497.350 1209.180 1642.210 ;
        RECT 1208.980 1497.030 1209.240 1497.350 ;
        RECT 1208.980 1449.090 1209.240 1449.410 ;
        RECT 1209.040 1400.790 1209.180 1449.090 ;
        RECT 1208.980 1400.470 1209.240 1400.790 ;
        RECT 1208.980 1352.530 1209.240 1352.850 ;
        RECT 1209.040 1304.230 1209.180 1352.530 ;
        RECT 1208.980 1303.910 1209.240 1304.230 ;
        RECT 1208.980 1255.970 1209.240 1256.290 ;
        RECT 1209.040 917.845 1209.180 1255.970 ;
        RECT 1208.970 917.475 1209.250 917.845 ;
        RECT 1209.890 917.475 1210.170 917.845 ;
        RECT 1209.960 869.710 1210.100 917.475 ;
        RECT 1208.980 869.390 1209.240 869.710 ;
        RECT 1209.900 869.390 1210.160 869.710 ;
        RECT 1209.040 627.970 1209.180 869.390 ;
        RECT 1208.980 627.650 1209.240 627.970 ;
        RECT 1209.900 627.650 1210.160 627.970 ;
        RECT 1209.960 579.885 1210.100 627.650 ;
        RECT 1208.970 579.515 1209.250 579.885 ;
        RECT 1209.890 579.515 1210.170 579.885 ;
        RECT 1209.040 531.410 1209.180 579.515 ;
        RECT 1208.980 531.090 1209.240 531.410 ;
        RECT 1209.900 531.090 1210.160 531.410 ;
        RECT 1209.960 483.325 1210.100 531.090 ;
        RECT 1208.970 482.955 1209.250 483.325 ;
        RECT 1209.890 482.955 1210.170 483.325 ;
        RECT 1209.040 434.850 1209.180 482.955 ;
        RECT 1208.980 434.530 1209.240 434.850 ;
        RECT 1208.980 386.250 1209.240 386.570 ;
        RECT 127.520 18.030 127.780 18.350 ;
        RECT 127.580 2.400 127.720 18.030 ;
        RECT 1209.040 17.670 1209.180 386.250 ;
        RECT 1208.980 17.350 1209.240 17.670 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 1208.970 917.520 1209.250 917.800 ;
        RECT 1209.890 917.520 1210.170 917.800 ;
        RECT 1208.970 579.560 1209.250 579.840 ;
        RECT 1209.890 579.560 1210.170 579.840 ;
        RECT 1208.970 483.000 1209.250 483.280 ;
        RECT 1209.890 483.000 1210.170 483.280 ;
      LAYER met3 ;
        RECT 1208.945 917.810 1209.275 917.825 ;
        RECT 1209.865 917.810 1210.195 917.825 ;
        RECT 1208.945 917.510 1210.195 917.810 ;
        RECT 1208.945 917.495 1209.275 917.510 ;
        RECT 1209.865 917.495 1210.195 917.510 ;
        RECT 1208.945 579.850 1209.275 579.865 ;
        RECT 1209.865 579.850 1210.195 579.865 ;
        RECT 1208.945 579.550 1210.195 579.850 ;
        RECT 1208.945 579.535 1209.275 579.550 ;
        RECT 1209.865 579.535 1210.195 579.550 ;
        RECT 1208.945 483.290 1209.275 483.305 ;
        RECT 1209.865 483.290 1210.195 483.305 ;
        RECT 1208.945 482.990 1210.195 483.290 ;
        RECT 1208.945 482.975 1209.275 482.990 ;
        RECT 1209.865 482.975 1210.195 482.990 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 51.590 17.240 51.910 17.300 ;
        RECT 26.290 17.100 51.910 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 51.590 17.040 51.910 17.100 ;
      LAYER via ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 51.620 17.040 51.880 17.300 ;
      LAYER met2 ;
        RECT 1161.980 1700.000 1162.260 1702.400 ;
        RECT 1162.120 1686.925 1162.260 1700.000 ;
        RECT 51.610 1686.555 51.890 1686.925 ;
        RECT 1162.050 1686.555 1162.330 1686.925 ;
        RECT 51.680 17.330 51.820 1686.555 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 51.620 17.010 51.880 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 51.610 1686.600 51.890 1686.880 ;
        RECT 1162.050 1686.600 1162.330 1686.880 ;
      LAYER met3 ;
        RECT 51.585 1686.890 51.915 1686.905 ;
        RECT 1162.025 1686.890 1162.355 1686.905 ;
        RECT 51.585 1686.590 1162.355 1686.890 ;
        RECT 51.585 1686.575 51.915 1686.590 ;
        RECT 1162.025 1686.575 1162.355 1686.590 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1159.805 1490.645 1159.975 1579.895 ;
        RECT 1159.345 1297.185 1159.515 1318.095 ;
        RECT 1160.725 814.385 1160.895 903.975 ;
        RECT 1160.725 758.965 1160.895 807.075 ;
        RECT 1159.805 620.925 1159.975 710.515 ;
        RECT 1160.725 476.085 1160.895 524.195 ;
        RECT 1159.805 379.525 1159.975 427.635 ;
      LAYER mcon ;
        RECT 1159.805 1579.725 1159.975 1579.895 ;
        RECT 1159.345 1317.925 1159.515 1318.095 ;
        RECT 1160.725 903.805 1160.895 903.975 ;
        RECT 1160.725 806.905 1160.895 807.075 ;
        RECT 1159.805 710.345 1159.975 710.515 ;
        RECT 1160.725 524.025 1160.895 524.195 ;
        RECT 1159.805 427.465 1159.975 427.635 ;
      LAYER met1 ;
        RECT 1159.730 1656.380 1160.050 1656.440 ;
        RECT 1163.870 1656.380 1164.190 1656.440 ;
        RECT 1159.730 1656.240 1164.190 1656.380 ;
        RECT 1159.730 1656.180 1160.050 1656.240 ;
        RECT 1163.870 1656.180 1164.190 1656.240 ;
        RECT 1159.730 1607.900 1160.050 1608.160 ;
        RECT 1159.820 1607.420 1159.960 1607.900 ;
        RECT 1160.190 1607.420 1160.510 1607.480 ;
        RECT 1159.820 1607.280 1160.510 1607.420 ;
        RECT 1160.190 1607.220 1160.510 1607.280 ;
        RECT 1159.745 1579.880 1160.035 1579.925 ;
        RECT 1160.190 1579.880 1160.510 1579.940 ;
        RECT 1159.745 1579.740 1160.510 1579.880 ;
        RECT 1159.745 1579.695 1160.035 1579.740 ;
        RECT 1160.190 1579.680 1160.510 1579.740 ;
        RECT 1159.745 1490.800 1160.035 1490.845 ;
        RECT 1160.190 1490.800 1160.510 1490.860 ;
        RECT 1159.745 1490.660 1160.510 1490.800 ;
        RECT 1159.745 1490.615 1160.035 1490.660 ;
        RECT 1160.190 1490.600 1160.510 1490.660 ;
        RECT 1159.730 1429.600 1160.050 1429.660 ;
        RECT 1161.570 1429.600 1161.890 1429.660 ;
        RECT 1159.730 1429.460 1161.890 1429.600 ;
        RECT 1159.730 1429.400 1160.050 1429.460 ;
        RECT 1161.570 1429.400 1161.890 1429.460 ;
        RECT 1160.190 1352.760 1160.510 1352.820 ;
        RECT 1161.570 1352.760 1161.890 1352.820 ;
        RECT 1160.190 1352.620 1161.890 1352.760 ;
        RECT 1160.190 1352.560 1160.510 1352.620 ;
        RECT 1161.570 1352.560 1161.890 1352.620 ;
        RECT 1159.285 1318.080 1159.575 1318.125 ;
        RECT 1159.730 1318.080 1160.050 1318.140 ;
        RECT 1159.285 1317.940 1160.050 1318.080 ;
        RECT 1159.285 1317.895 1159.575 1317.940 ;
        RECT 1159.730 1317.880 1160.050 1317.940 ;
        RECT 1159.270 1297.340 1159.590 1297.400 ;
        RECT 1159.075 1297.200 1159.590 1297.340 ;
        RECT 1159.270 1297.140 1159.590 1297.200 ;
        RECT 1159.270 1273.200 1159.590 1273.260 ;
        RECT 1160.190 1273.200 1160.510 1273.260 ;
        RECT 1159.270 1273.060 1160.510 1273.200 ;
        RECT 1159.270 1273.000 1159.590 1273.060 ;
        RECT 1160.190 1273.000 1160.510 1273.060 ;
        RECT 1160.190 1221.860 1160.510 1221.920 ;
        RECT 1159.820 1221.720 1160.510 1221.860 ;
        RECT 1159.820 1221.240 1159.960 1221.720 ;
        RECT 1160.190 1221.660 1160.510 1221.720 ;
        RECT 1159.730 1220.980 1160.050 1221.240 ;
        RECT 1159.730 1200.440 1160.050 1200.500 ;
        RECT 1161.110 1200.440 1161.430 1200.500 ;
        RECT 1159.730 1200.300 1161.430 1200.440 ;
        RECT 1159.730 1200.240 1160.050 1200.300 ;
        RECT 1161.110 1200.240 1161.430 1200.300 ;
        RECT 1159.730 1111.360 1160.050 1111.420 ;
        RECT 1161.110 1111.360 1161.430 1111.420 ;
        RECT 1159.730 1111.220 1161.430 1111.360 ;
        RECT 1159.730 1111.160 1160.050 1111.220 ;
        RECT 1161.110 1111.160 1161.430 1111.220 ;
        RECT 1158.810 1076.340 1159.130 1076.400 ;
        RECT 1159.730 1076.340 1160.050 1076.400 ;
        RECT 1158.810 1076.200 1160.050 1076.340 ;
        RECT 1158.810 1076.140 1159.130 1076.200 ;
        RECT 1159.730 1076.140 1160.050 1076.200 ;
        RECT 1159.730 1014.460 1160.050 1014.520 ;
        RECT 1160.190 1014.460 1160.510 1014.520 ;
        RECT 1159.730 1014.320 1160.510 1014.460 ;
        RECT 1159.730 1014.260 1160.050 1014.320 ;
        RECT 1160.190 1014.260 1160.510 1014.320 ;
        RECT 1160.650 903.960 1160.970 904.020 ;
        RECT 1160.455 903.820 1160.970 903.960 ;
        RECT 1160.650 903.760 1160.970 903.820 ;
        RECT 1160.650 814.540 1160.970 814.600 ;
        RECT 1160.455 814.400 1160.970 814.540 ;
        RECT 1160.650 814.340 1160.970 814.400 ;
        RECT 1160.650 807.060 1160.970 807.120 ;
        RECT 1160.455 806.920 1160.970 807.060 ;
        RECT 1160.650 806.860 1160.970 806.920 ;
        RECT 1160.665 759.120 1160.955 759.165 ;
        RECT 1161.110 759.120 1161.430 759.180 ;
        RECT 1160.665 758.980 1161.430 759.120 ;
        RECT 1160.665 758.935 1160.955 758.980 ;
        RECT 1161.110 758.920 1161.430 758.980 ;
        RECT 1159.730 717.640 1160.050 717.700 ;
        RECT 1160.190 717.640 1160.510 717.700 ;
        RECT 1159.730 717.500 1160.510 717.640 ;
        RECT 1159.730 717.440 1160.050 717.500 ;
        RECT 1160.190 717.440 1160.510 717.500 ;
        RECT 1159.745 710.500 1160.035 710.545 ;
        RECT 1160.190 710.500 1160.510 710.560 ;
        RECT 1159.745 710.360 1160.510 710.500 ;
        RECT 1159.745 710.315 1160.035 710.360 ;
        RECT 1160.190 710.300 1160.510 710.360 ;
        RECT 1159.730 621.080 1160.050 621.140 ;
        RECT 1159.535 620.940 1160.050 621.080 ;
        RECT 1159.730 620.880 1160.050 620.940 ;
        RECT 1159.730 530.980 1160.050 531.040 ;
        RECT 1160.650 530.980 1160.970 531.040 ;
        RECT 1159.730 530.840 1160.970 530.980 ;
        RECT 1159.730 530.780 1160.050 530.840 ;
        RECT 1160.650 530.780 1160.970 530.840 ;
        RECT 1160.650 524.180 1160.970 524.240 ;
        RECT 1160.455 524.040 1160.970 524.180 ;
        RECT 1160.650 523.980 1160.970 524.040 ;
        RECT 1160.665 476.240 1160.955 476.285 ;
        RECT 1161.110 476.240 1161.430 476.300 ;
        RECT 1160.665 476.100 1161.430 476.240 ;
        RECT 1160.665 476.055 1160.955 476.100 ;
        RECT 1161.110 476.040 1161.430 476.100 ;
        RECT 1159.730 427.620 1160.050 427.680 ;
        RECT 1159.535 427.480 1160.050 427.620 ;
        RECT 1159.730 427.420 1160.050 427.480 ;
        RECT 1159.730 379.680 1160.050 379.740 ;
        RECT 1159.535 379.540 1160.050 379.680 ;
        RECT 1159.730 379.480 1160.050 379.540 ;
        RECT 1159.270 338.200 1159.590 338.260 ;
        RECT 1159.730 338.200 1160.050 338.260 ;
        RECT 1159.270 338.060 1160.050 338.200 ;
        RECT 1159.270 338.000 1159.590 338.060 ;
        RECT 1159.730 338.000 1160.050 338.060 ;
        RECT 1159.270 234.500 1159.590 234.560 ;
        RECT 1160.190 234.500 1160.510 234.560 ;
        RECT 1159.270 234.360 1160.510 234.500 ;
        RECT 1159.270 234.300 1159.590 234.360 ;
        RECT 1160.190 234.300 1160.510 234.360 ;
        RECT 1159.270 144.740 1159.590 144.800 ;
        RECT 1160.190 144.740 1160.510 144.800 ;
        RECT 1159.270 144.600 1160.510 144.740 ;
        RECT 1159.270 144.540 1159.590 144.600 ;
        RECT 1160.190 144.540 1160.510 144.600 ;
        RECT 1159.270 96.260 1159.590 96.520 ;
        RECT 1159.360 96.120 1159.500 96.260 ;
        RECT 1159.730 96.120 1160.050 96.180 ;
        RECT 1159.360 95.980 1160.050 96.120 ;
        RECT 1159.730 95.920 1160.050 95.980 ;
      LAYER via ;
        RECT 1159.760 1656.180 1160.020 1656.440 ;
        RECT 1163.900 1656.180 1164.160 1656.440 ;
        RECT 1159.760 1607.900 1160.020 1608.160 ;
        RECT 1160.220 1607.220 1160.480 1607.480 ;
        RECT 1160.220 1579.680 1160.480 1579.940 ;
        RECT 1160.220 1490.600 1160.480 1490.860 ;
        RECT 1159.760 1429.400 1160.020 1429.660 ;
        RECT 1161.600 1429.400 1161.860 1429.660 ;
        RECT 1160.220 1352.560 1160.480 1352.820 ;
        RECT 1161.600 1352.560 1161.860 1352.820 ;
        RECT 1159.760 1317.880 1160.020 1318.140 ;
        RECT 1159.300 1297.140 1159.560 1297.400 ;
        RECT 1159.300 1273.000 1159.560 1273.260 ;
        RECT 1160.220 1273.000 1160.480 1273.260 ;
        RECT 1160.220 1221.660 1160.480 1221.920 ;
        RECT 1159.760 1220.980 1160.020 1221.240 ;
        RECT 1159.760 1200.240 1160.020 1200.500 ;
        RECT 1161.140 1200.240 1161.400 1200.500 ;
        RECT 1159.760 1111.160 1160.020 1111.420 ;
        RECT 1161.140 1111.160 1161.400 1111.420 ;
        RECT 1158.840 1076.140 1159.100 1076.400 ;
        RECT 1159.760 1076.140 1160.020 1076.400 ;
        RECT 1159.760 1014.260 1160.020 1014.520 ;
        RECT 1160.220 1014.260 1160.480 1014.520 ;
        RECT 1160.680 903.760 1160.940 904.020 ;
        RECT 1160.680 814.340 1160.940 814.600 ;
        RECT 1160.680 806.860 1160.940 807.120 ;
        RECT 1161.140 758.920 1161.400 759.180 ;
        RECT 1159.760 717.440 1160.020 717.700 ;
        RECT 1160.220 717.440 1160.480 717.700 ;
        RECT 1160.220 710.300 1160.480 710.560 ;
        RECT 1159.760 620.880 1160.020 621.140 ;
        RECT 1159.760 530.780 1160.020 531.040 ;
        RECT 1160.680 530.780 1160.940 531.040 ;
        RECT 1160.680 523.980 1160.940 524.240 ;
        RECT 1161.140 476.040 1161.400 476.300 ;
        RECT 1159.760 427.420 1160.020 427.680 ;
        RECT 1159.760 379.480 1160.020 379.740 ;
        RECT 1159.300 338.000 1159.560 338.260 ;
        RECT 1159.760 338.000 1160.020 338.260 ;
        RECT 1159.300 234.300 1159.560 234.560 ;
        RECT 1160.220 234.300 1160.480 234.560 ;
        RECT 1159.300 144.540 1159.560 144.800 ;
        RECT 1160.220 144.540 1160.480 144.800 ;
        RECT 1159.300 96.260 1159.560 96.520 ;
        RECT 1159.760 95.920 1160.020 96.180 ;
      LAYER met2 ;
        RECT 1165.200 1700.410 1165.480 1702.400 ;
        RECT 1163.960 1700.270 1165.480 1700.410 ;
        RECT 1163.960 1656.470 1164.100 1700.270 ;
        RECT 1165.200 1700.000 1165.480 1700.270 ;
        RECT 1159.760 1656.150 1160.020 1656.470 ;
        RECT 1163.900 1656.150 1164.160 1656.470 ;
        RECT 1159.820 1608.190 1159.960 1656.150 ;
        RECT 1159.760 1607.870 1160.020 1608.190 ;
        RECT 1160.220 1607.190 1160.480 1607.510 ;
        RECT 1160.280 1579.970 1160.420 1607.190 ;
        RECT 1160.220 1579.650 1160.480 1579.970 ;
        RECT 1160.220 1490.570 1160.480 1490.890 ;
        RECT 1160.280 1490.290 1160.420 1490.570 ;
        RECT 1160.280 1490.150 1160.880 1490.290 ;
        RECT 1160.740 1462.410 1160.880 1490.150 ;
        RECT 1159.820 1462.270 1160.880 1462.410 ;
        RECT 1159.820 1429.690 1159.960 1462.270 ;
        RECT 1159.760 1429.370 1160.020 1429.690 ;
        RECT 1161.600 1429.370 1161.860 1429.690 ;
        RECT 1161.660 1352.850 1161.800 1429.370 ;
        RECT 1160.220 1352.530 1160.480 1352.850 ;
        RECT 1161.600 1352.530 1161.860 1352.850 ;
        RECT 1160.280 1345.450 1160.420 1352.530 ;
        RECT 1159.820 1345.310 1160.420 1345.450 ;
        RECT 1159.820 1318.170 1159.960 1345.310 ;
        RECT 1159.760 1317.850 1160.020 1318.170 ;
        RECT 1159.300 1297.110 1159.560 1297.430 ;
        RECT 1159.360 1273.290 1159.500 1297.110 ;
        RECT 1159.300 1272.970 1159.560 1273.290 ;
        RECT 1160.220 1272.970 1160.480 1273.290 ;
        RECT 1160.280 1221.950 1160.420 1272.970 ;
        RECT 1160.220 1221.630 1160.480 1221.950 ;
        RECT 1159.760 1220.950 1160.020 1221.270 ;
        RECT 1159.820 1200.530 1159.960 1220.950 ;
        RECT 1159.760 1200.210 1160.020 1200.530 ;
        RECT 1161.140 1200.210 1161.400 1200.530 ;
        RECT 1161.200 1111.450 1161.340 1200.210 ;
        RECT 1159.760 1111.130 1160.020 1111.450 ;
        RECT 1161.140 1111.130 1161.400 1111.450 ;
        RECT 1159.820 1104.165 1159.960 1111.130 ;
        RECT 1158.830 1103.795 1159.110 1104.165 ;
        RECT 1159.750 1103.795 1160.030 1104.165 ;
        RECT 1158.900 1076.430 1159.040 1103.795 ;
        RECT 1158.840 1076.110 1159.100 1076.430 ;
        RECT 1159.760 1076.110 1160.020 1076.430 ;
        RECT 1159.820 1055.770 1159.960 1076.110 ;
        RECT 1159.820 1055.630 1160.420 1055.770 ;
        RECT 1160.280 1014.550 1160.420 1055.630 ;
        RECT 1159.760 1014.230 1160.020 1014.550 ;
        RECT 1160.220 1014.230 1160.480 1014.550 ;
        RECT 1159.820 931.330 1159.960 1014.230 ;
        RECT 1159.820 931.190 1160.420 931.330 ;
        RECT 1160.280 910.930 1160.420 931.190 ;
        RECT 1160.280 910.790 1160.880 910.930 ;
        RECT 1160.740 904.050 1160.880 910.790 ;
        RECT 1160.680 903.730 1160.940 904.050 ;
        RECT 1160.680 814.310 1160.940 814.630 ;
        RECT 1160.740 807.150 1160.880 814.310 ;
        RECT 1160.680 806.830 1160.940 807.150 ;
        RECT 1161.140 758.890 1161.400 759.210 ;
        RECT 1161.200 717.925 1161.340 758.890 ;
        RECT 1159.750 717.555 1160.030 717.925 ;
        RECT 1159.760 717.410 1160.020 717.555 ;
        RECT 1160.220 717.410 1160.480 717.730 ;
        RECT 1161.130 717.555 1161.410 717.925 ;
        RECT 1160.280 710.590 1160.420 717.410 ;
        RECT 1160.220 710.270 1160.480 710.590 ;
        RECT 1159.760 620.850 1160.020 621.170 ;
        RECT 1159.820 531.070 1159.960 620.850 ;
        RECT 1159.760 530.750 1160.020 531.070 ;
        RECT 1160.680 530.750 1160.940 531.070 ;
        RECT 1160.740 524.270 1160.880 530.750 ;
        RECT 1160.680 523.950 1160.940 524.270 ;
        RECT 1161.140 476.010 1161.400 476.330 ;
        RECT 1161.200 435.045 1161.340 476.010 ;
        RECT 1159.750 434.675 1160.030 435.045 ;
        RECT 1161.130 434.675 1161.410 435.045 ;
        RECT 1159.820 427.710 1159.960 434.675 ;
        RECT 1159.760 427.390 1160.020 427.710 ;
        RECT 1159.760 379.450 1160.020 379.770 ;
        RECT 1159.820 362.850 1159.960 379.450 ;
        RECT 1159.360 362.710 1159.960 362.850 ;
        RECT 1159.360 338.290 1159.500 362.710 ;
        RECT 1159.300 337.970 1159.560 338.290 ;
        RECT 1159.760 337.970 1160.020 338.290 ;
        RECT 1159.820 290.090 1159.960 337.970 ;
        RECT 1159.820 289.950 1160.420 290.090 ;
        RECT 1160.280 283.290 1160.420 289.950 ;
        RECT 1159.360 283.150 1160.420 283.290 ;
        RECT 1159.360 234.590 1159.500 283.150 ;
        RECT 1159.300 234.270 1159.560 234.590 ;
        RECT 1160.220 234.270 1160.480 234.590 ;
        RECT 1160.280 144.830 1160.420 234.270 ;
        RECT 1159.300 144.510 1159.560 144.830 ;
        RECT 1160.220 144.510 1160.480 144.830 ;
        RECT 1159.360 96.550 1159.500 144.510 ;
        RECT 1159.300 96.230 1159.560 96.550 ;
        RECT 1159.760 95.890 1160.020 96.210 ;
        RECT 1159.820 16.845 1159.960 95.890 ;
        RECT 32.290 16.475 32.570 16.845 ;
        RECT 1159.750 16.475 1160.030 16.845 ;
        RECT 32.360 2.400 32.500 16.475 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 1158.830 1103.840 1159.110 1104.120 ;
        RECT 1159.750 1103.840 1160.030 1104.120 ;
        RECT 1159.750 717.600 1160.030 717.880 ;
        RECT 1161.130 717.600 1161.410 717.880 ;
        RECT 1159.750 434.720 1160.030 435.000 ;
        RECT 1161.130 434.720 1161.410 435.000 ;
        RECT 32.290 16.520 32.570 16.800 ;
        RECT 1159.750 16.520 1160.030 16.800 ;
      LAYER met3 ;
        RECT 1158.805 1104.130 1159.135 1104.145 ;
        RECT 1159.725 1104.130 1160.055 1104.145 ;
        RECT 1158.805 1103.830 1160.055 1104.130 ;
        RECT 1158.805 1103.815 1159.135 1103.830 ;
        RECT 1159.725 1103.815 1160.055 1103.830 ;
        RECT 1159.725 717.890 1160.055 717.905 ;
        RECT 1161.105 717.890 1161.435 717.905 ;
        RECT 1159.725 717.590 1161.435 717.890 ;
        RECT 1159.725 717.575 1160.055 717.590 ;
        RECT 1161.105 717.575 1161.435 717.590 ;
        RECT 1159.725 435.010 1160.055 435.025 ;
        RECT 1161.105 435.010 1161.435 435.025 ;
        RECT 1159.725 434.710 1161.435 435.010 ;
        RECT 1159.725 434.695 1160.055 434.710 ;
        RECT 1161.105 434.695 1161.435 434.710 ;
        RECT 32.265 16.810 32.595 16.825 ;
        RECT 1159.725 16.810 1160.055 16.825 ;
        RECT 32.265 16.510 1160.055 16.810 ;
        RECT 32.265 16.495 32.595 16.510 ;
        RECT 1159.725 16.495 1160.055 16.510 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 -9.220 907.020 3528.900 ;
        RECT 1084.020 -9.220 1087.020 3528.900 ;
        RECT 1264.020 -9.220 1267.020 3528.900 ;
        RECT 1444.020 -9.220 1447.020 3528.900 ;
        RECT 1624.020 -9.220 1627.020 3528.900 ;
        RECT 1804.020 -9.220 1807.020 3528.900 ;
        RECT 1984.020 -9.220 1987.020 3528.900 ;
        RECT 2164.020 -9.220 2167.020 3528.900 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 -9.220 817.020 3528.900 ;
        RECT 994.020 -9.220 997.020 3528.900 ;
        RECT 1174.020 -9.220 1177.020 3528.900 ;
        RECT 1354.020 -9.220 1357.020 3528.900 ;
        RECT 1534.020 -9.220 1537.020 3528.900 ;
        RECT 1714.020 -9.220 1717.020 3528.900 ;
        RECT 1894.020 -9.220 1897.020 3528.900 ;
        RECT 2074.020 -9.220 2077.020 3528.900 ;
        RECT 2254.020 -9.220 2257.020 3528.900 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 -18.420 745.020 3538.100 ;
        RECT 922.020 -18.420 925.020 3538.100 ;
        RECT 1102.020 -18.420 1105.020 3538.100 ;
        RECT 1282.020 -18.420 1285.020 3538.100 ;
        RECT 1462.020 -18.420 1465.020 3538.100 ;
        RECT 1642.020 -18.420 1645.020 3538.100 ;
        RECT 1822.020 -18.420 1825.020 3538.100 ;
        RECT 2002.020 -18.420 2005.020 3538.100 ;
        RECT 2182.020 -18.420 2185.020 3538.100 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 -18.420 835.020 3538.100 ;
        RECT 1012.020 -18.420 1015.020 3538.100 ;
        RECT 1192.020 -18.420 1195.020 3538.100 ;
        RECT 1372.020 -18.420 1375.020 3538.100 ;
        RECT 1552.020 -18.420 1555.020 3538.100 ;
        RECT 1732.020 -18.420 1735.020 3538.100 ;
        RECT 1912.020 -18.420 1915.020 3538.100 ;
        RECT 2092.020 -18.420 2095.020 3538.100 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 -27.620 763.020 3547.300 ;
        RECT 940.020 -27.620 943.020 3547.300 ;
        RECT 1120.020 -27.620 1123.020 3547.300 ;
        RECT 1300.020 -27.620 1303.020 3547.300 ;
        RECT 1480.020 -27.620 1483.020 3547.300 ;
        RECT 1660.020 -27.620 1663.020 3547.300 ;
        RECT 1840.020 -27.620 1843.020 3547.300 ;
        RECT 2020.020 -27.620 2023.020 3547.300 ;
        RECT 2200.020 -27.620 2203.020 3547.300 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 -27.620 853.020 3547.300 ;
        RECT 1030.020 -27.620 1033.020 3547.300 ;
        RECT 1210.020 -27.620 1213.020 3547.300 ;
        RECT 1390.020 -27.620 1393.020 3547.300 ;
        RECT 1570.020 -27.620 1573.020 3547.300 ;
        RECT 1750.020 -27.620 1753.020 3547.300 ;
        RECT 1930.020 -27.620 1933.020 3547.300 ;
        RECT 2110.020 -27.620 2113.020 3547.300 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 -36.820 781.020 3556.500 ;
        RECT 958.020 -36.820 961.020 3556.500 ;
        RECT 1138.020 -36.820 1141.020 3556.500 ;
        RECT 1318.020 -36.820 1321.020 3556.500 ;
        RECT 1498.020 -36.820 1501.020 3556.500 ;
        RECT 1678.020 -36.820 1681.020 3556.500 ;
        RECT 1858.020 -36.820 1861.020 3556.500 ;
        RECT 2038.020 -36.820 2041.020 3556.500 ;
        RECT 2218.020 -36.820 2221.020 3556.500 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 -36.820 871.020 3556.500 ;
        RECT 1048.020 -36.820 1051.020 3556.500 ;
        RECT 1228.020 -36.820 1231.020 3556.500 ;
        RECT 1408.020 -36.820 1411.020 3556.500 ;
        RECT 1588.020 -36.820 1591.020 3556.500 ;
        RECT 1768.020 -36.820 1771.020 3556.500 ;
        RECT 1948.020 -36.820 1951.020 3556.500 ;
        RECT 2128.020 -36.820 2131.020 3556.500 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1154.070 1710.795 2642.630 3187.925 ;
      LAYER met1 ;
        RECT 1150.000 1702.760 2647.160 3197.320 ;
      LAYER met2 ;
        RECT 1150.030 3197.320 1154.800 3197.600 ;
        RECT 1155.640 3197.320 1167.680 3197.600 ;
        RECT 1168.520 3197.320 1181.020 3197.600 ;
        RECT 1181.860 3197.320 1193.900 3197.600 ;
        RECT 1194.740 3197.320 1207.240 3197.600 ;
        RECT 1208.080 3197.320 1220.580 3197.600 ;
        RECT 1221.420 3197.320 1233.460 3197.600 ;
        RECT 1234.300 3197.320 1246.800 3197.600 ;
        RECT 1247.640 3197.320 1259.680 3197.600 ;
        RECT 1260.520 3197.320 1273.020 3197.600 ;
        RECT 1273.860 3197.320 1286.360 3197.600 ;
        RECT 1287.200 3197.320 1299.240 3197.600 ;
        RECT 1300.080 3197.320 1312.580 3197.600 ;
        RECT 1313.420 3197.320 1325.460 3197.600 ;
        RECT 1326.300 3197.320 1338.800 3197.600 ;
        RECT 1339.640 3197.320 1352.140 3197.600 ;
        RECT 1352.980 3197.320 1365.020 3197.600 ;
        RECT 1365.860 3197.320 1378.360 3197.600 ;
        RECT 1379.200 3197.320 1391.240 3197.600 ;
        RECT 1392.080 3197.320 1404.580 3197.600 ;
        RECT 1405.420 3197.320 1417.920 3197.600 ;
        RECT 1418.760 3197.320 1430.800 3197.600 ;
        RECT 1431.640 3197.320 1444.140 3197.600 ;
        RECT 1444.980 3197.320 1457.020 3197.600 ;
        RECT 1457.860 3197.320 1470.360 3197.600 ;
        RECT 1471.200 3197.320 1483.700 3197.600 ;
        RECT 1484.540 3197.320 1496.580 3197.600 ;
        RECT 1497.420 3197.320 1509.920 3197.600 ;
        RECT 1510.760 3197.320 1522.800 3197.600 ;
        RECT 1523.640 3197.320 1536.140 3197.600 ;
        RECT 1536.980 3197.320 1549.480 3197.600 ;
        RECT 1550.320 3197.320 1562.360 3197.600 ;
        RECT 1563.200 3197.320 1575.700 3197.600 ;
        RECT 1576.540 3197.320 1588.580 3197.600 ;
        RECT 1589.420 3197.320 1601.920 3197.600 ;
        RECT 1602.760 3197.320 1615.260 3197.600 ;
        RECT 1616.100 3197.320 1628.140 3197.600 ;
        RECT 1628.980 3197.320 1641.480 3197.600 ;
        RECT 1642.320 3197.320 1654.820 3197.600 ;
        RECT 1655.660 3197.320 1667.700 3197.600 ;
        RECT 1668.540 3197.320 1681.040 3197.600 ;
        RECT 1681.880 3197.320 1693.920 3197.600 ;
        RECT 1694.760 3197.320 1707.260 3197.600 ;
        RECT 1708.100 3197.320 1720.600 3197.600 ;
        RECT 1721.440 3197.320 1733.480 3197.600 ;
        RECT 1734.320 3197.320 1746.820 3197.600 ;
        RECT 1747.660 3197.320 1759.700 3197.600 ;
        RECT 1760.540 3197.320 1773.040 3197.600 ;
        RECT 1773.880 3197.320 1786.380 3197.600 ;
        RECT 1787.220 3197.320 1799.260 3197.600 ;
        RECT 1800.100 3197.320 1812.600 3197.600 ;
        RECT 1813.440 3197.320 1825.480 3197.600 ;
        RECT 1826.320 3197.320 1838.820 3197.600 ;
        RECT 1839.660 3197.320 1852.160 3197.600 ;
        RECT 1853.000 3197.320 1865.040 3197.600 ;
        RECT 1865.880 3197.320 1878.380 3197.600 ;
        RECT 1879.220 3197.320 1891.260 3197.600 ;
        RECT 1892.100 3197.320 1904.600 3197.600 ;
        RECT 1905.440 3197.320 1917.940 3197.600 ;
        RECT 1918.780 3197.320 1930.820 3197.600 ;
        RECT 1931.660 3197.320 1944.160 3197.600 ;
        RECT 1945.000 3197.320 1957.040 3197.600 ;
        RECT 1957.880 3197.320 1970.380 3197.600 ;
        RECT 1971.220 3197.320 1983.720 3197.600 ;
        RECT 1984.560 3197.320 1996.600 3197.600 ;
        RECT 1997.440 3197.320 2009.940 3197.600 ;
        RECT 2010.780 3197.320 2022.820 3197.600 ;
        RECT 2023.660 3197.320 2036.160 3197.600 ;
        RECT 2037.000 3197.320 2049.500 3197.600 ;
        RECT 2050.340 3197.320 2062.380 3197.600 ;
        RECT 2063.220 3197.320 2075.720 3197.600 ;
        RECT 2076.560 3197.320 2088.600 3197.600 ;
        RECT 2089.440 3197.320 2101.940 3197.600 ;
        RECT 2102.780 3197.320 2115.280 3197.600 ;
        RECT 2116.120 3197.320 2128.160 3197.600 ;
        RECT 2129.000 3197.320 2141.500 3197.600 ;
        RECT 2142.340 3197.320 2154.840 3197.600 ;
        RECT 2155.680 3197.320 2167.720 3197.600 ;
        RECT 2168.560 3197.320 2181.060 3197.600 ;
        RECT 2181.900 3197.320 2193.940 3197.600 ;
        RECT 2194.780 3197.320 2207.280 3197.600 ;
        RECT 2208.120 3197.320 2220.620 3197.600 ;
        RECT 2221.460 3197.320 2233.500 3197.600 ;
        RECT 2234.340 3197.320 2246.840 3197.600 ;
        RECT 2247.680 3197.320 2259.720 3197.600 ;
        RECT 2260.560 3197.320 2273.060 3197.600 ;
        RECT 2273.900 3197.320 2286.400 3197.600 ;
        RECT 2287.240 3197.320 2299.280 3197.600 ;
        RECT 2300.120 3197.320 2312.620 3197.600 ;
        RECT 2313.460 3197.320 2325.500 3197.600 ;
        RECT 2326.340 3197.320 2338.840 3197.600 ;
        RECT 2339.680 3197.320 2352.180 3197.600 ;
        RECT 2353.020 3197.320 2365.060 3197.600 ;
        RECT 2365.900 3197.320 2378.400 3197.600 ;
        RECT 2379.240 3197.320 2391.280 3197.600 ;
        RECT 2392.120 3197.320 2404.620 3197.600 ;
        RECT 2405.460 3197.320 2417.960 3197.600 ;
        RECT 2418.800 3197.320 2430.840 3197.600 ;
        RECT 2431.680 3197.320 2444.180 3197.600 ;
        RECT 2445.020 3197.320 2457.060 3197.600 ;
        RECT 2457.900 3197.320 2470.400 3197.600 ;
        RECT 2471.240 3197.320 2483.740 3197.600 ;
        RECT 2484.580 3197.320 2496.620 3197.600 ;
        RECT 2497.460 3197.320 2509.960 3197.600 ;
        RECT 2510.800 3197.320 2522.840 3197.600 ;
        RECT 2523.680 3197.320 2536.180 3197.600 ;
        RECT 2537.020 3197.320 2549.520 3197.600 ;
        RECT 2550.360 3197.320 2562.400 3197.600 ;
        RECT 2563.240 3197.320 2575.740 3197.600 ;
        RECT 2576.580 3197.320 2588.620 3197.600 ;
        RECT 2589.460 3197.320 2601.960 3197.600 ;
        RECT 2602.800 3197.320 2615.300 3197.600 ;
        RECT 2616.140 3197.320 2628.180 3197.600 ;
        RECT 2629.020 3197.320 2641.520 3197.600 ;
        RECT 2642.360 3197.320 2647.130 3197.600 ;
        RECT 1150.030 1702.680 2647.130 3197.320 ;
        RECT 1150.580 1702.400 1152.500 1702.680 ;
        RECT 1153.340 1702.400 1155.720 1702.680 ;
        RECT 1156.560 1702.400 1158.480 1702.680 ;
        RECT 1159.320 1702.400 1161.700 1702.680 ;
        RECT 1162.540 1702.400 1164.920 1702.680 ;
        RECT 1165.760 1702.400 1167.680 1702.680 ;
        RECT 1168.520 1702.400 1170.900 1702.680 ;
        RECT 1171.740 1702.400 1174.120 1702.680 ;
        RECT 1174.960 1702.400 1176.880 1702.680 ;
        RECT 1177.720 1702.400 1180.100 1702.680 ;
        RECT 1180.940 1702.400 1183.320 1702.680 ;
        RECT 1184.160 1702.400 1186.080 1702.680 ;
        RECT 1186.920 1702.400 1189.300 1702.680 ;
        RECT 1190.140 1702.400 1192.520 1702.680 ;
        RECT 1193.360 1702.400 1195.280 1702.680 ;
        RECT 1196.120 1702.400 1198.500 1702.680 ;
        RECT 1199.340 1702.400 1201.720 1702.680 ;
        RECT 1202.560 1702.400 1204.480 1702.680 ;
        RECT 1205.320 1702.400 1207.700 1702.680 ;
        RECT 1208.540 1702.400 1210.920 1702.680 ;
        RECT 1211.760 1702.400 1213.680 1702.680 ;
        RECT 1214.520 1702.400 1216.900 1702.680 ;
        RECT 1217.740 1702.400 1220.120 1702.680 ;
        RECT 1220.960 1702.400 1222.880 1702.680 ;
        RECT 1223.720 1702.400 1226.100 1702.680 ;
        RECT 1226.940 1702.400 1229.320 1702.680 ;
        RECT 1230.160 1702.400 1232.080 1702.680 ;
        RECT 1232.920 1702.400 1235.300 1702.680 ;
        RECT 1236.140 1702.400 1238.060 1702.680 ;
        RECT 1238.900 1702.400 1241.280 1702.680 ;
        RECT 1242.120 1702.400 1244.500 1702.680 ;
        RECT 1245.340 1702.400 1247.260 1702.680 ;
        RECT 1248.100 1702.400 1250.480 1702.680 ;
        RECT 1251.320 1702.400 1253.700 1702.680 ;
        RECT 1254.540 1702.400 1256.460 1702.680 ;
        RECT 1257.300 1702.400 1259.680 1702.680 ;
        RECT 1260.520 1702.400 1262.900 1702.680 ;
        RECT 1263.740 1702.400 1265.660 1702.680 ;
        RECT 1266.500 1702.400 1268.880 1702.680 ;
        RECT 1269.720 1702.400 1272.100 1702.680 ;
        RECT 1272.940 1702.400 1274.860 1702.680 ;
        RECT 1275.700 1702.400 1278.080 1702.680 ;
        RECT 1278.920 1702.400 1281.300 1702.680 ;
        RECT 1282.140 1702.400 1284.060 1702.680 ;
        RECT 1284.900 1702.400 1287.280 1702.680 ;
        RECT 1288.120 1702.400 1290.500 1702.680 ;
        RECT 1291.340 1702.400 1293.260 1702.680 ;
        RECT 1294.100 1702.400 1296.480 1702.680 ;
        RECT 1297.320 1702.400 1299.700 1702.680 ;
        RECT 1300.540 1702.400 1302.460 1702.680 ;
        RECT 1303.300 1702.400 1305.680 1702.680 ;
        RECT 1306.520 1702.400 1308.900 1702.680 ;
        RECT 1309.740 1702.400 1311.660 1702.680 ;
        RECT 1312.500 1702.400 1314.880 1702.680 ;
        RECT 1315.720 1702.400 1318.100 1702.680 ;
        RECT 1318.940 1702.400 1320.860 1702.680 ;
        RECT 1321.700 1702.400 1324.080 1702.680 ;
        RECT 1324.920 1702.400 1326.840 1702.680 ;
        RECT 1327.680 1702.400 1330.060 1702.680 ;
        RECT 1330.900 1702.400 1333.280 1702.680 ;
        RECT 1334.120 1702.400 1336.040 1702.680 ;
        RECT 1336.880 1702.400 1339.260 1702.680 ;
        RECT 1340.100 1702.400 1342.480 1702.680 ;
        RECT 1343.320 1702.400 1345.240 1702.680 ;
        RECT 1346.080 1702.400 1348.460 1702.680 ;
        RECT 1349.300 1702.400 1351.680 1702.680 ;
        RECT 1352.520 1702.400 1354.440 1702.680 ;
        RECT 1355.280 1702.400 1357.660 1702.680 ;
        RECT 1358.500 1702.400 1360.880 1702.680 ;
        RECT 1361.720 1702.400 1363.640 1702.680 ;
        RECT 1364.480 1702.400 1366.860 1702.680 ;
        RECT 1367.700 1702.400 1370.080 1702.680 ;
        RECT 1370.920 1702.400 1372.840 1702.680 ;
        RECT 1373.680 1702.400 1376.060 1702.680 ;
        RECT 1376.900 1702.400 1379.280 1702.680 ;
        RECT 1380.120 1702.400 1382.040 1702.680 ;
        RECT 1382.880 1702.400 1385.260 1702.680 ;
        RECT 1386.100 1702.400 1388.480 1702.680 ;
        RECT 1389.320 1702.400 1391.240 1702.680 ;
        RECT 1392.080 1702.400 1394.460 1702.680 ;
        RECT 1395.300 1702.400 1397.680 1702.680 ;
        RECT 1398.520 1702.400 1400.440 1702.680 ;
        RECT 1401.280 1702.400 1403.660 1702.680 ;
        RECT 1404.500 1702.400 1406.880 1702.680 ;
        RECT 1407.720 1702.400 1409.640 1702.680 ;
        RECT 1410.480 1702.400 1412.860 1702.680 ;
        RECT 1413.700 1702.400 1415.620 1702.680 ;
        RECT 1416.460 1702.400 1418.840 1702.680 ;
        RECT 1419.680 1702.400 1422.060 1702.680 ;
        RECT 1422.900 1702.400 1424.820 1702.680 ;
        RECT 1425.660 1702.400 1428.040 1702.680 ;
        RECT 1428.880 1702.400 1431.260 1702.680 ;
        RECT 1432.100 1702.400 1434.020 1702.680 ;
        RECT 1434.860 1702.400 1437.240 1702.680 ;
        RECT 1438.080 1702.400 1440.460 1702.680 ;
        RECT 1441.300 1702.400 1443.220 1702.680 ;
        RECT 1444.060 1702.400 1446.440 1702.680 ;
        RECT 1447.280 1702.400 1449.660 1702.680 ;
        RECT 1450.500 1702.400 1452.420 1702.680 ;
        RECT 1453.260 1702.400 1455.640 1702.680 ;
        RECT 1456.480 1702.400 1458.860 1702.680 ;
        RECT 1459.700 1702.400 1461.620 1702.680 ;
        RECT 1462.460 1702.400 1464.840 1702.680 ;
        RECT 1465.680 1702.400 1468.060 1702.680 ;
        RECT 1468.900 1702.400 1470.820 1702.680 ;
        RECT 1471.660 1702.400 1474.040 1702.680 ;
        RECT 1474.880 1702.400 1477.260 1702.680 ;
        RECT 1478.100 1702.400 1480.020 1702.680 ;
        RECT 1480.860 1702.400 1483.240 1702.680 ;
        RECT 1484.080 1702.400 1486.460 1702.680 ;
        RECT 1487.300 1702.400 1489.220 1702.680 ;
        RECT 1490.060 1702.400 1492.440 1702.680 ;
        RECT 1493.280 1702.400 1495.660 1702.680 ;
        RECT 1496.500 1702.400 1498.420 1702.680 ;
        RECT 1499.260 1702.400 1501.640 1702.680 ;
        RECT 1502.480 1702.400 1504.400 1702.680 ;
        RECT 1505.240 1702.400 1507.620 1702.680 ;
        RECT 1508.460 1702.400 1510.840 1702.680 ;
        RECT 1511.680 1702.400 1513.600 1702.680 ;
        RECT 1514.440 1702.400 1516.820 1702.680 ;
        RECT 1517.660 1702.400 1520.040 1702.680 ;
        RECT 1520.880 1702.400 1522.800 1702.680 ;
        RECT 1523.640 1702.400 1526.020 1702.680 ;
        RECT 1526.860 1702.400 1529.240 1702.680 ;
        RECT 1530.080 1702.400 1532.000 1702.680 ;
        RECT 1532.840 1702.400 1535.220 1702.680 ;
        RECT 1536.060 1702.400 1538.440 1702.680 ;
        RECT 1539.280 1702.400 1541.200 1702.680 ;
        RECT 1542.040 1702.400 1544.420 1702.680 ;
        RECT 1545.260 1702.400 1547.640 1702.680 ;
        RECT 1548.480 1702.400 1550.400 1702.680 ;
        RECT 1551.240 1702.400 1553.620 1702.680 ;
        RECT 1554.460 1702.400 1556.840 1702.680 ;
        RECT 1557.680 1702.400 1559.600 1702.680 ;
        RECT 1560.440 1702.400 1562.820 1702.680 ;
        RECT 1563.660 1702.400 1566.040 1702.680 ;
        RECT 1566.880 1702.400 1568.800 1702.680 ;
        RECT 1569.640 1702.400 1572.020 1702.680 ;
        RECT 1572.860 1702.400 1575.240 1702.680 ;
        RECT 1576.080 1702.400 1578.000 1702.680 ;
        RECT 1578.840 1702.400 1581.220 1702.680 ;
        RECT 1582.060 1702.400 1584.440 1702.680 ;
        RECT 1585.280 1702.400 1587.200 1702.680 ;
        RECT 1588.040 1702.400 1590.420 1702.680 ;
        RECT 1591.260 1702.400 1593.180 1702.680 ;
        RECT 1594.020 1702.400 1596.400 1702.680 ;
        RECT 1597.240 1702.400 1599.620 1702.680 ;
        RECT 1600.460 1702.400 1602.380 1702.680 ;
        RECT 1603.220 1702.400 1605.600 1702.680 ;
        RECT 1606.440 1702.400 1608.820 1702.680 ;
        RECT 1609.660 1702.400 1611.580 1702.680 ;
        RECT 1612.420 1702.400 1614.800 1702.680 ;
        RECT 1615.640 1702.400 1618.020 1702.680 ;
        RECT 1618.860 1702.400 1620.780 1702.680 ;
        RECT 1621.620 1702.400 1624.000 1702.680 ;
        RECT 1624.840 1702.400 1627.220 1702.680 ;
        RECT 1628.060 1702.400 1629.980 1702.680 ;
        RECT 1630.820 1702.400 1633.200 1702.680 ;
        RECT 1634.040 1702.400 1636.420 1702.680 ;
        RECT 1637.260 1702.400 1639.180 1702.680 ;
        RECT 1640.020 1702.400 1642.400 1702.680 ;
        RECT 1643.240 1702.400 1645.620 1702.680 ;
        RECT 1646.460 1702.400 1648.380 1702.680 ;
        RECT 1649.220 1702.400 1651.600 1702.680 ;
        RECT 1652.440 1702.400 1654.820 1702.680 ;
        RECT 1655.660 1702.400 1657.580 1702.680 ;
        RECT 1658.420 1702.400 1660.800 1702.680 ;
        RECT 1661.640 1702.400 1664.020 1702.680 ;
        RECT 1664.860 1702.400 1666.780 1702.680 ;
        RECT 1667.620 1702.400 1670.000 1702.680 ;
        RECT 1670.840 1702.400 1673.220 1702.680 ;
        RECT 1674.060 1702.400 1675.980 1702.680 ;
        RECT 1676.820 1702.400 1679.200 1702.680 ;
        RECT 1680.040 1702.400 1681.960 1702.680 ;
        RECT 1682.800 1702.400 1685.180 1702.680 ;
        RECT 1686.020 1702.400 1688.400 1702.680 ;
        RECT 1689.240 1702.400 1691.160 1702.680 ;
        RECT 1692.000 1702.400 1694.380 1702.680 ;
        RECT 1695.220 1702.400 1697.600 1702.680 ;
        RECT 1698.440 1702.400 1700.360 1702.680 ;
        RECT 1701.200 1702.400 1703.580 1702.680 ;
        RECT 1704.420 1702.400 1706.800 1702.680 ;
        RECT 1707.640 1702.400 1709.560 1702.680 ;
        RECT 1710.400 1702.400 1712.780 1702.680 ;
        RECT 1713.620 1702.400 1716.000 1702.680 ;
        RECT 1716.840 1702.400 1718.760 1702.680 ;
        RECT 1719.600 1702.400 1721.980 1702.680 ;
        RECT 1722.820 1702.400 1725.200 1702.680 ;
        RECT 1726.040 1702.400 1727.960 1702.680 ;
        RECT 1728.800 1702.400 1731.180 1702.680 ;
        RECT 1732.020 1702.400 1734.400 1702.680 ;
        RECT 1735.240 1702.400 1737.160 1702.680 ;
        RECT 1738.000 1702.400 1740.380 1702.680 ;
        RECT 1741.220 1702.400 1743.600 1702.680 ;
        RECT 1744.440 1702.400 1746.360 1702.680 ;
        RECT 1747.200 1702.400 1749.580 1702.680 ;
        RECT 1750.420 1702.400 1752.800 1702.680 ;
        RECT 1753.640 1702.400 1755.560 1702.680 ;
        RECT 1756.400 1702.400 1758.780 1702.680 ;
        RECT 1759.620 1702.400 1762.000 1702.680 ;
        RECT 1762.840 1702.400 1764.760 1702.680 ;
        RECT 1765.600 1702.400 1767.980 1702.680 ;
        RECT 1768.820 1702.400 1770.740 1702.680 ;
        RECT 1771.580 1702.400 1773.960 1702.680 ;
        RECT 1774.800 1702.400 1777.180 1702.680 ;
        RECT 1778.020 1702.400 1779.940 1702.680 ;
        RECT 1780.780 1702.400 1783.160 1702.680 ;
        RECT 1784.000 1702.400 1786.380 1702.680 ;
        RECT 1787.220 1702.400 1789.140 1702.680 ;
        RECT 1789.980 1702.400 1792.360 1702.680 ;
        RECT 1793.200 1702.400 1795.580 1702.680 ;
        RECT 1796.420 1702.400 1798.340 1702.680 ;
        RECT 1799.180 1702.400 1801.560 1702.680 ;
        RECT 1802.400 1702.400 1804.780 1702.680 ;
        RECT 1805.620 1702.400 1807.540 1702.680 ;
        RECT 1808.380 1702.400 1810.760 1702.680 ;
        RECT 1811.600 1702.400 1813.980 1702.680 ;
        RECT 1814.820 1702.400 1816.740 1702.680 ;
        RECT 1817.580 1702.400 1819.960 1702.680 ;
        RECT 1820.800 1702.400 1823.180 1702.680 ;
        RECT 1824.020 1702.400 1825.940 1702.680 ;
        RECT 1826.780 1702.400 1829.160 1702.680 ;
        RECT 1830.000 1702.400 1832.380 1702.680 ;
        RECT 1833.220 1702.400 1835.140 1702.680 ;
        RECT 1835.980 1702.400 1838.360 1702.680 ;
        RECT 1839.200 1702.400 1841.580 1702.680 ;
        RECT 1842.420 1702.400 1844.340 1702.680 ;
        RECT 1845.180 1702.400 1847.560 1702.680 ;
        RECT 1848.400 1702.400 1850.780 1702.680 ;
        RECT 1851.620 1702.400 1853.540 1702.680 ;
        RECT 1854.380 1702.400 1856.760 1702.680 ;
        RECT 1857.600 1702.400 1859.520 1702.680 ;
        RECT 1860.360 1702.400 1862.740 1702.680 ;
        RECT 1863.580 1702.400 1865.960 1702.680 ;
        RECT 1866.800 1702.400 1868.720 1702.680 ;
        RECT 1869.560 1702.400 1871.940 1702.680 ;
        RECT 1872.780 1702.400 1875.160 1702.680 ;
        RECT 1876.000 1702.400 1877.920 1702.680 ;
        RECT 1878.760 1702.400 1881.140 1702.680 ;
        RECT 1881.980 1702.400 1884.360 1702.680 ;
        RECT 1885.200 1702.400 1887.120 1702.680 ;
        RECT 1887.960 1702.400 1890.340 1702.680 ;
        RECT 1891.180 1702.400 1893.560 1702.680 ;
        RECT 1894.400 1702.400 1896.320 1702.680 ;
        RECT 1897.160 1702.400 1899.540 1702.680 ;
        RECT 1900.380 1702.400 1902.760 1702.680 ;
        RECT 1903.600 1702.400 1905.520 1702.680 ;
        RECT 1906.360 1702.400 1908.740 1702.680 ;
        RECT 1909.580 1702.400 1911.960 1702.680 ;
        RECT 1912.800 1702.400 1914.720 1702.680 ;
        RECT 1915.560 1702.400 1917.940 1702.680 ;
        RECT 1918.780 1702.400 1921.160 1702.680 ;
        RECT 1922.000 1702.400 1923.920 1702.680 ;
        RECT 1924.760 1702.400 1927.140 1702.680 ;
        RECT 1927.980 1702.400 1930.360 1702.680 ;
        RECT 1931.200 1702.400 1933.120 1702.680 ;
        RECT 1933.960 1702.400 1936.340 1702.680 ;
        RECT 1937.180 1702.400 1939.560 1702.680 ;
        RECT 1940.400 1702.400 1942.320 1702.680 ;
        RECT 1943.160 1702.400 1945.540 1702.680 ;
        RECT 1946.380 1702.400 1948.300 1702.680 ;
        RECT 1949.140 1702.400 1951.520 1702.680 ;
        RECT 1952.360 1702.400 1954.740 1702.680 ;
        RECT 1955.580 1702.400 1957.500 1702.680 ;
        RECT 1958.340 1702.400 1960.720 1702.680 ;
        RECT 1961.560 1702.400 1963.940 1702.680 ;
        RECT 1964.780 1702.400 1966.700 1702.680 ;
        RECT 1967.540 1702.400 1969.920 1702.680 ;
        RECT 1970.760 1702.400 1973.140 1702.680 ;
        RECT 1973.980 1702.400 1975.900 1702.680 ;
        RECT 1976.740 1702.400 1979.120 1702.680 ;
        RECT 1979.960 1702.400 1982.340 1702.680 ;
        RECT 1983.180 1702.400 1985.100 1702.680 ;
        RECT 1985.940 1702.400 1988.320 1702.680 ;
        RECT 1989.160 1702.400 1991.540 1702.680 ;
        RECT 1992.380 1702.400 1994.300 1702.680 ;
        RECT 1995.140 1702.400 1997.520 1702.680 ;
        RECT 1998.360 1702.400 2000.740 1702.680 ;
        RECT 2001.580 1702.400 2003.500 1702.680 ;
        RECT 2004.340 1702.400 2006.720 1702.680 ;
        RECT 2007.560 1702.400 2009.940 1702.680 ;
        RECT 2010.780 1702.400 2012.700 1702.680 ;
        RECT 2013.540 1702.400 2015.920 1702.680 ;
        RECT 2016.760 1702.400 2019.140 1702.680 ;
        RECT 2019.980 1702.400 2021.900 1702.680 ;
        RECT 2022.740 1702.400 2025.120 1702.680 ;
        RECT 2025.960 1702.400 2028.340 1702.680 ;
        RECT 2029.180 1702.400 2031.100 1702.680 ;
        RECT 2031.940 1702.400 2034.320 1702.680 ;
        RECT 2035.160 1702.400 2037.080 1702.680 ;
        RECT 2037.920 1702.400 2040.300 1702.680 ;
        RECT 2041.140 1702.400 2043.520 1702.680 ;
        RECT 2044.360 1702.400 2046.280 1702.680 ;
        RECT 2047.120 1702.400 2049.500 1702.680 ;
        RECT 2050.340 1702.400 2052.720 1702.680 ;
        RECT 2053.560 1702.400 2055.480 1702.680 ;
        RECT 2056.320 1702.400 2058.700 1702.680 ;
        RECT 2059.540 1702.400 2061.920 1702.680 ;
        RECT 2062.760 1702.400 2064.680 1702.680 ;
        RECT 2065.520 1702.400 2067.900 1702.680 ;
        RECT 2068.740 1702.400 2071.120 1702.680 ;
        RECT 2071.960 1702.400 2073.880 1702.680 ;
        RECT 2074.720 1702.400 2077.100 1702.680 ;
        RECT 2077.940 1702.400 2080.320 1702.680 ;
        RECT 2081.160 1702.400 2083.080 1702.680 ;
        RECT 2083.920 1702.400 2086.300 1702.680 ;
        RECT 2087.140 1702.400 2089.520 1702.680 ;
        RECT 2090.360 1702.400 2092.280 1702.680 ;
        RECT 2093.120 1702.400 2095.500 1702.680 ;
        RECT 2096.340 1702.400 2098.720 1702.680 ;
        RECT 2099.560 1702.400 2101.480 1702.680 ;
        RECT 2102.320 1702.400 2104.700 1702.680 ;
        RECT 2105.540 1702.400 2107.920 1702.680 ;
        RECT 2108.760 1702.400 2110.680 1702.680 ;
        RECT 2111.520 1702.400 2113.900 1702.680 ;
        RECT 2114.740 1702.400 2117.120 1702.680 ;
        RECT 2117.960 1702.400 2119.880 1702.680 ;
        RECT 2120.720 1702.400 2123.100 1702.680 ;
        RECT 2123.940 1702.400 2125.860 1702.680 ;
        RECT 2126.700 1702.400 2129.080 1702.680 ;
        RECT 2129.920 1702.400 2132.300 1702.680 ;
        RECT 2133.140 1702.400 2135.060 1702.680 ;
        RECT 2135.900 1702.400 2138.280 1702.680 ;
        RECT 2139.120 1702.400 2141.500 1702.680 ;
        RECT 2142.340 1702.400 2144.260 1702.680 ;
        RECT 2145.100 1702.400 2147.480 1702.680 ;
        RECT 2148.320 1702.400 2150.700 1702.680 ;
        RECT 2151.540 1702.400 2153.460 1702.680 ;
        RECT 2154.300 1702.400 2156.680 1702.680 ;
        RECT 2157.520 1702.400 2159.900 1702.680 ;
        RECT 2160.740 1702.400 2162.660 1702.680 ;
        RECT 2163.500 1702.400 2165.880 1702.680 ;
        RECT 2166.720 1702.400 2169.100 1702.680 ;
        RECT 2169.940 1702.400 2171.860 1702.680 ;
        RECT 2172.700 1702.400 2175.080 1702.680 ;
        RECT 2175.920 1702.400 2178.300 1702.680 ;
        RECT 2179.140 1702.400 2181.060 1702.680 ;
        RECT 2181.900 1702.400 2184.280 1702.680 ;
        RECT 2185.120 1702.400 2187.500 1702.680 ;
        RECT 2188.340 1702.400 2190.260 1702.680 ;
        RECT 2191.100 1702.400 2193.480 1702.680 ;
        RECT 2194.320 1702.400 2196.700 1702.680 ;
        RECT 2197.540 1702.400 2199.460 1702.680 ;
        RECT 2200.300 1702.400 2202.680 1702.680 ;
        RECT 2203.520 1702.400 2205.900 1702.680 ;
        RECT 2206.740 1702.400 2208.660 1702.680 ;
        RECT 2209.500 1702.400 2211.880 1702.680 ;
        RECT 2212.720 1702.400 2214.640 1702.680 ;
        RECT 2215.480 1702.400 2217.860 1702.680 ;
        RECT 2218.700 1702.400 2221.080 1702.680 ;
        RECT 2221.920 1702.400 2223.840 1702.680 ;
        RECT 2224.680 1702.400 2227.060 1702.680 ;
        RECT 2227.900 1702.400 2230.280 1702.680 ;
        RECT 2231.120 1702.400 2233.040 1702.680 ;
        RECT 2233.880 1702.400 2236.260 1702.680 ;
        RECT 2237.100 1702.400 2239.480 1702.680 ;
        RECT 2240.320 1702.400 2242.240 1702.680 ;
        RECT 2243.080 1702.400 2245.460 1702.680 ;
        RECT 2246.300 1702.400 2248.680 1702.680 ;
        RECT 2249.520 1702.400 2251.440 1702.680 ;
        RECT 2252.280 1702.400 2254.660 1702.680 ;
        RECT 2255.500 1702.400 2257.880 1702.680 ;
        RECT 2258.720 1702.400 2260.640 1702.680 ;
        RECT 2261.480 1702.400 2263.860 1702.680 ;
        RECT 2264.700 1702.400 2267.080 1702.680 ;
        RECT 2267.920 1702.400 2269.840 1702.680 ;
        RECT 2270.680 1702.400 2273.060 1702.680 ;
        RECT 2273.900 1702.400 2276.280 1702.680 ;
        RECT 2277.120 1702.400 2279.040 1702.680 ;
        RECT 2279.880 1702.400 2282.260 1702.680 ;
        RECT 2283.100 1702.400 2285.480 1702.680 ;
        RECT 2286.320 1702.400 2288.240 1702.680 ;
        RECT 2289.080 1702.400 2291.460 1702.680 ;
        RECT 2292.300 1702.400 2294.680 1702.680 ;
        RECT 2295.520 1702.400 2297.440 1702.680 ;
        RECT 2298.280 1702.400 2300.660 1702.680 ;
        RECT 2301.500 1702.400 2303.420 1702.680 ;
        RECT 2304.260 1702.400 2306.640 1702.680 ;
        RECT 2307.480 1702.400 2309.860 1702.680 ;
        RECT 2310.700 1702.400 2312.620 1702.680 ;
        RECT 2313.460 1702.400 2315.840 1702.680 ;
        RECT 2316.680 1702.400 2319.060 1702.680 ;
        RECT 2319.900 1702.400 2321.820 1702.680 ;
        RECT 2322.660 1702.400 2325.040 1702.680 ;
        RECT 2325.880 1702.400 2328.260 1702.680 ;
        RECT 2329.100 1702.400 2331.020 1702.680 ;
        RECT 2331.860 1702.400 2334.240 1702.680 ;
        RECT 2335.080 1702.400 2337.460 1702.680 ;
        RECT 2338.300 1702.400 2340.220 1702.680 ;
        RECT 2341.060 1702.400 2343.440 1702.680 ;
        RECT 2344.280 1702.400 2346.660 1702.680 ;
        RECT 2347.500 1702.400 2349.420 1702.680 ;
        RECT 2350.260 1702.400 2352.640 1702.680 ;
        RECT 2353.480 1702.400 2355.860 1702.680 ;
        RECT 2356.700 1702.400 2358.620 1702.680 ;
        RECT 2359.460 1702.400 2361.840 1702.680 ;
        RECT 2362.680 1702.400 2365.060 1702.680 ;
        RECT 2365.900 1702.400 2367.820 1702.680 ;
        RECT 2368.660 1702.400 2371.040 1702.680 ;
        RECT 2371.880 1702.400 2374.260 1702.680 ;
        RECT 2375.100 1702.400 2377.020 1702.680 ;
        RECT 2377.860 1702.400 2380.240 1702.680 ;
        RECT 2381.080 1702.400 2383.460 1702.680 ;
        RECT 2384.300 1702.400 2386.220 1702.680 ;
        RECT 2387.060 1702.400 2389.440 1702.680 ;
        RECT 2390.280 1702.400 2392.200 1702.680 ;
        RECT 2393.040 1702.400 2395.420 1702.680 ;
        RECT 2396.260 1702.400 2398.640 1702.680 ;
        RECT 2399.480 1702.400 2401.400 1702.680 ;
        RECT 2402.240 1702.400 2404.620 1702.680 ;
        RECT 2405.460 1702.400 2407.840 1702.680 ;
        RECT 2408.680 1702.400 2410.600 1702.680 ;
        RECT 2411.440 1702.400 2413.820 1702.680 ;
        RECT 2414.660 1702.400 2417.040 1702.680 ;
        RECT 2417.880 1702.400 2419.800 1702.680 ;
        RECT 2420.640 1702.400 2423.020 1702.680 ;
        RECT 2423.860 1702.400 2426.240 1702.680 ;
        RECT 2427.080 1702.400 2429.000 1702.680 ;
        RECT 2429.840 1702.400 2432.220 1702.680 ;
        RECT 2433.060 1702.400 2435.440 1702.680 ;
        RECT 2436.280 1702.400 2438.200 1702.680 ;
        RECT 2439.040 1702.400 2441.420 1702.680 ;
        RECT 2442.260 1702.400 2444.640 1702.680 ;
        RECT 2445.480 1702.400 2447.400 1702.680 ;
        RECT 2448.240 1702.400 2450.620 1702.680 ;
        RECT 2451.460 1702.400 2453.840 1702.680 ;
        RECT 2454.680 1702.400 2456.600 1702.680 ;
        RECT 2457.440 1702.400 2459.820 1702.680 ;
        RECT 2460.660 1702.400 2463.040 1702.680 ;
        RECT 2463.880 1702.400 2465.800 1702.680 ;
        RECT 2466.640 1702.400 2469.020 1702.680 ;
        RECT 2469.860 1702.400 2472.240 1702.680 ;
        RECT 2473.080 1702.400 2475.000 1702.680 ;
        RECT 2475.840 1702.400 2478.220 1702.680 ;
        RECT 2479.060 1702.400 2480.980 1702.680 ;
        RECT 2481.820 1702.400 2484.200 1702.680 ;
        RECT 2485.040 1702.400 2487.420 1702.680 ;
        RECT 2488.260 1702.400 2490.180 1702.680 ;
        RECT 2491.020 1702.400 2493.400 1702.680 ;
        RECT 2494.240 1702.400 2496.620 1702.680 ;
        RECT 2497.460 1702.400 2499.380 1702.680 ;
        RECT 2500.220 1702.400 2502.600 1702.680 ;
        RECT 2503.440 1702.400 2505.820 1702.680 ;
        RECT 2506.660 1702.400 2508.580 1702.680 ;
        RECT 2509.420 1702.400 2511.800 1702.680 ;
        RECT 2512.640 1702.400 2515.020 1702.680 ;
        RECT 2515.860 1702.400 2517.780 1702.680 ;
        RECT 2518.620 1702.400 2521.000 1702.680 ;
        RECT 2521.840 1702.400 2524.220 1702.680 ;
        RECT 2525.060 1702.400 2526.980 1702.680 ;
        RECT 2527.820 1702.400 2530.200 1702.680 ;
        RECT 2531.040 1702.400 2533.420 1702.680 ;
        RECT 2534.260 1702.400 2536.180 1702.680 ;
        RECT 2537.020 1702.400 2539.400 1702.680 ;
        RECT 2540.240 1702.400 2542.620 1702.680 ;
        RECT 2543.460 1702.400 2545.380 1702.680 ;
        RECT 2546.220 1702.400 2548.600 1702.680 ;
        RECT 2549.440 1702.400 2551.820 1702.680 ;
        RECT 2552.660 1702.400 2554.580 1702.680 ;
        RECT 2555.420 1702.400 2557.800 1702.680 ;
        RECT 2558.640 1702.400 2561.020 1702.680 ;
        RECT 2561.860 1702.400 2563.780 1702.680 ;
        RECT 2564.620 1702.400 2567.000 1702.680 ;
        RECT 2567.840 1702.400 2569.760 1702.680 ;
        RECT 2570.600 1702.400 2572.980 1702.680 ;
        RECT 2573.820 1702.400 2576.200 1702.680 ;
        RECT 2577.040 1702.400 2578.960 1702.680 ;
        RECT 2579.800 1702.400 2582.180 1702.680 ;
        RECT 2583.020 1702.400 2585.400 1702.680 ;
        RECT 2586.240 1702.400 2588.160 1702.680 ;
        RECT 2589.000 1702.400 2591.380 1702.680 ;
        RECT 2592.220 1702.400 2594.600 1702.680 ;
        RECT 2595.440 1702.400 2597.360 1702.680 ;
        RECT 2598.200 1702.400 2600.580 1702.680 ;
        RECT 2601.420 1702.400 2603.800 1702.680 ;
        RECT 2604.640 1702.400 2606.560 1702.680 ;
        RECT 2607.400 1702.400 2609.780 1702.680 ;
        RECT 2610.620 1702.400 2613.000 1702.680 ;
        RECT 2613.840 1702.400 2615.760 1702.680 ;
        RECT 2616.600 1702.400 2618.980 1702.680 ;
        RECT 2619.820 1702.400 2622.200 1702.680 ;
        RECT 2623.040 1702.400 2624.960 1702.680 ;
        RECT 2625.800 1702.400 2628.180 1702.680 ;
        RECT 2629.020 1702.400 2631.400 1702.680 ;
        RECT 2632.240 1702.400 2634.160 1702.680 ;
        RECT 2635.000 1702.400 2637.380 1702.680 ;
        RECT 2638.220 1702.400 2640.600 1702.680 ;
        RECT 2641.440 1702.400 2643.360 1702.680 ;
        RECT 2644.200 1702.400 2646.580 1702.680 ;
      LAYER met3 ;
        RECT 1152.755 1710.715 2630.390 3188.005 ;
      LAYER met4 ;
        RECT 1169.590 1710.640 1171.190 3188.080 ;
      LAYER met4 ;
        RECT 1173.685 1710.640 1174.020 3188.080 ;
        RECT 1177.020 1710.640 1192.020 3188.080 ;
        RECT 1195.020 1710.640 1210.020 3188.080 ;
        RECT 1213.020 1710.640 1228.020 3188.080 ;
        RECT 1231.020 3045.290 1245.990 3188.080 ;
        RECT 1248.390 3150.690 1264.020 3188.080 ;
        RECT 1248.570 3149.510 1264.020 3150.690 ;
        RECT 1248.390 3075.890 1264.020 3149.510 ;
        RECT 1248.570 3074.710 1264.020 3075.890 ;
        RECT 1231.020 3044.110 1245.550 3045.290 ;
        RECT 1231.020 1710.640 1245.990 3044.110 ;
        RECT 1248.390 1712.490 1264.020 3074.710 ;
        RECT 1248.570 1711.310 1264.020 1712.490 ;
        RECT 1248.390 1710.640 1264.020 1711.310 ;
        RECT 1267.020 1710.640 1282.020 3188.080 ;
        RECT 1285.020 1710.640 1300.020 3188.080 ;
        RECT 1303.020 1710.640 1318.020 3188.080 ;
        RECT 1321.020 1710.640 1354.020 3188.080 ;
        RECT 1357.020 1710.640 1372.020 3188.080 ;
        RECT 1375.020 1710.640 1390.020 3188.080 ;
        RECT 1393.020 1710.640 1408.020 3188.080 ;
        RECT 1411.020 1710.640 1444.020 3188.080 ;
        RECT 1447.020 1710.640 1462.020 3188.080 ;
        RECT 1465.020 1710.640 1480.020 3188.080 ;
        RECT 1483.020 1710.640 1498.020 3188.080 ;
        RECT 1501.020 1710.640 1534.020 3188.080 ;
        RECT 1537.020 1710.640 1552.020 3188.080 ;
        RECT 1555.020 1710.640 1570.020 3188.080 ;
        RECT 1573.020 1710.640 1588.020 3188.080 ;
        RECT 1591.020 1710.640 1624.020 3188.080 ;
        RECT 1627.020 1710.640 1642.020 3188.080 ;
        RECT 1645.020 1710.640 1660.020 3188.080 ;
        RECT 1663.020 1710.640 1678.020 3188.080 ;
        RECT 1681.020 1710.640 1714.020 3188.080 ;
        RECT 1717.020 1710.640 1732.020 3188.080 ;
        RECT 1735.020 1710.640 1750.020 3188.080 ;
        RECT 1753.020 1710.640 1768.020 3188.080 ;
        RECT 1771.020 1710.640 1804.020 3188.080 ;
        RECT 1807.020 1710.640 1822.020 3188.080 ;
        RECT 1825.020 1710.640 1840.020 3188.080 ;
        RECT 1843.020 1710.640 1858.020 3188.080 ;
        RECT 1861.020 1710.640 1894.020 3188.080 ;
        RECT 1897.020 1710.640 1912.020 3188.080 ;
        RECT 1915.020 1710.640 1930.020 3188.080 ;
        RECT 1933.020 1710.640 1948.020 3188.080 ;
        RECT 1951.020 1710.640 1984.020 3188.080 ;
        RECT 1987.020 1710.640 2002.020 3188.080 ;
        RECT 2005.020 1710.640 2020.020 3188.080 ;
        RECT 2023.020 1710.640 2038.020 3188.080 ;
        RECT 2041.020 1710.640 2074.020 3188.080 ;
        RECT 2077.020 1710.640 2092.020 3188.080 ;
        RECT 2095.020 1710.640 2110.020 3188.080 ;
        RECT 2113.020 1710.640 2128.020 3188.080 ;
        RECT 2131.020 1710.640 2164.020 3188.080 ;
        RECT 2167.020 1710.640 2182.020 3188.080 ;
        RECT 2185.020 1710.640 2200.020 3188.080 ;
        RECT 2203.020 1710.640 2218.020 3188.080 ;
        RECT 2221.020 1710.640 2254.020 3188.080 ;
        RECT 2257.020 1710.640 2272.020 3188.080 ;
        RECT 2275.020 1710.640 2290.020 3188.080 ;
        RECT 2293.020 1710.640 2308.020 3188.080 ;
        RECT 2311.020 1710.640 2344.020 3188.080 ;
        RECT 2347.020 1710.640 2362.020 3188.080 ;
        RECT 2365.020 1710.640 2380.020 3188.080 ;
        RECT 2383.020 1710.640 2398.020 3188.080 ;
        RECT 2401.020 1710.640 2434.020 3188.080 ;
        RECT 2437.020 1710.640 2452.020 3188.080 ;
        RECT 2455.020 1710.640 2470.020 3188.080 ;
        RECT 2473.020 1710.640 2488.020 3188.080 ;
        RECT 2491.020 1710.640 2524.020 3188.080 ;
        RECT 2527.020 1710.640 2542.020 3188.080 ;
        RECT 2545.020 1710.640 2560.020 3188.080 ;
        RECT 2563.020 1710.640 2578.020 3188.080 ;
        RECT 2581.020 1710.640 2614.020 3188.080 ;
        RECT 2617.020 1710.640 2630.390 3188.080 ;
  END
END user_project_wrapper
END LIBRARY

